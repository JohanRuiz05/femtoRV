* GTKWave TIM to ngspice PWL converter
* Source: femto.tim
* Time Scale: 1e-12 seconds
* VDD Level: 3.3V
* Signals: 4

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt 
.tran 10000ns 200us
.print tran format=raw file=femto_cir.raw  v(*)
* Fuentes de alimentación
Vvdd VPWR 0 DC 3.3
Vgnd VGND 0 DC 0

* clk - 89369 transitions
V_clk clk 0 PWL(0 0 -8e-08 0 2e-08 3.3 -6e-08 3.3 4e-08 0 -4e-08 0 6e-08 3.3 -1.9999999999999994e-08 3.3 8e-08 0 0.0 0 1e-07 3.3 1.9999999999999994e-08 3.3 1.2e-07 0 4.0000000000000014e-08 0 1.4e-07 3.3 6.000000000000001e-08 3.3 1.6e-07 0 8e-08 0 1.8e-07 3.3 1e-07 3.3 2e-07 0 1.2e-07 0 2.1999999999999998e-07 3.3 1.3999999999999998e-07 3.3 2.4e-07 0 1.6e-07 0 2.6e-07 3.3 1.8000000000000002e-07 3.3 2.8e-07 0 2e-07 0 3e-07 3.3 2.2e-07 3.3 3.2e-07 0 2.4e-07 0 3.4e-07 3.3 2.6e-07 3.3 3.6e-07 0 2.8e-07 0 3.8e-07 3.3 3e-07 3.3 4e-07 0 3.2e-07 0 4.2e-07 3.3 3.4e-07 3.3 4.3999999999999997e-07 0 3.6e-07 0 4.6e-07 3.3 3.7999999999999996e-07 3.3 4.8e-07 0 4e-07 0 5e-07 3.3 4.2e-07 3.3 5.2e-07 0 4.4e-07 0 5.4e-07 3.3 4.6000000000000004e-07 3.3 5.6e-07 0 4.8e-07 0 5.8e-07 3.3 5e-07 3.3 6e-07 0 5.2e-07 0 6.2e-07 3.3 5.4e-07 3.3 6.4e-07 0 5.6e-07 0 6.6e-07 3.3 5.8e-07 3.3 6.8e-07 0 6e-07 0 7e-07 3.3 6.2e-07 3.3 7.2e-07 0 6.4e-07 0 7.4e-07 3.3 6.6e-07 3.3 7.6e-07 0 6.8e-07 0 7.799999999999999e-07 3.3 7e-07 3.3 8e-07 0 7.2e-07 0 8.2e-07 3.3 7.4e-07 3.3 8.4e-07 0 7.6e-07 0 8.6e-07 3.3 7.799999999999999e-07 3.3 8.799999999999999e-07 0 8e-07 0 9e-07 3.3 8.2e-07 3.3 9.2e-07 0 8.4e-07 0 9.4e-07 3.3 8.599999999999999e-07 3.3 9.6e-07 0 8.799999999999999e-07 0 9.8e-07 3.3 9e-07 3.3 1e-06 0 9.2e-07 0 1.02e-06 3.3 9.4e-07 3.3 1.04e-06 0 9.600000000000001e-07 0 1.06e-06 3.3 9.8e-07 3.3 1.08e-06 0 1.0000000000000002e-06 0 1.1e-06 3.3 1.02e-06 3.3 1.12e-06 0 1.0399999999999998e-06 0 1.1399999999999999e-06 3.3 1.06e-06 3.3 1.16e-06 0 1.0799999999999998e-06 0 1.18e-06 3.3 1.1e-06 3.3 1.2e-06 0 1.1199999999999999e-06 0 1.22e-06 3.3 1.14e-06 3.3 1.24e-06 0 1.16e-06 0 1.26e-06 3.3 1.1800000000000001e-06 3.3 1.28e-06 0 1.2e-06 0 1.3e-06 3.3 1.2200000000000002e-06 3.3 1.32e-06 0 1.24e-06 0 1.3399999999999999e-06 3.3 1.2599999999999998e-06 3.3 1.36e-06 0 1.28e-06 0 1.38e-06 3.3 1.2999999999999998e-06 3.3 1.4e-06 0 1.32e-06 0 1.42e-06 3.3 1.3399999999999999e-06 3.3 1.44e-06 0 1.3600000000000001e-06 0 1.46e-06 3.3 1.38e-06 3.3 1.48e-06 0 1.4000000000000001e-06 0 1.5e-06 3.3 1.42e-06 3.3 1.52e-06 0 1.4399999999999998e-06 0 1.5399999999999999e-06 3.3 1.46e-06 3.3 1.5599999999999999e-06 0 1.4799999999999998e-06 0 1.58e-06 3.3 1.5e-06 3.3 1.6e-06 0 1.5199999999999998e-06 0 1.62e-06 3.3 1.54e-06 3.3 1.64e-06 0 1.5599999999999999e-06 0 1.66e-06 3.3 1.5800000000000001e-06 3.3 1.68e-06 0 1.6e-06 0 1.7e-06 3.3 1.6200000000000002e-06 3.3 1.72e-06 0 1.64e-06 0 1.74e-06 3.3 1.6599999999999998e-06 3.3 1.7599999999999999e-06 0 1.68e-06 0 1.78e-06 3.3 1.6999999999999998e-06 3.3 1.8e-06 0 1.72e-06 0 1.82e-06 3.3 1.7399999999999999e-06 3.3 1.84e-06 0 1.76e-06 0 1.86e-06 3.3 1.78e-06 3.3 1.88e-06 0 1.8000000000000001e-06 0 1.9e-06 3.3 1.82e-06 3.3 1.92e-06 0 1.8400000000000002e-06 0 1.94e-06 3.3 1.86e-06 3.3 1.96e-06 0 1.8800000000000002e-06 0 1.98e-06 3.3 1.9e-06 3.3 2e-06 0 1.9200000000000003e-06 0 2.02e-06 3.3 1.94e-06 3.3 2.04e-06 0 1.96e-06 0 2.0599999999999998e-06 3.3 1.98e-06 3.3 2.08e-06 0 2e-06 0 2.1e-06 3.3 2.02e-06 3.3 2.12e-06 0 2.04e-06 0 2.14e-06 3.3 2.06e-06 3.3 2.16e-06 0 2.08e-06 0 2.18e-06 3.3 2.1000000000000002e-06 3.3 2.2e-06 0 2.12e-06 0 2.22e-06 3.3 2.1400000000000003e-06 3.3 2.24e-06 0 2.16e-06 0 2.26e-06 3.3 2.18e-06 3.3 2.2799999999999998e-06 0 2.2e-06 0 2.3e-06 3.3 2.22e-06 3.3 2.32e-06 0 2.24e-06 0 2.34e-06 3.3 2.26e-06 3.3 2.36e-06 0 2.28e-06 0 2.38e-06 3.3 2.3e-06 3.3 2.4e-06 0 2.3200000000000002e-06 0 2.42e-06 3.3 2.34e-06 3.3 2.44e-06 0 2.36e-06 0 2.4599999999999997e-06 3.3 2.38e-06 3.3 2.48e-06 0 2.4e-06 0 2.4999999999999998e-06 3.3 2.42e-06 3.3 2.52e-06 0 2.44e-06 0 2.54e-06 3.3 2.46e-06 3.3 2.56e-06 0 2.48e-06 0 2.58e-06 3.3 2.5e-06 3.3 2.6e-06 0 2.52e-06 0 2.62e-06 3.3 2.5400000000000002e-06 3.3 2.64e-06 0 2.56e-06 0 2.66e-06 3.3 2.58e-06 3.3 2.6799999999999998e-06 0 2.6e-06 0 2.7e-06 3.3 2.62e-06 3.3 2.72e-06 0 2.64e-06 0 2.74e-06 3.3 2.66e-06 3.3 2.76e-06 0 2.68e-06 0 2.78e-06 3.3 2.7e-06 3.3 2.8e-06 0 2.7200000000000002e-06 0 2.82e-06 3.3 2.74e-06 3.3 2.84e-06 0 2.7600000000000003e-06 0 2.86e-06 3.3 2.78e-06 3.3 2.88e-06 0 2.8e-06 0 2.8999999999999998e-06 3.3 2.82e-06 3.3 2.92e-06 0 2.84e-06 0 2.94e-06 3.3 2.86e-06 3.3 2.96e-06 0 2.88e-06 0 2.98e-06 3.3 2.9e-06 3.3 3e-06 0 2.92e-06 0 3.02e-06 3.3 2.9400000000000002e-06 3.3 3.04e-06 0 2.96e-06 0 3.06e-06 3.3 2.98e-06 3.3 3.0799999999999997e-06 0 3e-06 0 3.1e-06 3.3 3.02e-06 3.3 3.1199999999999998e-06 0 3.04e-06 0 3.14e-06 3.3 3.06e-06 3.3 3.16e-06 0 3.08e-06 0 3.18e-06 3.3 3.1e-06 3.3 3.2e-06 0 3.12e-06 0 3.22e-06 3.3 3.14e-06 3.3 3.24e-06 0 3.1600000000000002e-06 0 3.26e-06 3.3 3.18e-06 3.3 3.28e-06 0 3.2e-06 0 3.2999999999999997e-06 3.3 3.22e-06 3.3 3.32e-06 0 3.24e-06 0 3.3399999999999998e-06 3.3 3.26e-06 3.3 3.36e-06 0 3.28e-06 0 3.38e-06 3.3 3.3e-06 3.3 3.4e-06 0 3.32e-06 0 3.42e-06 3.3 3.34e-06 3.3 3.44e-06 0 3.36e-06 0 3.46e-06 3.3 3.3800000000000002e-06 3.3 3.48e-06 0 3.4e-06 0 3.5e-06 3.3 3.42e-06 3.3 3.5199999999999998e-06 0 3.44e-06 0 3.54e-06 3.3 3.46e-06 3.3 3.56e-06 0 3.48e-06 0 3.58e-06 3.3 3.5e-06 3.3 3.6e-06 0 3.52e-06 0 3.62e-06 3.3 3.54e-06 3.3 3.64e-06 0 3.5600000000000002e-06 0 3.66e-06 3.3 3.58e-06 3.3 3.68e-06 0 3.6e-06 0 3.6999999999999997e-06 3.3 3.62e-06 3.3 3.72e-06 0 3.64e-06 0 3.7399999999999998e-06 3.3 3.66e-06 3.3 3.76e-06 0 3.68e-06 0 3.78e-06 3.3 3.7e-06 3.3 3.8e-06 0 3.72e-06 0 3.82e-06 3.3 3.7399999999999998e-06 3.3 3.84e-06 0 3.7600000000000004e-06 0 3.86e-06 3.3 3.7800000000000002e-06 3.3 3.88e-06 0 3.8e-06 0 3.9e-06 3.3 3.82e-06 3.3 3.92e-06 0 3.84e-06 0 3.9399999999999995e-06 3.3 3.86e-06 3.3 3.96e-06 0 3.88e-06 0 3.98e-06 3.3 3.9e-06 3.3 4e-06 0 3.92e-06 0 4.02e-06 3.3 3.94e-06 3.3 4.04e-06 0 3.96e-06 0 4.06e-06 3.3 3.98e-06 3.3 4.08e-06 0 4e-06 0 4.1e-06 3.3 4.02e-06 3.3 4.1199999999999995e-06 0 4.04e-06 0 4.14e-06 3.3 4.06e-06 3.3 4.16e-06 0 4.08e-06 0 4.18e-06 3.3 4.1e-06 3.3 4.2e-06 0 4.12e-06 0 4.22e-06 3.3 4.14e-06 3.3 4.24e-06 0 4.16e-06 0 4.26e-06 3.3 4.18e-06 3.3 4.28e-06 0 4.2000000000000004e-06 0 4.3e-06 3.3 4.22e-06 3.3 4.32e-06 0 4.24e-06 0 4.34e-06 3.3 4.26e-06 3.3 4.36e-06 0 4.28e-06 0 4.3799999999999996e-06 3.3 4.3e-06 3.3 4.4e-06 0 4.32e-06 0 4.42e-06 3.3 4.34e-06 3.3 4.44e-06 0 4.36e-06 0 4.46e-06 3.3 4.38e-06 3.3 4.48e-06 0 4.4e-06 0 4.5e-06 3.3 4.42e-06 3.3 4.52e-06 0 4.44e-06 0 4.54e-06 3.3 4.46e-06 3.3 4.5599999999999995e-06 0 4.48e-06 0 4.58e-06 3.3 4.5e-06 3.3 4.6e-06 0 4.52e-06 0 4.62e-06 3.3 4.54e-06 3.3 4.64e-06 0 4.56e-06 0 4.66e-06 3.3 4.58e-06 3.3 4.68e-06 0 4.6e-06 0 4.7e-06 3.3 4.62e-06 3.3 4.72e-06 0 4.64e-06 0 4.7399999999999995e-06 3.3 4.66e-06 3.3 4.76e-06 0 4.68e-06 0 4.78e-06 3.3 4.7e-06 3.3 4.8e-06 0 4.72e-06 0 4.82e-06 3.3 4.74e-06 3.3 4.84e-06 0 4.76e-06 0 4.86e-06 3.3 4.78e-06 3.3 4.88e-06 0 4.8e-06 0 4.9e-06 3.3 4.82e-06 3.3 4.9199999999999995e-06 0 4.84e-06 0 4.94e-06 3.3 4.86e-06 3.3 4.96e-06 0 4.88e-06 0 4.98e-06 3.3 4.9e-06 3.3 4.9999999999999996e-06 0 4.92e-06 0 5.02e-06 3.3 4.94e-06 3.3 5.04e-06 0 4.96e-06 0 5.06e-06 3.3 4.98e-06 3.3 5.08e-06 0 5e-06 0 5.1e-06 3.3 5.02e-06 3.3 5.12e-06 0 5.04e-06 0 5.14e-06 3.3 5.06e-06 3.3 5.16e-06 0 5.08e-06 0 5.1799999999999995e-06 3.3 5.1e-06 3.3 5.2e-06 0 5.12e-06 0 5.22e-06 3.3 5.14e-06 3.3 5.24e-06 0 5.16e-06 0 5.26e-06 3.3 5.18e-06 3.3 5.28e-06 0 5.2e-06 0 5.3e-06 3.3 5.22e-06 3.3 5.32e-06 0 5.24e-06 0 5.34e-06 3.3 5.26e-06 3.3 5.3599999999999995e-06 0 5.28e-06 0 5.38e-06 3.3 5.3e-06 3.3 5.4e-06 0 5.32e-06 0 5.42e-06 3.3 5.34e-06 3.3 5.44e-06 0 5.36e-06 0 5.46e-06 3.3 5.38e-06 3.3 5.48e-06 0 5.4e-06 0 5.5e-06 3.3 5.42e-06 3.3 5.52e-06 0 5.44e-06 0 5.5399999999999995e-06 3.3 5.46e-06 3.3 5.56e-06 0 5.48e-06 0 5.58e-06 3.3 5.5e-06 3.3 5.6e-06 0 5.52e-06 0 5.6199999999999996e-06 3.3 5.54e-06 3.3 5.64e-06 0 5.56e-06 0 5.66e-06 3.3 5.58e-06 3.3 5.68e-06 0 5.6e-06 0 5.7e-06 3.3 5.62e-06 3.3 5.72e-06 0 5.64e-06 0 5.74e-06 3.3 5.66e-06 3.3 5.76e-06 0 5.68e-06 0 5.78e-06 3.3 5.7e-06 3.3 5.7999999999999995e-06 0 5.72e-06 0 5.82e-06 3.3 5.74e-06 3.3 5.84e-06 0 5.76e-06 0 5.86e-06 3.3 5.78e-06 3.3 5.88e-06 0 5.8e-06 0 5.9e-06 3.3 5.82e-06 3.3 5.92e-06 0 5.84e-06 0 5.94e-06 3.3 5.86e-06 3.3 5.96e-06 0 5.88e-06 0 5.9799999999999995e-06 3.3 5.9e-06 3.3 6e-06 0 5.92e-06 0 6.02e-06 3.3 5.94e-06 3.3 6.04e-06 0 5.96e-06 0 6.06e-06 3.3 5.98e-06 3.3 6.08e-06 0 6e-06 0 6.1e-06 3.3 6.02e-06 3.3 6.12e-06 0 6.04e-06 0 6.14e-06 3.3 6.06e-06 3.3 6.1599999999999995e-06 0 6.08e-06 0 6.18e-06 3.3 6.1e-06 3.3 6.2e-06 0 6.12e-06 0 6.22e-06 3.3 6.14e-06 3.3 6.2399999999999995e-06 0 6.16e-06 0 6.26e-06 3.3 6.18e-06 3.3 6.28e-06 0 6.2e-06 0 6.3e-06 3.3 6.22e-06 3.3 6.32e-06 0 6.24e-06 0 6.34e-06 3.3 6.26e-06 3.3 6.36e-06 0 6.28e-06 0 6.38e-06 3.3 6.3e-06 3.3 6.4e-06 0 6.32e-06 0 6.4199999999999995e-06 3.3 6.34e-06 3.3 6.44e-06 0 6.36e-06 0 6.46e-06 3.3 6.38e-06 3.3 6.48e-06 0 6.4e-06 0 6.5e-06 3.3 6.42e-06 3.3 6.52e-06 0 6.44e-06 0 6.54e-06 3.3 6.46e-06 3.3 6.56e-06 0 6.48e-06 0 6.58e-06 3.3 6.5e-06 3.3 6.5999999999999995e-06 0 6.52e-06 0 6.62e-06 3.3 6.54e-06 3.3 6.64e-06 0 6.56e-06 0 6.66e-06 3.3 6.58e-06 3.3 6.6799999999999996e-06 0 6.6e-06 0 6.7e-06 3.3 6.62e-06 3.3 6.72e-06 0 6.64e-06 0 6.74e-06 3.3 6.66e-06 3.3 6.76e-06 0 6.6799999999999996e-06 0 6.7799999999999995e-06 3.3 6.7e-06 3.3 6.8e-06 0 6.72e-06 0 6.82e-06 3.3 6.74e-06 3.3 6.84e-06 0 6.76e-06 0 6.8599999999999995e-06 3.3 6.78e-06 3.3 6.88e-06 0 6.8e-06 0 6.9e-06 3.3 6.82e-06 3.3 6.92e-06 0 6.84e-06 0 6.94e-06 3.3 6.86e-06 3.3 6.96e-06 0 6.88e-06 0 6.98e-06 3.3 6.9e-06 3.3 7e-06 0 6.92e-06 0 7.02e-06 3.3 6.94e-06 3.3 7.0399999999999995e-06 0 6.96e-06 0 7.06e-06 3.3 6.98e-06 3.3 7.08e-06 0 7e-06 0 7.1e-06 3.3 7.02e-06 3.3 7.12e-06 0 7.04e-06 0 7.14e-06 3.3 7.06e-06 3.3 7.16e-06 0 7.08e-06 0 7.18e-06 3.3 7.1e-06 3.3 7.2e-06 0 7.12e-06 0 7.2199999999999995e-06 3.3 7.14e-06 3.3 7.24e-06 0 7.16e-06 0 7.26e-06 3.3 7.18e-06 3.3 7.28e-06 0 7.2e-06 0 7.2999999999999996e-06 3.3 7.22e-06 3.3 7.32e-06 0 7.24e-06 0 7.34e-06 3.3 7.26e-06 3.3 7.36e-06 0 7.28e-06 0 7.38e-06 3.3 7.2999999999999996e-06 3.3 7.3999999999999995e-06 0 7.32e-06 0 7.42e-06 3.3 7.34e-06 3.3 7.44e-06 0 7.36e-06 0 7.46e-06 3.3 7.38e-06 3.3 7.4799999999999995e-06 0 7.4e-06 0 7.5e-06 3.3 7.42e-06 3.3 7.52e-06 0 7.44e-06 0 7.54e-06 3.3 7.46e-06 3.3 7.56e-06 0 7.4799999999999995e-06 0 7.5799999999999994e-06 3.3 7.5e-06 3.3 7.6e-06 0 7.52e-06 0 7.62e-06 3.3 7.54e-06 3.3 7.64e-06 0 7.56e-06 0 7.66e-06 3.3 7.5799999999999994e-06 3.3 7.68e-06 0 7.599999999999999e-06 0 7.699999999999999e-06 3.3 7.620000000000001e-06 3.3 7.72e-06 0 7.64e-06 0 7.74e-06 3.3 7.66e-06 3.3 7.76e-06 0 7.68e-06 0 7.78e-06 3.3 7.699999999999999e-06 3.3 7.8e-06 0 7.719999999999999e-06 0 7.82e-06 3.3 7.739999999999999e-06 3.3 7.84e-06 0 7.759999999999999e-06 0 7.86e-06 3.3 7.779999999999998e-06 3.3 7.879999999999999e-06 0 7.8e-06 0 7.9e-06 3.3 7.82e-06 3.3 7.92e-06 0 7.84e-06 0 7.94e-06 3.3 7.86e-06 3.3 7.96e-06 0 7.879999999999999e-06 0 7.98e-06 3.3 7.899999999999999e-06 3.3 8e-06 0 7.919999999999999e-06 0 8.02e-06 3.3 7.939999999999999e-06 3.3 8.04e-06 0 7.959999999999998e-06 0 8.059999999999999e-06 3.3 7.98e-06 3.3 8.08e-06 0 8e-06 0 8.1e-06 3.3 8.02e-06 3.3 8.12e-06 0 8.04e-06 0 8.14e-06 3.3 8.059999999999999e-06 3.3 8.16e-06 0 8.079999999999999e-06 0 8.18e-06 3.3 8.099999999999999e-06 3.3 8.2e-06 0 8.119999999999998e-06 0 8.22e-06 3.3 8.139999999999998e-06 3.3 8.239999999999999e-06 0 8.16e-06 0 8.26e-06 3.3 8.18e-06 3.3 8.28e-06 0 8.2e-06 0 8.3e-06 3.3 8.22e-06 3.3 8.32e-06 0 8.239999999999999e-06 0 8.34e-06 3.3 8.259999999999999e-06 3.3 8.36e-06 0 8.279999999999999e-06 0 8.38e-06 3.3 8.299999999999998e-06 3.3 8.4e-06 0 8.319999999999998e-06 0 8.419999999999999e-06 3.3 8.34e-06 3.3 8.44e-06 0 8.36e-06 0 8.46e-06 3.3 8.38e-06 3.3 8.48e-06 0 8.4e-06 0 8.5e-06 3.3 8.419999999999999e-06 3.3 8.52e-06 0 8.439999999999999e-06 0 8.54e-06 3.3 8.459999999999999e-06 3.3 8.56e-06 0 8.479999999999998e-06 0 8.58e-06 3.3 8.5e-06 3.3 8.6e-06 0 8.52e-06 0 8.62e-06 3.3 8.54e-06 3.3 8.64e-06 0 8.56e-06 0 8.66e-06 3.3 8.58e-06 3.3 8.68e-06 0 8.599999999999999e-06 0 8.7e-06 3.3 8.619999999999999e-06 3.3 8.72e-06 0 8.639999999999999e-06 0 8.74e-06 3.3 8.659999999999998e-06 3.3 8.759999999999999e-06 0 8.68e-06 0 8.78e-06 3.3 8.7e-06 3.3 8.8e-06 0 8.72e-06 0 8.82e-06 3.3 8.74e-06 3.3 8.84e-06 0 8.759999999999999e-06 0 8.86e-06 3.3 8.779999999999999e-06 3.3 8.88e-06 0 8.799999999999999e-06 0 8.9e-06 3.3 8.819999999999999e-06 3.3 8.92e-06 0 8.839999999999998e-06 0 8.939999999999999e-06 3.3 8.86e-06 3.3 8.96e-06 0 8.88e-06 0 8.98e-06 3.3 8.9e-06 3.3 9e-06 0 8.92e-06 0 9.02e-06 3.3 8.939999999999999e-06 3.3 9.04e-06 0 8.959999999999999e-06 0 9.06e-06 3.3 8.979999999999999e-06 3.3 9.08e-06 0 8.999999999999999e-06 0 9.1e-06 3.3 9.019999999999998e-06 3.3 9.119999999999999e-06 0 9.04e-06 0 9.14e-06 3.3 9.06e-06 3.3 9.16e-06 0 9.08e-06 0 9.18e-06 3.3 9.1e-06 3.3 9.2e-06 0 9.119999999999999e-06 0 9.22e-06 3.3 9.139999999999999e-06 3.3 9.24e-06 0 9.159999999999999e-06 0 9.26e-06 3.3 9.179999999999999e-06 3.3 9.28e-06 0 9.199999999999998e-06 0 9.299999999999999e-06 3.3 9.22e-06 3.3 9.32e-06 0 9.24e-06 0 9.34e-06 3.3 9.26e-06 3.3 9.36e-06 0 9.28e-06 0 9.38e-06 3.3 9.299999999999999e-06 3.3 9.4e-06 0 9.319999999999999e-06 0 9.42e-06 3.3 9.339999999999999e-06 3.3 9.44e-06 0 9.359999999999998e-06 0 9.46e-06 3.3 9.379999999999998e-06 3.3 9.479999999999999e-06 0 9.4e-06 0 9.5e-06 3.3 9.42e-06 3.3 9.52e-06 0 9.44e-06 0 9.54e-06 3.3 9.46e-06 3.3 9.56e-06 0 9.479999999999999e-06 0 9.58e-06 3.3 9.499999999999999e-06 3.3 9.6e-06 0 9.519999999999999e-06 0 9.62e-06 3.3 9.539999999999998e-06 3.3 9.64e-06 0 9.559999999999998e-06 0 9.659999999999999e-06 3.3 9.58e-06 3.3 9.68e-06 0 9.6e-06 0 9.7e-06 3.3 9.62e-06 3.3 9.72e-06 0 9.64e-06 0 9.74e-06 3.3 9.659999999999999e-06 3.3 9.76e-06 0 9.679999999999999e-06 0 9.78e-06 3.3 9.699999999999999e-06 3.3 9.8e-06 0 9.719999999999998e-06 0 9.82e-06 3.3 9.739999999999998e-06 3.3 9.839999999999999e-06 0 9.76e-06 0 9.86e-06 3.3 9.78e-06 3.3 9.88e-06 0 9.8e-06 0 9.9e-06 3.3 9.82e-06 3.3 9.92e-06 0 9.839999999999999e-06 0 9.94e-06 3.3 9.859999999999999e-06 3.3 9.96e-06 0 9.879999999999999e-06 0 9.98e-06 3.3 9.899999999999998e-06 3.3 9.999999999999999e-06 0 9.92e-06 0 1.002e-05 3.3 9.94e-06 3.3 1.004e-05 0 9.96e-06 0 1.006e-05 3.3 9.98e-06 3.3 1.008e-05 0 9.999999999999999e-06 0 1.01e-05 3.3 1.0019999999999999e-05 3.3 1.012e-05 0 1.0039999999999999e-05 0 1.014e-05 3.3 1.0059999999999999e-05 3.3 1.016e-05 0 1.0079999999999998e-05 0 1.0179999999999999e-05 3.3 1.01e-05 3.3 1.02e-05 0 1.012e-05 0 1.022e-05 3.3 1.014e-05 3.3 1.024e-05 0 1.016e-05 0 1.026e-05 3.3 1.0179999999999999e-05 3.3 1.028e-05 0 1.0199999999999999e-05 0 1.03e-05 3.3 1.0219999999999999e-05 3.3 1.032e-05 0 1.0239999999999999e-05 0 1.034e-05 3.3 1.0259999999999998e-05 3.3 1.0359999999999999e-05 0 1.028e-05 0 1.038e-05 3.3 1.03e-05 3.3 1.04e-05 0 1.032e-05 0 1.042e-05 3.3 1.034e-05 3.3 1.044e-05 0 1.0359999999999999e-05 0 1.046e-05 3.3 1.0379999999999999e-05 3.3 1.048e-05 0 1.0399999999999999e-05 0 1.05e-05 3.3 1.0419999999999998e-05 3.3 1.052e-05 0 1.0439999999999998e-05 0 1.0539999999999999e-05 3.3 1.046e-05 3.3 1.056e-05 0 1.048e-05 0 1.058e-05 3.3 1.05e-05 3.3 1.06e-05 0 1.052e-05 0 1.062e-05 3.3 1.0539999999999999e-05 3.3 1.064e-05 0 1.0559999999999999e-05 0 1.066e-05 3.3 1.0579999999999999e-05 3.3 1.068e-05 0 1.0599999999999998e-05 0 1.07e-05 3.3 1.0619999999999998e-05 3.3 1.0719999999999999e-05 0 1.064e-05 0 1.074e-05 3.3 1.066e-05 3.3 1.076e-05 0 1.068e-05 0 1.078e-05 3.3 1.07e-05 3.3 1.08e-05 0 1.0719999999999999e-05 0 1.082e-05 3.3 1.0739999999999999e-05 3.3 1.084e-05 0 1.0759999999999999e-05 0 1.086e-05 3.3 1.0779999999999998e-05 3.3 1.088e-05 0 1.0799999999999998e-05 0 1.0899999999999999e-05 3.3 1.082e-05 3.3 1.092e-05 0 1.084e-05 0 1.094e-05 3.3 1.086e-05 3.3 1.096e-05 0 1.088e-05 0 1.098e-05 3.3 1.0899999999999999e-05 3.3 1.1e-05 0 1.0919999999999999e-05 0 1.102e-05 3.3 1.0939999999999999e-05 3.3 1.104e-05 0 1.0959999999999998e-05 0 1.1059999999999999e-05 3.3 1.0979999999999998e-05 3.3 1.1079999999999999e-05 0 1.1e-05 0 1.11e-05 3.3 1.102e-05 3.3 1.112e-05 0 1.104e-05 0 1.114e-05 3.3 1.1059999999999999e-05 3.3 1.116e-05 0 1.1079999999999999e-05 0 1.118e-05 3.3 1.1099999999999999e-05 3.3 1.12e-05 0 1.1119999999999999e-05 0 1.122e-05 3.3 1.1139999999999998e-05 3.3 1.1239999999999999e-05 0 1.116e-05 0 1.126e-05 3.3 1.118e-05 3.3 1.128e-05 0 1.12e-05 0 1.13e-05 3.3 1.122e-05 3.3 1.132e-05 0 1.1239999999999999e-05 0 1.134e-05 3.3 1.1259999999999999e-05 3.3 1.136e-05 0 1.1279999999999999e-05 0 1.138e-05 3.3 1.1299999999999999e-05 3.3 1.14e-05 0 1.1319999999999998e-05 0 1.1419999999999999e-05 3.3 1.134e-05 3.3 1.144e-05 0 1.136e-05 0 1.146e-05 3.3 1.138e-05 3.3 1.148e-05 0 1.14e-05 0 1.15e-05 3.3 1.1419999999999999e-05 3.3 1.152e-05 0 1.1439999999999999e-05 0 1.154e-05 3.3 1.1459999999999999e-05 3.3 1.156e-05 0 1.1479999999999999e-05 0 1.158e-05 3.3 1.1499999999999998e-05 3.3 1.1599999999999999e-05 0 1.152e-05 0 1.162e-05 3.3 1.154e-05 3.3 1.164e-05 0 1.156e-05 0 1.166e-05 3.3 1.158e-05 3.3 1.168e-05 0 1.1599999999999999e-05 0 1.17e-05 3.3 1.1619999999999999e-05 3.3 1.172e-05 0 1.1639999999999999e-05 0 1.174e-05 3.3 1.1659999999999998e-05 3.3 1.176e-05 0 1.1679999999999998e-05 0 1.1779999999999999e-05 3.3 1.17e-05 3.3 1.18e-05 0 1.172e-05 0 1.182e-05 3.3 1.174e-05 3.3 1.184e-05 0 1.176e-05 0 1.186e-05 3.3 1.1779999999999999e-05 3.3 1.188e-05 0 1.1799999999999999e-05 0 1.19e-05 3.3 1.1819999999999999e-05 3.3 1.192e-05 0 1.1839999999999998e-05 0 1.194e-05 3.3 1.1859999999999998e-05 3.3 1.1959999999999999e-05 0 1.188e-05 0 1.198e-05 3.3 1.19e-05 3.3 1.2e-05 0 1.192e-05 0 1.202e-05 3.3 1.194e-05 3.3 1.204e-05 0 1.1959999999999999e-05 0 1.206e-05 3.3 1.1979999999999999e-05 3.3 1.208e-05 0 1.1999999999999999e-05 0 1.21e-05 3.3 1.2019999999999998e-05 3.3 1.212e-05 0 1.2039999999999998e-05 0 1.2139999999999999e-05 3.3 1.206e-05 3.3 1.216e-05 0 1.208e-05 0 1.218e-05 3.3 1.21e-05 3.3 1.22e-05 0 1.212e-05 0 1.222e-05 3.3 1.2139999999999999e-05 3.3 1.224e-05 0 1.2159999999999999e-05 0 1.226e-05 3.3 1.2179999999999999e-05 3.3 1.228e-05 0 1.2199999999999998e-05 0 1.2299999999999999e-05 3.3 1.2219999999999998e-05 3.3 1.2319999999999999e-05 0 1.224e-05 0 1.234e-05 3.3 1.226e-05 3.3 1.236e-05 0 1.228e-05 0 1.238e-05 3.3 1.2299999999999999e-05 3.3 1.24e-05 0 1.2319999999999999e-05 0 1.242e-05 3.3 1.2339999999999999e-05 3.3 1.244e-05 0 1.2359999999999999e-05 0 1.246e-05 3.3 1.2379999999999998e-05 3.3 1.2479999999999999e-05 0 1.2399999999999998e-05 0 1.2499999999999999e-05 3.3 1.242e-05 3.3 1.252e-05 0 1.244e-05 0 1.254e-05 3.3 1.246e-05 3.3 1.256e-05 0 1.2479999999999999e-05 0 1.258e-05 3.3 1.2499999999999999e-05 3.3 1.26e-05 0 1.2519999999999999e-05 0 1.262e-05 3.3 1.2539999999999999e-05 3.3 1.264e-05 0 1.2559999999999998e-05 0 1.2659999999999999e-05 3.3 1.258e-05 3.3 1.268e-05 0 1.26e-05 0 1.27e-05 3.3 1.262e-05 3.3 1.272e-05 0 1.264e-05 0 1.274e-05 3.3 1.2659999999999999e-05 3.3 1.276e-05 0 1.2679999999999999e-05 0 1.278e-05 3.3 1.2699999999999999e-05 3.3 1.28e-05 0 1.2719999999999998e-05 0 1.282e-05 3.3 1.2739999999999998e-05 3.3 1.2839999999999999e-05 0 1.276e-05 0 1.286e-05 3.3 1.278e-05 3.3 1.288e-05 0 1.28e-05 0 1.29e-05 3.3 1.282e-05 3.3 1.292e-05 0 1.2839999999999999e-05 0 1.294e-05 3.3 1.2859999999999999e-05 3.3 1.296e-05 0 1.2879999999999999e-05 0 1.298e-05 3.3 1.2899999999999998e-05 3.3 1.3e-05 0 1.2919999999999998e-05 0 1.3019999999999999e-05 3.3 1.294e-05 3.3 1.304e-05 0 1.296e-05 0 1.306e-05 3.3 1.298e-05 3.3 1.308e-05 0 1.3e-05 0 1.31e-05 3.3 1.3019999999999999e-05 3.3 1.312e-05 0 1.3039999999999999e-05 0 1.314e-05 3.3 1.3059999999999999e-05 3.3 1.316e-05 0 1.3079999999999998e-05 0 1.318e-05 3.3 1.3099999999999998e-05 3.3 1.3199999999999999e-05 0 1.312e-05 0 1.322e-05 3.3 1.314e-05 3.3 1.324e-05 0 1.316e-05 0 1.326e-05 3.3 1.318e-05 3.3 1.328e-05 0 1.3199999999999999e-05 0 1.33e-05 3.3 1.3219999999999999e-05 3.3 1.332e-05 0 1.3239999999999999e-05 0 1.334e-05 3.3 1.3259999999999998e-05 3.3 1.3359999999999999e-05 0 1.3279999999999998e-05 0 1.3379999999999999e-05 3.3 1.33e-05 3.3 1.34e-05 0 1.332e-05 0 1.342e-05 3.3 1.334e-05 3.3 1.344e-05 0 1.3359999999999999e-05 0 1.346e-05 3.3 1.3379999999999999e-05 3.3 1.348e-05 0 1.3399999999999999e-05 0 1.35e-05 3.3 1.3419999999999999e-05 3.3 1.352e-05 0 1.3439999999999998e-05 0 1.3539999999999999e-05 3.3 1.3459999999999998e-05 3.3 1.3559999999999999e-05 0 1.348e-05 0 1.358e-05 3.3 1.35e-05 3.3 1.36e-05 0 1.352e-05 0 1.362e-05 3.3 1.3539999999999999e-05 3.3 1.364e-05 0 1.3559999999999999e-05 0 1.366e-05 3.3 1.3579999999999999e-05 3.3 1.368e-05 0 1.3599999999999999e-05 0 1.37e-05 3.3 1.3619999999999998e-05 3.3 1.3719999999999999e-05 0 1.3639999999999998e-05 0 1.3739999999999999e-05 3.3 1.366e-05 3.3 1.376e-05 0 1.368e-05 0 1.378e-05 3.3 1.37e-05 3.3 1.38e-05 0 1.3719999999999999e-05 0 1.382e-05 3.3 1.3739999999999999e-05 3.3 1.384e-05 0 1.3759999999999999e-05 0 1.386e-05 3.3 1.3779999999999999e-05 3.3 1.388e-05 0 1.3799999999999998e-05 0 1.3899999999999999e-05 3.3 1.382e-05 3.3 1.392e-05 0 1.384e-05 0 1.394e-05 3.3 1.386e-05 3.3 1.396e-05 0 1.388e-05 0 1.398e-05 3.3 1.3899999999999999e-05 3.3 1.4e-05 0 1.3919999999999999e-05 0 1.402e-05 3.3 1.3939999999999999e-05 3.3 1.404e-05 0 1.3959999999999998e-05 0 1.406e-05 3.3 1.3979999999999998e-05 3.3 1.4079999999999999e-05 0 1.4e-05 0 1.41e-05 3.3 1.402e-05 3.3 1.412e-05 0 1.404e-05 0 1.414e-05 3.3 1.406e-05 3.3 1.416e-05 0 1.4079999999999999e-05 0 1.418e-05 3.3 1.4099999999999999e-05 3.3 1.42e-05 0 1.4119999999999999e-05 0 1.422e-05 3.3 1.4139999999999998e-05 3.3 1.424e-05 0 1.4159999999999998e-05 0 1.4259999999999999e-05 3.3 1.418e-05 3.3 1.428e-05 0 1.42e-05 0 1.43e-05 3.3 1.422e-05 3.3 1.432e-05 0 1.424e-05 0 1.434e-05 3.3 1.4259999999999999e-05 3.3 1.436e-05 0 1.4279999999999999e-05 0 1.438e-05 3.3 1.4299999999999999e-05 3.3 1.44e-05 0 1.4319999999999998e-05 0 1.442e-05 3.3 1.4339999999999998e-05 3.3 1.4439999999999999e-05 0 1.436e-05 0 1.446e-05 3.3 1.438e-05 3.3 1.448e-05 0 1.44e-05 0 1.45e-05 3.3 1.442e-05 3.3 1.452e-05 0 1.4439999999999999e-05 0 1.454e-05 3.3 1.4459999999999999e-05 3.3 1.456e-05 0 1.4479999999999999e-05 0 1.458e-05 3.3 1.4499999999999998e-05 3.3 1.4599999999999999e-05 0 1.4519999999999998e-05 0 1.4619999999999999e-05 3.3 1.454e-05 3.3 1.464e-05 0 1.456e-05 0 1.466e-05 3.3 1.458e-05 3.3 1.468e-05 0 1.4599999999999999e-05 0 1.47e-05 3.3 1.4619999999999999e-05 3.3 1.472e-05 0 1.4639999999999999e-05 0 1.474e-05 3.3 1.4659999999999999e-05 3.3 1.476e-05 0 1.4679999999999998e-05 0 1.4779999999999999e-05 3.3 1.4699999999999998e-05 3.3 1.4799999999999999e-05 0 1.472e-05 0 1.482e-05 3.3 1.474e-05 3.3 1.484e-05 0 1.476e-05 0 1.486e-05 3.3 1.4779999999999999e-05 3.3 1.488e-05 0 1.4799999999999999e-05 0 1.49e-05 3.3 1.4819999999999999e-05 3.3 1.492e-05 0 1.4839999999999999e-05 0 1.494e-05 3.3 1.4859999999999998e-05 3.3 1.4959999999999999e-05 0 1.4879999999999998e-05 0 1.4979999999999999e-05 3.3 1.49e-05 3.3 1.5e-05 0 1.492e-05 0 1.502e-05 3.3 1.494e-05 3.3 1.504e-05 0 1.4959999999999999e-05 0 1.506e-05 3.3 1.4979999999999999e-05 3.3 1.508e-05 0 1.4999999999999999e-05 0 1.51e-05 3.3 1.5019999999999998e-05 3.3 1.512e-05 0 1.5039999999999998e-05 0 1.5139999999999999e-05 3.3 1.5059999999999998e-05 3.3 1.5159999999999999e-05 0 1.508e-05 0 1.518e-05 3.3 1.51e-05 3.3 1.52e-05 0 1.512e-05 0 1.522e-05 3.3 1.5139999999999999e-05 3.3 1.524e-05 0 1.5159999999999999e-05 0 1.526e-05 3.3 1.5179999999999999e-05 3.3 1.528e-05 0 1.5199999999999998e-05 0 1.53e-05 3.3 1.5219999999999998e-05 3.3 1.532e-05 0 1.5239999999999998e-05 0 1.534e-05 3.3 1.526e-05 3.3 1.536e-05 0 1.528e-05 0 1.538e-05 3.3 1.53e-05 3.3 1.5399999999999998e-05 0 1.532e-05 0 1.5419999999999998e-05 3.3 1.5340000000000002e-05 3.3 1.544e-05 0 1.5360000000000002e-05 0 1.546e-05 3.3 1.5380000000000002e-05 3.3 1.548e-05 0 1.54e-05 0 1.55e-05 3.3 1.542e-05 3.3 1.552e-05 0 1.544e-05 0 1.554e-05 3.3 1.546e-05 3.3 1.556e-05 0 1.548e-05 0 1.558e-05 3.3 1.55e-05 3.3 1.56e-05 0 1.552e-05 0 1.562e-05 3.3 1.554e-05 3.3 1.564e-05 0 1.556e-05 0 1.566e-05 3.3 1.558e-05 3.3 1.568e-05 0 1.56e-05 0 1.57e-05 3.3 1.562e-05 3.3 1.572e-05 0 1.564e-05 0 1.574e-05 3.3 1.566e-05 3.3 1.5759999999999998e-05 0 1.568e-05 0 1.5779999999999998e-05 3.3 1.5700000000000002e-05 3.3 1.58e-05 0 1.5720000000000002e-05 0 1.582e-05 3.3 1.5740000000000002e-05 3.3 1.584e-05 0 1.576e-05 0 1.586e-05 3.3 1.578e-05 3.3 1.588e-05 0 1.58e-05 0 1.59e-05 3.3 1.582e-05 3.3 1.592e-05 0 1.584e-05 0 1.594e-05 3.3 1.586e-05 3.3 1.596e-05 0 1.588e-05 0 1.598e-05 3.3 1.59e-05 3.3 1.6e-05 0 1.592e-05 0 1.602e-05 3.3 1.594e-05 3.3 1.604e-05 0 1.596e-05 0 1.606e-05 3.3 1.598e-05 3.3 1.608e-05 0 1.6e-05 0 1.61e-05 3.3 1.602e-05 3.3 1.6119999999999998e-05 0 1.6040000000000002e-05 0 1.614e-05 3.3 1.6060000000000002e-05 3.3 1.616e-05 0 1.6080000000000002e-05 0 1.618e-05 3.3 1.6100000000000002e-05 3.3 1.62e-05 0 1.612e-05 0 1.622e-05 3.3 1.614e-05 3.3 1.624e-05 0 1.616e-05 0 1.626e-05 3.3 1.618e-05 3.3 1.628e-05 0 1.62e-05 0 1.63e-05 3.3 1.622e-05 3.3 1.632e-05 0 1.624e-05 0 1.634e-05 3.3 1.626e-05 3.3 1.636e-05 0 1.628e-05 0 1.638e-05 3.3 1.63e-05 3.3 1.64e-05 0 1.632e-05 0 1.642e-05 3.3 1.634e-05 3.3 1.644e-05 0 1.636e-05 0 1.6459999999999998e-05 3.3 1.638e-05 3.3 1.6479999999999998e-05 0 1.6400000000000002e-05 0 1.65e-05 3.3 1.6420000000000002e-05 3.3 1.652e-05 0 1.6440000000000002e-05 0 1.654e-05 3.3 1.646e-05 3.3 1.656e-05 0 1.648e-05 0 1.658e-05 3.3 1.65e-05 3.3 1.66e-05 0 1.652e-05 0 1.662e-05 3.3 1.654e-05 3.3 1.664e-05 0 1.656e-05 0 1.666e-05 3.3 1.658e-05 3.3 1.668e-05 0 1.66e-05 0 1.67e-05 3.3 1.662e-05 3.3 1.672e-05 0 1.664e-05 0 1.674e-05 3.3 1.666e-05 3.3 1.676e-05 0 1.668e-05 0 1.678e-05 3.3 1.67e-05 3.3 1.68e-05 0 1.672e-05 0 1.6819999999999998e-05 3.3 1.674e-05 3.3 1.6839999999999998e-05 0 1.6760000000000002e-05 0 1.686e-05 3.3 1.6780000000000002e-05 3.3 1.688e-05 0 1.6800000000000002e-05 0 1.69e-05 3.3 1.682e-05 3.3 1.692e-05 0 1.684e-05 0 1.694e-05 3.3 1.686e-05 3.3 1.696e-05 0 1.688e-05 0 1.698e-05 3.3 1.69e-05 3.3 1.7e-05 0 1.692e-05 0 1.702e-05 3.3 1.694e-05 3.3 1.704e-05 0 1.696e-05 0 1.706e-05 3.3 1.698e-05 3.3 1.708e-05 0 1.7e-05 0 1.71e-05 3.3 1.702e-05 3.3 1.712e-05 0 1.704e-05 0 1.714e-05 3.3 1.706e-05 3.3 1.716e-05 0 1.708e-05 0 1.7179999999999998e-05 3.3 1.7100000000000002e-05 3.3 1.72e-05 0 1.7120000000000002e-05 0 1.722e-05 3.3 1.7140000000000002e-05 3.3 1.724e-05 0 1.7160000000000002e-05 0 1.726e-05 3.3 1.718e-05 3.3 1.728e-05 0 1.72e-05 0 1.73e-05 3.3 1.722e-05 3.3 1.732e-05 0 1.724e-05 0 1.734e-05 3.3 1.726e-05 3.3 1.736e-05 0 1.728e-05 0 1.738e-05 3.3 1.73e-05 3.3 1.74e-05 0 1.732e-05 0 1.742e-05 3.3 1.734e-05 3.3 1.744e-05 0 1.736e-05 0 1.746e-05 3.3 1.738e-05 3.3 1.748e-05 0 1.74e-05 0 1.75e-05 3.3 1.742e-05 3.3 1.7519999999999998e-05 0 1.744e-05 0 1.7539999999999998e-05 3.3 1.7460000000000002e-05 3.3 1.756e-05 0 1.7480000000000002e-05 0 1.758e-05 3.3 1.7500000000000002e-05 3.3 1.76e-05 0 1.752e-05 0 1.762e-05 3.3 1.754e-05 3.3 1.764e-05 0 1.756e-05 0 1.766e-05 3.3 1.758e-05 3.3 1.768e-05 0 1.76e-05 0 1.77e-05 3.3 1.762e-05 3.3 1.772e-05 0 1.764e-05 0 1.774e-05 3.3 1.766e-05 3.3 1.776e-05 0 1.768e-05 0 1.778e-05 3.3 1.77e-05 3.3 1.78e-05 0 1.772e-05 0 1.782e-05 3.3 1.774e-05 3.3 1.784e-05 0 1.776e-05 0 1.786e-05 3.3 1.778e-05 3.3 1.7879999999999998e-05 0 1.78e-05 0 1.7899999999999998e-05 3.3 1.7820000000000002e-05 3.3 1.792e-05 0 1.7840000000000002e-05 0 1.794e-05 3.3 1.7860000000000002e-05 3.3 1.796e-05 0 1.788e-05 0 1.798e-05 3.3 1.79e-05 3.3 1.8e-05 0 1.792e-05 0 1.802e-05 3.3 1.794e-05 3.3 1.804e-05 0 1.796e-05 0 1.806e-05 3.3 1.798e-05 3.3 1.808e-05 0 1.8e-05 0 1.81e-05 3.3 1.802e-05 3.3 1.812e-05 0 1.804e-05 0 1.814e-05 3.3 1.806e-05 3.3 1.816e-05 0 1.808e-05 0 1.818e-05 3.3 1.81e-05 3.3 1.82e-05 0 1.812e-05 0 1.822e-05 3.3 1.814e-05 3.3 1.8239999999999998e-05 0 1.816e-05 0 1.8259999999999998e-05 3.3 1.8180000000000002e-05 3.3 1.828e-05 0 1.8200000000000002e-05 0 1.83e-05 3.3 1.8220000000000002e-05 3.3 1.832e-05 0 1.824e-05 0 1.834e-05 3.3 1.826e-05 3.3 1.836e-05 0 1.828e-05 0 1.838e-05 3.3 1.83e-05 3.3 1.84e-05 0 1.832e-05 0 1.842e-05 3.3 1.834e-05 3.3 1.844e-05 0 1.836e-05 0 1.846e-05 3.3 1.838e-05 3.3 1.848e-05 0 1.84e-05 0 1.85e-05 3.3 1.842e-05 3.3 1.852e-05 0 1.844e-05 0 1.854e-05 3.3 1.846e-05 3.3 1.856e-05 0 1.848e-05 0 1.8579999999999998e-05 3.3 1.85e-05 3.3 1.8599999999999998e-05 0 1.8520000000000002e-05 0 1.862e-05 3.3 1.8540000000000002e-05 3.3 1.864e-05 0 1.8560000000000002e-05 0 1.866e-05 3.3 1.858e-05 3.3 1.868e-05 0 1.86e-05 0 1.87e-05 3.3 1.862e-05 3.3 1.872e-05 0 1.864e-05 0 1.874e-05 3.3 1.866e-05 3.3 1.876e-05 0 1.868e-05 0 1.878e-05 3.3 1.87e-05 3.3 1.88e-05 0 1.872e-05 0 1.882e-05 3.3 1.874e-05 3.3 1.884e-05 0 1.876e-05 0 1.886e-05 3.3 1.878e-05 3.3 1.888e-05 0 1.88e-05 0 1.89e-05 3.3 1.882e-05 3.3 1.892e-05 0 1.884e-05 0 1.8939999999999998e-05 3.3 1.886e-05 3.3 1.8959999999999998e-05 0 1.8880000000000002e-05 0 1.898e-05 3.3 1.8900000000000002e-05 3.3 1.9e-05 0 1.8920000000000002e-05 0 1.902e-05 3.3 1.894e-05 3.3 1.904e-05 0 1.896e-05 0 1.906e-05 3.3 1.898e-05 3.3 1.908e-05 0 1.9e-05 0 1.91e-05 3.3 1.902e-05 3.3 1.912e-05 0 1.904e-05 0 1.914e-05 3.3 1.906e-05 3.3 1.916e-05 0 1.908e-05 0 1.918e-05 3.3 1.91e-05 3.3 1.92e-05 0 1.912e-05 0 1.922e-05 3.3 1.914e-05 3.3 1.924e-05 0 1.916e-05 0 1.926e-05 3.3 1.918e-05 3.3 1.928e-05 0 1.92e-05 0 1.9299999999999998e-05 3.3 1.922e-05 3.3 1.9319999999999998e-05 0 1.9240000000000002e-05 0 1.934e-05 3.3 1.9260000000000002e-05 3.3 1.936e-05 0 1.9280000000000002e-05 0 1.938e-05 3.3 1.93e-05 3.3 1.94e-05 0 1.932e-05 0 1.942e-05 3.3 1.934e-05 3.3 1.944e-05 0 1.936e-05 0 1.946e-05 3.3 1.938e-05 3.3 1.948e-05 0 1.94e-05 0 1.95e-05 3.3 1.942e-05 3.3 1.952e-05 0 1.944e-05 0 1.954e-05 3.3 1.946e-05 3.3 1.956e-05 0 1.948e-05 0 1.958e-05 3.3 1.95e-05 3.3 1.96e-05 0 1.952e-05 0 1.962e-05 3.3 1.954e-05 3.3 1.964e-05 0 1.956e-05 0 1.9659999999999998e-05 3.3 1.958e-05 3.3 1.9679999999999998e-05 0 1.9600000000000002e-05 0 1.97e-05 3.3 1.9620000000000002e-05 3.3 1.972e-05 0 1.9640000000000002e-05 0 1.974e-05 3.3 1.966e-05 3.3 1.976e-05 0 1.968e-05 0 1.978e-05 3.3 1.97e-05 3.3 1.98e-05 0 1.972e-05 0 1.982e-05 3.3 1.974e-05 3.3 1.984e-05 0 1.976e-05 0 1.986e-05 3.3 1.978e-05 3.3 1.988e-05 0 1.98e-05 0 1.99e-05 3.3 1.982e-05 3.3 1.992e-05 0 1.984e-05 0 1.994e-05 3.3 1.986e-05 3.3 1.996e-05 0 1.988e-05 0 1.998e-05 3.3 1.99e-05 3.3 1.9999999999999998e-05 0 1.992e-05 0 2.0019999999999998e-05 3.3 1.9940000000000002e-05 3.3 2.004e-05 0 1.9960000000000002e-05 0 2.006e-05 3.3 1.9980000000000002e-05 3.3 2.008e-05 0 2e-05 0 2.01e-05 3.3 2.002e-05 3.3 2.012e-05 0 2.004e-05 0 2.014e-05 3.3 2.006e-05 3.3 2.016e-05 0 2.008e-05 0 2.018e-05 3.3 2.01e-05 3.3 2.02e-05 0 2.012e-05 0 2.022e-05 3.3 2.014e-05 3.3 2.024e-05 0 2.016e-05 0 2.026e-05 3.3 2.018e-05 3.3 2.028e-05 0 2.02e-05 0 2.03e-05 3.3 2.022e-05 3.3 2.032e-05 0 2.024e-05 0 2.034e-05 3.3 2.026e-05 3.3 2.0359999999999998e-05 0 2.028e-05 0 2.0379999999999998e-05 3.3 2.0300000000000002e-05 3.3 2.04e-05 0 2.0320000000000002e-05 0 2.042e-05 3.3 2.0340000000000002e-05 3.3 2.044e-05 0 2.036e-05 0 2.046e-05 3.3 2.038e-05 3.3 2.048e-05 0 2.04e-05 0 2.05e-05 3.3 2.042e-05 3.3 2.052e-05 0 2.044e-05 0 2.054e-05 3.3 2.046e-05 3.3 2.056e-05 0 2.048e-05 0 2.058e-05 3.3 2.05e-05 3.3 2.06e-05 0 2.052e-05 0 2.062e-05 3.3 2.054e-05 3.3 2.064e-05 0 2.056e-05 0 2.066e-05 3.3 2.058e-05 3.3 2.068e-05 0 2.06e-05 0 2.07e-05 3.3 2.062e-05 3.3 2.0719999999999998e-05 0 2.064e-05 0 2.0739999999999998e-05 3.3 2.0660000000000002e-05 3.3 2.076e-05 0 2.0680000000000002e-05 0 2.078e-05 3.3 2.0700000000000002e-05 3.3 2.08e-05 0 2.072e-05 0 2.082e-05 3.3 2.074e-05 3.3 2.084e-05 0 2.076e-05 0 2.086e-05 3.3 2.078e-05 3.3 2.088e-05 0 2.08e-05 0 2.09e-05 3.3 2.082e-05 3.3 2.092e-05 0 2.084e-05 0 2.094e-05 3.3 2.086e-05 3.3 2.096e-05 0 2.088e-05 0 2.098e-05 3.3 2.09e-05 3.3 2.1e-05 0 2.092e-05 0 2.102e-05 3.3 2.094e-05 3.3 2.104e-05 0 2.096e-05 0 2.1059999999999998e-05 3.3 2.098e-05 3.3 2.1079999999999998e-05 0 2.1000000000000002e-05 0 2.11e-05 3.3 2.1020000000000002e-05 3.3 2.112e-05 0 2.1040000000000002e-05 0 2.114e-05 3.3 2.106e-05 3.3 2.116e-05 0 2.108e-05 0 2.118e-05 3.3 2.11e-05 3.3 2.12e-05 0 2.112e-05 0 2.122e-05 3.3 2.114e-05 3.3 2.124e-05 0 2.116e-05 0 2.126e-05 3.3 2.118e-05 3.3 2.128e-05 0 2.12e-05 0 2.13e-05 3.3 2.122e-05 3.3 2.132e-05 0 2.124e-05 0 2.134e-05 3.3 2.126e-05 3.3 2.136e-05 0 2.128e-05 0 2.138e-05 3.3 2.13e-05 3.3 2.14e-05 0 2.132e-05 0 2.1419999999999998e-05 3.3 2.134e-05 3.3 2.1439999999999998e-05 0 2.1360000000000002e-05 0 2.146e-05 3.3 2.1380000000000002e-05 3.3 2.148e-05 0 2.1400000000000002e-05 0 2.15e-05 3.3 2.142e-05 3.3 2.152e-05 0 2.144e-05 0 2.154e-05 3.3 2.146e-05 3.3 2.156e-05 0 2.148e-05 0 2.158e-05 3.3 2.15e-05 3.3 2.16e-05 0 2.152e-05 0 2.162e-05 3.3 2.154e-05 3.3 2.164e-05 0 2.156e-05 0 2.166e-05 3.3 2.158e-05 3.3 2.168e-05 0 2.16e-05 0 2.17e-05 3.3 2.162e-05 3.3 2.172e-05 0 2.164e-05 0 2.174e-05 3.3 2.166e-05 3.3 2.176e-05 0 2.168e-05 0 2.1779999999999998e-05 3.3 2.17e-05 3.3 2.1799999999999998e-05 0 2.1720000000000002e-05 0 2.182e-05 3.3 2.1740000000000002e-05 3.3 2.184e-05 0 2.1760000000000002e-05 0 2.186e-05 3.3 2.178e-05 3.3 2.188e-05 0 2.18e-05 0 2.19e-05 3.3 2.182e-05 3.3 2.192e-05 0 2.184e-05 0 2.194e-05 3.3 2.186e-05 3.3 2.196e-05 0 2.188e-05 0 2.198e-05 3.3 2.19e-05 3.3 2.2e-05 0 2.192e-05 0 2.202e-05 3.3 2.194e-05 3.3 2.204e-05 0 2.196e-05 0 2.206e-05 3.3 2.198e-05 3.3 2.208e-05 0 2.2e-05 0 2.21e-05 3.3 2.202e-05 3.3 2.2119999999999998e-05 0 2.204e-05 0 2.2139999999999998e-05 3.3 2.206e-05 3.3 2.2159999999999998e-05 0 2.2080000000000002e-05 0 2.218e-05 3.3 2.2100000000000002e-05 3.3 2.22e-05 0 2.212e-05 0 2.222e-05 3.3 2.214e-05 3.3 2.224e-05 0 2.216e-05 0 2.226e-05 3.3 2.218e-05 3.3 2.228e-05 0 2.22e-05 0 2.23e-05 3.3 2.222e-05 3.3 2.232e-05 0 2.224e-05 0 2.234e-05 3.3 2.226e-05 3.3 2.236e-05 0 2.228e-05 0 2.238e-05 3.3 2.23e-05 3.3 2.24e-05 0 2.232e-05 0 2.242e-05 3.3 2.234e-05 3.3 2.244e-05 0 2.236e-05 0 2.246e-05 3.3 2.238e-05 3.3 2.2479999999999998e-05 0 2.24e-05 0 2.2499999999999998e-05 3.3 2.2420000000000002e-05 3.3 2.252e-05 0 2.2440000000000002e-05 0 2.254e-05 3.3 2.2460000000000002e-05 3.3 2.256e-05 0 2.248e-05 0 2.258e-05 3.3 2.25e-05 3.3 2.26e-05 0 2.252e-05 0 2.262e-05 3.3 2.254e-05 3.3 2.264e-05 0 2.256e-05 0 2.266e-05 3.3 2.258e-05 3.3 2.268e-05 0 2.26e-05 0 2.27e-05 3.3 2.262e-05 3.3 2.272e-05 0 2.264e-05 0 2.274e-05 3.3 2.266e-05 3.3 2.276e-05 0 2.268e-05 0 2.278e-05 3.3 2.27e-05 3.3 2.28e-05 0 2.272e-05 0 2.282e-05 3.3 2.274e-05 3.3 2.2839999999999998e-05 0 2.276e-05 0 2.2859999999999998e-05 3.3 2.2780000000000002e-05 3.3 2.288e-05 0 2.2800000000000002e-05 0 2.29e-05 3.3 2.2820000000000002e-05 3.3 2.292e-05 0 2.284e-05 0 2.294e-05 3.3 2.286e-05 3.3 2.296e-05 0 2.288e-05 0 2.298e-05 3.3 2.29e-05 3.3 2.3e-05 0 2.292e-05 0 2.302e-05 3.3 2.294e-05 3.3 2.304e-05 0 2.296e-05 0 2.306e-05 3.3 2.298e-05 3.3 2.308e-05 0 2.3e-05 0 2.31e-05 3.3 2.302e-05 3.3 2.312e-05 0 2.304e-05 0 2.314e-05 3.3 2.306e-05 3.3 2.316e-05 0 2.308e-05 0 2.3179999999999998e-05 3.3 2.31e-05 3.3 2.3199999999999998e-05 0 2.312e-05 0 2.3219999999999998e-05 3.3 2.3140000000000002e-05 3.3 2.324e-05 0 2.3160000000000002e-05 0 2.326e-05 3.3 2.318e-05 3.3 2.328e-05 0 2.32e-05 0 2.33e-05 3.3 2.322e-05 3.3 2.332e-05 0 2.324e-05 0 2.334e-05 3.3 2.326e-05 3.3 2.336e-05 0 2.328e-05 0 2.338e-05 3.3 2.33e-05 3.3 2.34e-05 0 2.332e-05 0 2.342e-05 3.3 2.334e-05 3.3 2.344e-05 0 2.336e-05 0 2.346e-05 3.3 2.338e-05 3.3 2.348e-05 0 2.34e-05 0 2.35e-05 3.3 2.342e-05 3.3 2.352e-05 0 2.344e-05 0 2.3539999999999998e-05 3.3 2.346e-05 3.3 2.3559999999999998e-05 0 2.348e-05 0 2.3579999999999998e-05 3.3 2.3500000000000002e-05 3.3 2.36e-05 0 2.3520000000000002e-05 0 2.362e-05 3.3 2.354e-05 3.3 2.364e-05 0 2.356e-05 0 2.366e-05 3.3 2.358e-05 3.3 2.368e-05 0 2.36e-05 0 2.37e-05 3.3 2.362e-05 3.3 2.372e-05 0 2.364e-05 0 2.374e-05 3.3 2.366e-05 3.3 2.376e-05 0 2.368e-05 0 2.378e-05 3.3 2.37e-05 3.3 2.38e-05 0 2.372e-05 0 2.382e-05 3.3 2.374e-05 3.3 2.384e-05 0 2.376e-05 0 2.386e-05 3.3 2.378e-05 3.3 2.388e-05 0 2.38e-05 0 2.3899999999999998e-05 3.3 2.382e-05 3.3 2.3919999999999998e-05 0 2.3840000000000002e-05 0 2.394e-05 3.3 2.3860000000000002e-05 3.3 2.396e-05 0 2.3880000000000002e-05 0 2.398e-05 3.3 2.39e-05 3.3 2.4e-05 0 2.392e-05 0 2.402e-05 3.3 2.394e-05 3.3 2.404e-05 0 2.396e-05 0 2.406e-05 3.3 2.398e-05 3.3 2.408e-05 0 2.4e-05 0 2.41e-05 3.3 2.402e-05 3.3 2.412e-05 0 2.404e-05 0 2.414e-05 3.3 2.406e-05 3.3 2.416e-05 0 2.408e-05 0 2.418e-05 3.3 2.41e-05 3.3 2.42e-05 0 2.412e-05 0 2.422e-05 3.3 2.414e-05 3.3 2.424e-05 0 2.416e-05 0 2.4259999999999998e-05 3.3 2.418e-05 3.3 2.4279999999999998e-05 0 2.4200000000000002e-05 0 2.43e-05 3.3 2.4220000000000002e-05 3.3 2.432e-05 0 2.4240000000000002e-05 0 2.434e-05 3.3 2.426e-05 3.3 2.436e-05 0 2.428e-05 0 2.438e-05 3.3 2.43e-05 3.3 2.44e-05 0 2.432e-05 0 2.442e-05 3.3 2.434e-05 3.3 2.444e-05 0 2.436e-05 0 2.446e-05 3.3 2.438e-05 3.3 2.448e-05 0 2.44e-05 0 2.45e-05 3.3 2.442e-05 3.3 2.452e-05 0 2.444e-05 0 2.454e-05 3.3 2.446e-05 3.3 2.456e-05 0 2.448e-05 0 2.458e-05 3.3 2.45e-05 3.3 2.4599999999999998e-05 0 2.452e-05 0 2.4619999999999998e-05 3.3 2.454e-05 3.3 2.4639999999999998e-05 0 2.4560000000000002e-05 0 2.466e-05 3.3 2.4580000000000002e-05 3.3 2.468e-05 0 2.46e-05 0 2.47e-05 3.3 2.462e-05 3.3 2.472e-05 0 2.464e-05 0 2.474e-05 3.3 2.466e-05 3.3 2.476e-05 0 2.468e-05 0 2.478e-05 3.3 2.47e-05 3.3 2.48e-05 0 2.472e-05 0 2.482e-05 3.3 2.474e-05 3.3 2.484e-05 0 2.476e-05 0 2.486e-05 3.3 2.478e-05 3.3 2.488e-05 0 2.48e-05 0 2.49e-05 3.3 2.482e-05 3.3 2.492e-05 0 2.484e-05 0 2.494e-05 3.3 2.486e-05 3.3 2.4959999999999998e-05 0 2.488e-05 0 2.4979999999999998e-05 3.3 2.49e-05 3.3 2.4999999999999998e-05 0 2.4920000000000002e-05 0 2.502e-05 3.3 2.4940000000000002e-05 3.3 2.504e-05 0 2.496e-05 0 2.506e-05 3.3 2.498e-05 3.3 2.508e-05 0 2.5e-05 0 2.51e-05 3.3 2.502e-05 3.3 2.512e-05 0 2.504e-05 0 2.514e-05 3.3 2.506e-05 3.3 2.516e-05 0 2.508e-05 0 2.518e-05 3.3 2.51e-05 3.3 2.52e-05 0 2.512e-05 0 2.522e-05 3.3 2.514e-05 3.3 2.524e-05 0 2.516e-05 0 2.526e-05 3.3 2.518e-05 3.3 2.528e-05 0 2.52e-05 0 2.53e-05 3.3 2.522e-05 3.3 2.5319999999999998e-05 0 2.524e-05 0 2.5339999999999998e-05 3.3 2.5260000000000002e-05 3.3 2.536e-05 0 2.5280000000000002e-05 0 2.538e-05 3.3 2.5300000000000002e-05 3.3 2.54e-05 0 2.532e-05 0 2.542e-05 3.3 2.534e-05 3.3 2.544e-05 0 2.536e-05 0 2.546e-05 3.3 2.538e-05 3.3 2.548e-05 0 2.54e-05 0 2.55e-05 3.3 2.542e-05 3.3 2.552e-05 0 2.544e-05 0 2.554e-05 3.3 2.546e-05 3.3 2.556e-05 0 2.548e-05 0 2.558e-05 3.3 2.55e-05 3.3 2.56e-05 0 2.552e-05 0 2.562e-05 3.3 2.554e-05 3.3 2.564e-05 0 2.556e-05 0 2.5659999999999998e-05 3.3 2.558e-05 3.3 2.5679999999999998e-05 0 2.56e-05 0 2.5699999999999998e-05 3.3 2.5620000000000002e-05 3.3 2.572e-05 0 2.5640000000000002e-05 0 2.574e-05 3.3 2.566e-05 3.3 2.576e-05 0 2.568e-05 0 2.578e-05 3.3 2.57e-05 3.3 2.58e-05 0 2.572e-05 0 2.582e-05 3.3 2.574e-05 3.3 2.584e-05 0 2.576e-05 0 2.586e-05 3.3 2.578e-05 3.3 2.588e-05 0 2.58e-05 0 2.59e-05 3.3 2.582e-05 3.3 2.592e-05 0 2.584e-05 0 2.594e-05 3.3 2.586e-05 3.3 2.596e-05 0 2.588e-05 0 2.598e-05 3.3 2.59e-05 3.3 2.6e-05 0 2.592e-05 0 2.6019999999999998e-05 3.3 2.594e-05 3.3 2.6039999999999998e-05 0 2.596e-05 0 2.6059999999999998e-05 3.3 2.5980000000000002e-05 3.3 2.608e-05 0 2.6000000000000002e-05 0 2.61e-05 3.3 2.602e-05 3.3 2.612e-05 0 2.604e-05 0 2.614e-05 3.3 2.606e-05 3.3 2.616e-05 0 2.608e-05 0 2.618e-05 3.3 2.61e-05 3.3 2.62e-05 0 2.612e-05 0 2.622e-05 3.3 2.614e-05 3.3 2.624e-05 0 2.616e-05 0 2.626e-05 3.3 2.618e-05 3.3 2.628e-05 0 2.62e-05 0 2.63e-05 3.3 2.622e-05 3.3 2.632e-05 0 2.624e-05 0 2.634e-05 3.3 2.626e-05 3.3 2.636e-05 0 2.628e-05 0 2.6379999999999998e-05 3.3 2.63e-05 3.3 2.6399999999999998e-05 0 2.6320000000000002e-05 0 2.642e-05 3.3 2.6340000000000002e-05 3.3 2.644e-05 0 2.6360000000000002e-05 0 2.646e-05 3.3 2.638e-05 3.3 2.648e-05 0 2.64e-05 0 2.65e-05 3.3 2.642e-05 3.3 2.652e-05 0 2.644e-05 0 2.654e-05 3.3 2.646e-05 3.3 2.656e-05 0 2.648e-05 0 2.658e-05 3.3 2.65e-05 3.3 2.66e-05 0 2.652e-05 0 2.662e-05 3.3 2.654e-05 3.3 2.664e-05 0 2.656e-05 0 2.666e-05 3.3 2.658e-05 3.3 2.668e-05 0 2.66e-05 0 2.67e-05 3.3 2.662e-05 3.3 2.6719999999999998e-05 0 2.664e-05 0 2.6739999999999998e-05 3.3 2.666e-05 3.3 2.6759999999999998e-05 0 2.6680000000000002e-05 0 2.678e-05 3.3 2.6700000000000002e-05 3.3 2.68e-05 0 2.672e-05 0 2.682e-05 3.3 2.674e-05 3.3 2.684e-05 0 2.676e-05 0 2.686e-05 3.3 2.678e-05 3.3 2.688e-05 0 2.68e-05 0 2.69e-05 3.3 2.682e-05 3.3 2.692e-05 0 2.684e-05 0 2.694e-05 3.3 2.686e-05 3.3 2.696e-05 0 2.688e-05 0 2.698e-05 3.3 2.69e-05 3.3 2.7e-05 0 2.692e-05 0 2.702e-05 3.3 2.694e-05 3.3 2.704e-05 0 2.696e-05 0 2.706e-05 3.3 2.698e-05 3.3 2.7079999999999998e-05 0 2.7e-05 0 2.7099999999999998e-05 3.3 2.702e-05 3.3 2.7119999999999998e-05 0 2.7040000000000002e-05 0 2.714e-05 3.3 2.7060000000000002e-05 3.3 2.716e-05 0 2.708e-05 0 2.718e-05 3.3 2.71e-05 3.3 2.72e-05 0 2.712e-05 0 2.722e-05 3.3 2.714e-05 3.3 2.724e-05 0 2.716e-05 0 2.726e-05 3.3 2.718e-05 3.3 2.728e-05 0 2.72e-05 0 2.73e-05 3.3 2.722e-05 3.3 2.732e-05 0 2.724e-05 0 2.734e-05 3.3 2.726e-05 3.3 2.736e-05 0 2.728e-05 0 2.738e-05 3.3 2.73e-05 3.3 2.74e-05 0 2.732e-05 0 2.742e-05 3.3 2.734e-05 3.3 2.7439999999999998e-05 0 2.736e-05 0 2.7459999999999998e-05 3.3 2.738e-05 3.3 2.7479999999999998e-05 0 2.7400000000000002e-05 0 2.75e-05 3.3 2.7420000000000002e-05 3.3 2.752e-05 0 2.744e-05 0 2.754e-05 3.3 2.746e-05 3.3 2.756e-05 0 2.748e-05 0 2.758e-05 3.3 2.75e-05 3.3 2.76e-05 0 2.752e-05 0 2.762e-05 3.3 2.754e-05 3.3 2.764e-05 0 2.756e-05 0 2.766e-05 3.3 2.758e-05 3.3 2.768e-05 0 2.76e-05 0 2.77e-05 3.3 2.762e-05 3.3 2.772e-05 0 2.764e-05 0 2.774e-05 3.3 2.766e-05 3.3 2.776e-05 0 2.768e-05 0 2.7779999999999998e-05 3.3 2.77e-05 3.3 2.7799999999999998e-05 0 2.772e-05 0 2.7819999999999998e-05 3.3 2.7740000000000002e-05 3.3 2.784e-05 0 2.7760000000000002e-05 0 2.786e-05 3.3 2.778e-05 3.3 2.788e-05 0 2.78e-05 0 2.79e-05 3.3 2.782e-05 3.3 2.792e-05 0 2.784e-05 0 2.794e-05 3.3 2.786e-05 3.3 2.796e-05 0 2.788e-05 0 2.798e-05 3.3 2.79e-05 3.3 2.8e-05 0 2.792e-05 0 2.802e-05 3.3 2.794e-05 3.3 2.804e-05 0 2.796e-05 0 2.806e-05 3.3 2.798e-05 3.3 2.808e-05 0 2.8e-05 0 2.81e-05 3.3 2.802e-05 3.3 2.812e-05 0 2.804e-05 0 2.8139999999999998e-05 3.3 2.806e-05 3.3 2.8159999999999998e-05 0 2.808e-05 0 2.8179999999999998e-05 3.3 2.8100000000000002e-05 3.3 2.82e-05 0 2.8120000000000002e-05 0 2.822e-05 3.3 2.814e-05 3.3 2.824e-05 0 2.816e-05 0 2.826e-05 3.3 2.818e-05 3.3 2.828e-05 0 2.82e-05 0 2.83e-05 3.3 2.822e-05 3.3 2.832e-05 0 2.824e-05 0 2.834e-05 3.3 2.826e-05 3.3 2.836e-05 0 2.828e-05 0 2.838e-05 3.3 2.83e-05 3.3 2.84e-05 0 2.832e-05 0 2.842e-05 3.3 2.834e-05 3.3 2.844e-05 0 2.836e-05 0 2.846e-05 3.3 2.838e-05 3.3 2.848e-05 0 2.84e-05 0 2.8499999999999998e-05 3.3 2.842e-05 3.3 2.8519999999999998e-05 0 2.844e-05 0 2.8539999999999998e-05 3.3 2.8460000000000002e-05 3.3 2.856e-05 0 2.8480000000000002e-05 0 2.858e-05 3.3 2.85e-05 3.3 2.86e-05 0 2.852e-05 0 2.862e-05 3.3 2.854e-05 3.3 2.864e-05 0 2.856e-05 0 2.866e-05 3.3 2.858e-05 3.3 2.868e-05 0 2.86e-05 0 2.87e-05 3.3 2.862e-05 3.3 2.872e-05 0 2.864e-05 0 2.874e-05 3.3 2.866e-05 3.3 2.876e-05 0 2.868e-05 0 2.878e-05 3.3 2.87e-05 3.3 2.88e-05 0 2.872e-05 0 2.882e-05 3.3 2.874e-05 3.3 2.884e-05 0 2.876e-05 0 2.8859999999999998e-05 3.3 2.878e-05 3.3 2.8879999999999998e-05 0 2.88e-05 0 2.8899999999999998e-05 3.3 2.8820000000000002e-05 3.3 2.892e-05 0 2.8840000000000002e-05 0 2.894e-05 3.3 2.886e-05 3.3 2.896e-05 0 2.888e-05 0 2.898e-05 3.3 2.89e-05 3.3 2.9e-05 0 2.892e-05 0 2.902e-05 3.3 2.894e-05 3.3 2.904e-05 0 2.896e-05 0 2.906e-05 3.3 2.898e-05 3.3 2.908e-05 0 2.9e-05 0 2.91e-05 3.3 2.902e-05 3.3 2.912e-05 0 2.904e-05 0 2.914e-05 3.3 2.906e-05 3.3 2.916e-05 0 2.908e-05 0 2.918e-05 3.3 2.91e-05 3.3 2.9199999999999998e-05 0 2.912e-05 0 2.9219999999999998e-05 3.3 2.914e-05 3.3 2.9239999999999998e-05 0 2.9160000000000002e-05 0 2.926e-05 3.3 2.9180000000000002e-05 3.3 2.928e-05 0 2.92e-05 0 2.93e-05 3.3 2.922e-05 3.3 2.932e-05 0 2.924e-05 0 2.934e-05 3.3 2.926e-05 3.3 2.936e-05 0 2.928e-05 0 2.938e-05 3.3 2.93e-05 3.3 2.94e-05 0 2.932e-05 0 2.942e-05 3.3 2.934e-05 3.3 2.944e-05 0 2.936e-05 0 2.946e-05 3.3 2.938e-05 3.3 2.948e-05 0 2.94e-05 0 2.95e-05 3.3 2.942e-05 3.3 2.952e-05 0 2.944e-05 0 2.954e-05 3.3 2.946e-05 3.3 2.9559999999999998e-05 0 2.948e-05 0 2.9579999999999998e-05 3.3 2.95e-05 3.3 2.9599999999999998e-05 0 2.9520000000000002e-05 0 2.962e-05 3.3 2.9540000000000002e-05 3.3 2.964e-05 0 2.956e-05 0 2.966e-05 3.3 2.958e-05 3.3 2.968e-05 0 2.96e-05 0 2.97e-05 3.3 2.962e-05 3.3 2.972e-05 0 2.964e-05 0 2.974e-05 3.3 2.966e-05 3.3 2.976e-05 0 2.968e-05 0 2.978e-05 3.3 2.97e-05 3.3 2.98e-05 0 2.972e-05 0 2.982e-05 3.3 2.974e-05 3.3 2.984e-05 0 2.976e-05 0 2.986e-05 3.3 2.978e-05 3.3 2.988e-05 0 2.98e-05 0 2.99e-05 3.3 2.982e-05 3.3 2.9919999999999998e-05 0 2.984e-05 0 2.9939999999999998e-05 3.3 2.986e-05 3.3 2.9959999999999998e-05 0 2.9880000000000002e-05 0 2.998e-05 3.3 2.9900000000000002e-05 3.3 3e-05 0 2.992e-05 0 3.002e-05 3.3 2.994e-05 3.3 3.004e-05 0 2.996e-05 0 3.006e-05 3.3 2.998e-05 3.3 3.008e-05 0 3e-05 0 3.01e-05 3.3 3.002e-05 3.3 3.012e-05 0 3.004e-05 0 3.014e-05 3.3 3.006e-05 3.3 3.016e-05 0 3.008e-05 0 3.018e-05 3.3 3.01e-05 3.3 3.02e-05 0 3.012e-05 0 3.022e-05 3.3 3.014e-05 3.3 3.024e-05 0 3.016e-05 0 3.0259999999999998e-05 3.3 3.018e-05 3.3 3.0279999999999998e-05 0 3.02e-05 0 3.0299999999999998e-05 3.3 3.022e-05 3.3 3.0319999999999998e-05 0 3.0240000000000002e-05 0 3.034e-05 3.3 3.026e-05 3.3 3.036e-05 0 3.028e-05 0 3.038e-05 3.3 3.03e-05 3.3 3.04e-05 0 3.032e-05 0 3.042e-05 3.3 3.034e-05 3.3 3.044e-05 0 3.036e-05 0 3.046e-05 3.3 3.038e-05 3.3 3.048e-05 0 3.04e-05 0 3.05e-05 3.3 3.042e-05 3.3 3.052e-05 0 3.0440000000000003e-05 0 3.054e-05 3.3 3.046e-05 3.3 3.056e-05 0 3.0480000000000003e-05 0 3.058e-05 3.3 3.05e-05 3.3 3.06e-05 0 3.052e-05 0 3.062e-05 3.3 3.0539999999999996e-05 3.3 3.064e-05 0 3.056e-05 0 3.066e-05 3.3 3.0579999999999995e-05 3.3 3.068e-05 0 3.06e-05 0 3.07e-05 3.3 3.0619999999999995e-05 3.3 3.072e-05 0 3.064e-05 0 3.074e-05 3.3 3.0659999999999994e-05 3.3 3.076e-05 0 3.068e-05 0 3.078e-05 3.3 3.0699999999999994e-05 3.3 3.0799999999999996e-05 0 3.072e-05 0 3.082e-05 3.3 3.0739999999999994e-05 3.3 3.0839999999999996e-05 0 3.076e-05 0 3.086e-05 3.3 3.078e-05 3.3 3.088e-05 0 3.0799999999999996e-05 0 3.09e-05 3.3 3.082e-05 3.3 3.092e-05 0 3.0839999999999996e-05 0 3.094e-05 3.3 3.086e-05 3.3 3.096e-05 0 3.0879999999999996e-05 0 3.098e-05 3.3 3.09e-05 3.3 3.1e-05 0 3.0919999999999995e-05 0 3.102e-05 3.3 3.094e-05 3.3 3.104e-05 0 3.0959999999999995e-05 0 3.106e-05 3.3 3.098e-05 3.3 3.108e-05 0 3.0999999999999995e-05 0 3.11e-05 3.3 3.102e-05 3.3 3.112e-05 0 3.1039999999999994e-05 0 3.114e-05 3.3 3.106e-05 3.3 3.116e-05 0 3.1079999999999994e-05 0 3.1179999999999996e-05 3.3 3.11e-05 3.3 3.12e-05 0 3.112e-05 0 3.122e-05 3.3 3.114e-05 3.3 3.124e-05 0 3.116e-05 0 3.126e-05 3.3 3.1179999999999996e-05 3.3 3.128e-05 0 3.12e-05 0 3.13e-05 3.3 3.1219999999999996e-05 3.3 3.132e-05 0 3.124e-05 0 3.134e-05 3.3 3.1259999999999995e-05 3.3 3.136e-05 0 3.128e-05 0 3.138e-05 3.3 3.1299999999999995e-05 3.3 3.14e-05 0 3.132e-05 0 3.142e-05 3.3 3.1339999999999995e-05 3.3 3.144e-05 0 3.136e-05 0 3.146e-05 3.3 3.1379999999999994e-05 3.3 3.148e-05 0 3.14e-05 0 3.15e-05 3.3 3.1419999999999994e-05 3.3 3.1519999999999996e-05 0 3.144e-05 0 3.154e-05 3.3 3.1459999999999994e-05 3.3 3.1559999999999996e-05 0 3.148e-05 0 3.158e-05 3.3 3.15e-05 3.3 3.16e-05 0 3.1519999999999996e-05 0 3.162e-05 3.3 3.154e-05 3.3 3.164e-05 0 3.1559999999999996e-05 0 3.166e-05 3.3 3.158e-05 3.3 3.168e-05 0 3.1599999999999996e-05 0 3.17e-05 3.3 3.162e-05 3.3 3.172e-05 0 3.1639999999999995e-05 0 3.174e-05 3.3 3.166e-05 3.3 3.176e-05 0 3.1679999999999995e-05 0 3.178e-05 3.3 3.17e-05 3.3 3.18e-05 0 3.1719999999999994e-05 0 3.182e-05 3.3 3.174e-05 3.3 3.184e-05 0 3.1759999999999994e-05 0 3.1859999999999997e-05 3.3 3.178e-05 3.3 3.188e-05 0 3.1799999999999994e-05 0 3.1899999999999996e-05 3.3 3.182e-05 3.3 3.192e-05 0 3.184e-05 0 3.194e-05 3.3 3.1859999999999997e-05 3.3 3.196e-05 0 3.188e-05 0 3.198e-05 3.3 3.1899999999999996e-05 3.3 3.2e-05 0 3.192e-05 0 3.202e-05 3.3 3.1939999999999996e-05 3.3 3.204e-05 0 3.196e-05 0 3.206e-05 3.3 3.1979999999999995e-05 3.3 3.208e-05 0 3.2e-05 0 3.21e-05 3.3 3.2019999999999995e-05 3.3 3.212e-05 0 3.204e-05 0 3.214e-05 3.3 3.2059999999999995e-05 3.3 3.216e-05 0 3.208e-05 0 3.218e-05 3.3 3.2099999999999994e-05 3.3 3.22e-05 0 3.212e-05 0 3.222e-05 3.3 3.2139999999999994e-05 3.3 3.2239999999999996e-05 0 3.216e-05 0 3.226e-05 3.3 3.218e-05 3.3 3.228e-05 0 3.22e-05 0 3.23e-05 3.3 3.222e-05 3.3 3.232e-05 0 3.2239999999999996e-05 0 3.234e-05 3.3 3.226e-05 3.3 3.236e-05 0 3.2279999999999996e-05 0 3.238e-05 3.3 3.23e-05 3.3 3.24e-05 0 3.2319999999999995e-05 0 3.242e-05 3.3 3.234e-05 3.3 3.244e-05 0 3.2359999999999995e-05 0 3.246e-05 3.3 3.238e-05 3.3 3.248e-05 0 3.2399999999999995e-05 0 3.25e-05 3.3 3.242e-05 3.3 3.252e-05 0 3.2439999999999994e-05 0 3.254e-05 3.3 3.246e-05 3.3 3.256e-05 0 3.2479999999999994e-05 0 3.2579999999999996e-05 3.3 3.25e-05 3.3 3.26e-05 0 3.2519999999999994e-05 0 3.2619999999999996e-05 3.3 3.254e-05 3.3 3.264e-05 0 3.256e-05 0 3.266e-05 3.3 3.2579999999999996e-05 3.3 3.268e-05 0 3.26e-05 0 3.27e-05 3.3 3.2619999999999996e-05 3.3 3.272e-05 0 3.264e-05 0 3.274e-05 3.3 3.2659999999999996e-05 3.3 3.276e-05 0 3.268e-05 0 3.278e-05 3.3 3.2699999999999995e-05 3.3 3.28e-05 0 3.272e-05 0 3.282e-05 3.3 3.2739999999999995e-05 3.3 3.284e-05 0 3.276e-05 0 3.286e-05 3.3 3.2779999999999994e-05 3.3 3.288e-05 0 3.28e-05 0 3.29e-05 3.3 3.2819999999999994e-05 3.3 3.2919999999999997e-05 0 3.284e-05 0 3.294e-05 3.3 3.2859999999999994e-05 3.3 3.2959999999999996e-05 0 3.288e-05 0 3.298e-05 3.3 3.29e-05 3.3 3.3e-05 0 3.2919999999999997e-05 0 3.302e-05 3.3 3.294e-05 3.3 3.304e-05 0 3.2959999999999996e-05 0 3.306e-05 3.3 3.298e-05 3.3 3.308e-05 0 3.2999999999999996e-05 0 3.31e-05 3.3 3.302e-05 3.3 3.312e-05 0 3.3039999999999995e-05 0 3.314e-05 3.3 3.306e-05 3.3 3.316e-05 0 3.3079999999999995e-05 0 3.318e-05 3.3 3.31e-05 3.3 3.32e-05 0 3.3119999999999995e-05 0 3.322e-05 3.3 3.314e-05 3.3 3.324e-05 0 3.3159999999999994e-05 0 3.326e-05 3.3 3.318e-05 3.3 3.328e-05 0 3.3199999999999994e-05 0 3.3299999999999996e-05 3.3 3.322e-05 3.3 3.332e-05 0 3.324e-05 0 3.334e-05 3.3 3.326e-05 3.3 3.336e-05 0 3.328e-05 0 3.338e-05 3.3 3.3299999999999996e-05 3.3 3.34e-05 0 3.332e-05 0 3.342e-05 3.3 3.3339999999999996e-05 3.3 3.344e-05 0 3.336e-05 0 3.346e-05 3.3 3.3379999999999996e-05 3.3 3.348e-05 0 3.34e-05 0 3.35e-05 3.3 3.3419999999999995e-05 3.3 3.352e-05 0 3.344e-05 0 3.354e-05 3.3 3.3459999999999995e-05 3.3 3.356e-05 0 3.348e-05 0 3.358e-05 3.3 3.3499999999999994e-05 3.3 3.36e-05 0 3.352e-05 0 3.362e-05 3.3 3.3539999999999994e-05 3.3 3.3639999999999996e-05 0 3.356e-05 0 3.366e-05 3.3 3.3579999999999994e-05 3.3 3.3679999999999996e-05 0 3.36e-05 0 3.37e-05 3.3 3.362e-05 3.3 3.372e-05 0 3.3639999999999996e-05 0 3.374e-05 3.3 3.366e-05 3.3 3.376e-05 0 3.3679999999999996e-05 0 3.378e-05 3.3 3.37e-05 3.3 3.38e-05 0 3.3719999999999996e-05 0 3.382e-05 3.3 3.374e-05 3.3 3.384e-05 0 3.3759999999999995e-05 0 3.386e-05 3.3 3.378e-05 3.3 3.388e-05 0 3.3799999999999995e-05 0 3.39e-05 3.3 3.382e-05 3.3 3.392e-05 0 3.3839999999999994e-05 0 3.394e-05 3.3 3.386e-05 3.3 3.396e-05 0 3.3879999999999994e-05 0 3.3979999999999997e-05 3.3 3.39e-05 3.3 3.4e-05 0 3.3919999999999994e-05 0 3.4019999999999996e-05 3.3 3.394e-05 3.3 3.404e-05 0 3.396e-05 0 3.406e-05 3.3 3.3979999999999997e-05 3.3 3.408e-05 0 3.4e-05 0 3.41e-05 3.3 3.4019999999999996e-05 3.3 3.412e-05 0 3.404e-05 0 3.414e-05 3.3 3.4059999999999996e-05 3.3 3.416e-05 0 3.408e-05 0 3.418e-05 3.3 3.4099999999999995e-05 3.3 3.42e-05 0 3.412e-05 0 3.422e-05 3.3 3.4139999999999995e-05 3.3 3.424e-05 0 3.416e-05 0 3.426e-05 3.3 3.4179999999999995e-05 3.3 3.428e-05 0 3.42e-05 0 3.43e-05 3.3 3.4219999999999994e-05 3.3 3.432e-05 0 3.424e-05 0 3.434e-05 3.3 3.4259999999999994e-05 3.3 3.4359999999999996e-05 0 3.428e-05 0 3.438e-05 3.3 3.43e-05 3.3 3.44e-05 0 3.432e-05 0 3.442e-05 3.3 3.434e-05 3.3 3.444e-05 0 3.4359999999999996e-05 0 3.446e-05 3.3 3.438e-05 3.3 3.448e-05 0 3.4399999999999996e-05 0 3.45e-05 3.3 3.442e-05 3.3 3.452e-05 0 3.4439999999999996e-05 0 3.454e-05 3.3 3.446e-05 3.3 3.456e-05 0 3.4479999999999995e-05 0 3.458e-05 3.3 3.45e-05 3.3 3.46e-05 0 3.4519999999999995e-05 0 3.462e-05 3.3 3.454e-05 3.3 3.464e-05 0 3.4559999999999994e-05 0 3.466e-05 3.3 3.458e-05 3.3 3.468e-05 0 3.4599999999999994e-05 0 3.4699999999999996e-05 3.3 3.462e-05 3.3 3.472e-05 0 3.4639999999999994e-05 0 3.4739999999999996e-05 3.3 3.466e-05 3.3 3.476e-05 0 3.468e-05 0 3.478e-05 3.3 3.4699999999999996e-05 3.3 3.48e-05 0 3.472e-05 0 3.482e-05 3.3 3.4739999999999996e-05 3.3 3.484e-05 0 3.476e-05 0 3.486e-05 3.3 3.4779999999999996e-05 3.3 3.488e-05 0 3.48e-05 0 3.49e-05 3.3 3.4819999999999995e-05 3.3 3.492e-05 0 3.484e-05 0 3.494e-05 3.3 3.4859999999999995e-05 3.3 3.496e-05 0 3.488e-05 0 3.498e-05 3.3 3.4899999999999995e-05 3.3 3.5e-05 0 3.492e-05 0 3.502e-05 3.3 3.4939999999999994e-05 3.3 3.5039999999999997e-05 0 3.496e-05 0 3.506e-05 3.3 3.4979999999999994e-05 3.3 3.5079999999999996e-05 0 3.5e-05 0 3.51e-05 3.3 3.502e-05 3.3 3.512e-05 0 3.5039999999999997e-05 0 3.514e-05 3.3 3.506e-05 3.3 3.516e-05 0 3.5079999999999996e-05 0 3.518e-05 3.3 3.51e-05 3.3 3.52e-05 0 3.5119999999999996e-05 0 3.522e-05 3.3 3.514e-05 3.3 3.524e-05 0 3.5159999999999995e-05 0 3.526e-05 3.3 3.518e-05 3.3 3.528e-05 0 3.5199999999999995e-05 0 3.53e-05 3.3 3.522e-05 3.3 3.532e-05 0 3.5239999999999995e-05 0 3.534e-05 3.3 3.526e-05 3.3 3.536e-05 0 3.5279999999999994e-05 0 3.538e-05 3.3 3.53e-05 3.3 3.54e-05 0 3.5319999999999994e-05 0 3.5419999999999996e-05 3.3 3.534e-05 3.3 3.544e-05 0 3.5359999999999993e-05 0 3.5459999999999996e-05 3.3 3.538e-05 3.3 3.548e-05 0 3.54e-05 0 3.55e-05 3.3 3.5419999999999996e-05 3.3 3.552e-05 0 3.544e-05 0 3.554e-05 3.3 3.5459999999999996e-05 3.3 3.556e-05 0 3.548e-05 0 3.558e-05 3.3 3.5499999999999996e-05 3.3 3.56e-05 0 3.552e-05 0 3.562e-05 3.3 3.5539999999999995e-05 3.3 3.564e-05 0 3.556e-05 0 3.566e-05 3.3 3.5579999999999995e-05 3.3 3.568e-05 0 3.56e-05 0 3.57e-05 3.3 3.5619999999999994e-05 3.3 3.572e-05 0 3.564e-05 0 3.574e-05 3.3 3.5659999999999994e-05 3.3 3.5759999999999996e-05 0 3.568e-05 0 3.578e-05 3.3 3.5699999999999994e-05 3.3 3.5799999999999996e-05 0 3.572e-05 0 3.582e-05 3.3 3.574e-05 3.3 3.584e-05 0 3.5759999999999996e-05 0 3.586e-05 3.3 3.578e-05 3.3 3.588e-05 0 3.5799999999999996e-05 0 3.59e-05 3.3 3.582e-05 3.3 3.592e-05 0 3.5839999999999996e-05 0 3.594e-05 3.3 3.586e-05 3.3 3.596e-05 0 3.5879999999999995e-05 0 3.598e-05 3.3 3.59e-05 3.3 3.6e-05 0 3.5919999999999995e-05 0 3.602e-05 3.3 3.594e-05 3.3 3.604e-05 0 3.5959999999999995e-05 0 3.606e-05 3.3 3.598e-05 3.3 3.608e-05 0 3.5999999999999994e-05 0 3.6099999999999997e-05 3.3 3.602e-05 3.3 3.612e-05 0 3.6039999999999994e-05 0 3.6139999999999996e-05 3.3 3.606e-05 3.3 3.616e-05 0 3.608e-05 0 3.618e-05 3.3 3.6099999999999997e-05 3.3 3.62e-05 0 3.612e-05 0 3.622e-05 3.3 3.6139999999999996e-05 3.3 3.624e-05 0 3.616e-05 0 3.626e-05 3.3 3.6179999999999996e-05 3.3 3.628e-05 0 3.62e-05 0 3.63e-05 3.3 3.6219999999999995e-05 3.3 3.632e-05 0 3.624e-05 0 3.634e-05 3.3 3.6259999999999995e-05 3.3 3.636e-05 0 3.628e-05 0 3.638e-05 3.3 3.6299999999999995e-05 3.3 3.64e-05 0 3.632e-05 0 3.642e-05 3.3 3.6339999999999994e-05 3.3 3.644e-05 0 3.636e-05 0 3.646e-05 3.3 3.6379999999999994e-05 3.3 3.6479999999999996e-05 0 3.64e-05 0 3.65e-05 3.3 3.6419999999999994e-05 3.3 3.6519999999999996e-05 0 3.644e-05 0 3.654e-05 3.3 3.646e-05 3.3 3.656e-05 0 3.6479999999999996e-05 0 3.658e-05 3.3 3.65e-05 3.3 3.66e-05 0 3.6519999999999996e-05 0 3.662e-05 3.3 3.654e-05 3.3 3.664e-05 0 3.6559999999999996e-05 0 3.666e-05 3.3 3.658e-05 3.3 3.668e-05 0 3.6599999999999995e-05 0 3.67e-05 3.3 3.662e-05 3.3 3.672e-05 0 3.6639999999999995e-05 0 3.674e-05 3.3 3.666e-05 3.3 3.676e-05 0 3.6679999999999994e-05 0 3.678e-05 3.3 3.67e-05 3.3 3.68e-05 0 3.6719999999999994e-05 0 3.6819999999999996e-05 3.3 3.674e-05 3.3 3.684e-05 0 3.6759999999999994e-05 0 3.6859999999999996e-05 3.3 3.678e-05 3.3 3.688e-05 0 3.68e-05 0 3.69e-05 3.3 3.6819999999999996e-05 3.3 3.692e-05 0 3.684e-05 0 3.694e-05 3.3 3.6859999999999996e-05 3.3 3.696e-05 0 3.688e-05 0 3.698e-05 3.3 3.6899999999999996e-05 3.3 3.7e-05 0 3.692e-05 0 3.702e-05 3.3 3.6939999999999995e-05 3.3 3.704e-05 0 3.696e-05 0 3.706e-05 3.3 3.6979999999999995e-05 3.3 3.708e-05 0 3.7e-05 0 3.71e-05 3.3 3.7019999999999995e-05 3.3 3.712e-05 0 3.704e-05 0 3.714e-05 3.3 3.7059999999999994e-05 3.3 3.7159999999999997e-05 0 3.708e-05 0 3.718e-05 3.3 3.7099999999999994e-05 3.3 3.7199999999999996e-05 0 3.712e-05 0 3.722e-05 3.3 3.714e-05 3.3 3.724e-05 0 3.7159999999999997e-05 0 3.726e-05 3.3 3.718e-05 3.3 3.728e-05 0 3.7199999999999996e-05 0 3.73e-05 3.3 3.722e-05 3.3 3.732e-05 0 3.7239999999999996e-05 0 3.734e-05 3.3 3.726e-05 3.3 3.736e-05 0 3.7279999999999995e-05 0 3.738e-05 3.3 3.73e-05 3.3 3.74e-05 0 3.7319999999999995e-05 0 3.742e-05 3.3 3.734e-05 3.3 3.744e-05 0 3.7359999999999995e-05 0 3.746e-05 3.3 3.738e-05 3.3 3.748e-05 0 3.7399999999999994e-05 0 3.75e-05 3.3 3.742e-05 3.3 3.752e-05 0 3.7439999999999994e-05 0 3.7539999999999996e-05 3.3 3.746e-05 3.3 3.756e-05 0 3.7479999999999994e-05 0 3.7579999999999996e-05 3.3 3.75e-05 3.3 3.76e-05 0 3.752e-05 0 3.762e-05 3.3 3.7539999999999996e-05 3.3 3.764e-05 0 3.756e-05 0 3.766e-05 3.3 3.7579999999999996e-05 3.3 3.768e-05 0 3.76e-05 0 3.77e-05 3.3 3.7619999999999996e-05 3.3 3.772e-05 0 3.764e-05 0 3.774e-05 3.3 3.7659999999999995e-05 3.3 3.776e-05 0 3.768e-05 0 3.778e-05 3.3 3.7699999999999995e-05 3.3 3.78e-05 0 3.772e-05 0 3.782e-05 3.3 3.7739999999999994e-05 3.3 3.784e-05 0 3.776e-05 0 3.786e-05 3.3 3.7779999999999994e-05 3.3 3.7879999999999996e-05 0 3.78e-05 0 3.79e-05 3.3 3.7819999999999994e-05 3.3 3.7919999999999996e-05 0 3.784e-05 0 3.794e-05 3.3 3.786e-05 3.3 3.796e-05 0 3.7879999999999996e-05 0 3.798e-05 3.3 3.79e-05 3.3 3.8e-05 0 3.7919999999999996e-05 0 3.802e-05 3.3 3.794e-05 3.3 3.804e-05 0 3.7959999999999996e-05 0 3.806e-05 3.3 3.798e-05 3.3 3.808e-05 0 3.7999999999999995e-05 0 3.81e-05 3.3 3.802e-05 3.3 3.812e-05 0 3.8039999999999995e-05 0 3.814e-05 3.3 3.806e-05 3.3 3.816e-05 0 3.8079999999999995e-05 0 3.818e-05 3.3 3.81e-05 3.3 3.82e-05 0 3.8119999999999994e-05 0 3.8219999999999997e-05 3.3 3.814e-05 3.3 3.824e-05 0 3.8159999999999994e-05 0 3.8259999999999996e-05 3.3 3.818e-05 3.3 3.828e-05 0 3.82e-05 0 3.83e-05 3.3 3.8219999999999997e-05 3.3 3.832e-05 0 3.824e-05 0 3.834e-05 3.3 3.8259999999999996e-05 3.3 3.836e-05 0 3.828e-05 0 3.838e-05 3.3 3.8299999999999996e-05 3.3 3.84e-05 0 3.832e-05 0 3.842e-05 3.3 3.8339999999999995e-05 3.3 3.844e-05 0 3.836e-05 0 3.846e-05 3.3 3.8379999999999995e-05 3.3 3.848e-05 0 3.84e-05 0 3.85e-05 3.3 3.8419999999999995e-05 3.3 3.852e-05 0 3.844e-05 0 3.854e-05 3.3 3.8459999999999994e-05 3.3 3.856e-05 0 3.848e-05 0 3.858e-05 3.3 3.8499999999999994e-05 3.3 3.8599999999999996e-05 0 3.852e-05 0 3.862e-05 3.3 3.8539999999999994e-05 3.3 3.8639999999999996e-05 0 3.856e-05 0 3.866e-05 3.3 3.858e-05 3.3 3.868e-05 0 3.8599999999999996e-05 0 3.87e-05 3.3 3.862e-05 3.3 3.872e-05 0 3.8639999999999996e-05 0 3.874e-05 3.3 3.866e-05 3.3 3.876e-05 0 3.8679999999999996e-05 0 3.878e-05 3.3 3.87e-05 3.3 3.88e-05 0 3.8719999999999995e-05 0 3.882e-05 3.3 3.874e-05 3.3 3.884e-05 0 3.8759999999999995e-05 0 3.886e-05 3.3 3.878e-05 3.3 3.888e-05 0 3.8799999999999994e-05 0 3.89e-05 3.3 3.882e-05 3.3 3.892e-05 0 3.8839999999999994e-05 0 3.8939999999999996e-05 3.3 3.886e-05 3.3 3.896e-05 0 3.8879999999999994e-05 0 3.8979999999999996e-05 3.3 3.89e-05 3.3 3.9e-05 0 3.892e-05 0 3.902e-05 3.3 3.8939999999999996e-05 3.3 3.904e-05 0 3.896e-05 0 3.906e-05 3.3 3.8979999999999996e-05 3.3 3.908e-05 0 3.9e-05 0 3.91e-05 3.3 3.9019999999999996e-05 3.3 3.912e-05 0 3.904e-05 0 3.914e-05 3.3 3.9059999999999995e-05 3.3 3.916e-05 0 3.908e-05 0 3.918e-05 3.3 3.9099999999999995e-05 3.3 3.92e-05 0 3.912e-05 0 3.922e-05 3.3 3.9139999999999995e-05 3.3 3.924e-05 0 3.916e-05 0 3.926e-05 3.3 3.9179999999999994e-05 3.3 3.928e-05 0 3.92e-05 0 3.93e-05 3.3 3.9219999999999994e-05 3.3 3.9319999999999996e-05 0 3.924e-05 0 3.934e-05 3.3 3.9259999999999993e-05 3.3 3.9359999999999996e-05 0 3.928e-05 0 3.938e-05 3.3 3.93e-05 3.3 3.94e-05 0 3.9319999999999996e-05 0 3.942e-05 3.3 3.934e-05 3.3 3.944e-05 0 3.9359999999999996e-05 0 3.946e-05 3.3 3.938e-05 3.3 3.948e-05 0 3.9399999999999995e-05 0 3.95e-05 3.3 3.942e-05 3.3 3.952e-05 0 3.9439999999999995e-05 0 3.954e-05 3.3 3.946e-05 3.3 3.956e-05 0 3.9479999999999995e-05 0 3.958e-05 3.3 3.95e-05 3.3 3.96e-05 0 3.9519999999999994e-05 0 3.962e-05 3.3 3.954e-05 3.3 3.964e-05 0 3.9559999999999994e-05 0 3.9659999999999996e-05 3.3 3.958e-05 3.3 3.968e-05 0 3.9599999999999994e-05 0 3.9699999999999996e-05 3.3 3.962e-05 3.3 3.972e-05 0 3.964e-05 0 3.974e-05 3.3 3.9659999999999996e-05 3.3 3.976e-05 0 3.968e-05 0 3.978e-05 3.3 3.9699999999999996e-05 3.3 3.98e-05 0 3.972e-05 0 3.982e-05 3.3 3.9739999999999996e-05 3.3 3.984e-05 0 3.976e-05 0 3.986e-05 3.3 3.9779999999999995e-05 3.3 3.988e-05 0 3.98e-05 0 3.99e-05 3.3 3.9819999999999995e-05 3.3 3.992e-05 0 3.984e-05 0 3.994e-05 3.3 3.9859999999999994e-05 3.3 3.996e-05 0 3.988e-05 0 3.998e-05 3.3 3.9899999999999994e-05 3.3 3.9999999999999996e-05 0 3.992e-05 0 4.002e-05 3.3 3.9939999999999994e-05 3.3 4.0039999999999996e-05 0 3.996e-05 0 4.006e-05 3.3 3.998e-05 3.3 4.008e-05 0 3.9999999999999996e-05 0 4.01e-05 3.3 4.002e-05 3.3 4.012e-05 0 4.0039999999999996e-05 0 4.014e-05 3.3 4.006e-05 3.3 4.016e-05 0 4.0079999999999996e-05 0 4.018e-05 3.3 4.01e-05 3.3 4.02e-05 0 4.0119999999999995e-05 0 4.022e-05 3.3 4.014e-05 3.3 4.024e-05 0 4.0159999999999995e-05 0 4.026e-05 3.3 4.018e-05 3.3 4.028e-05 0 4.0199999999999995e-05 0 4.03e-05 3.3 4.022e-05 3.3 4.032e-05 0 4.0239999999999994e-05 0 4.034e-05 3.3 4.026e-05 3.3 4.036e-05 0 4.0279999999999994e-05 0 4.0379999999999996e-05 3.3 4.03e-05 3.3 4.04e-05 0 4.0319999999999993e-05 0 4.0419999999999996e-05 3.3 4.034e-05 3.3 4.044e-05 0 4.036e-05 0 4.046e-05 3.3 4.0379999999999996e-05 3.3 4.048e-05 0 4.04e-05 0 4.05e-05 3.3 4.0419999999999996e-05 3.3 4.052e-05 0 4.044e-05 0 4.054e-05 3.3 4.0459999999999995e-05 3.3 4.056e-05 0 4.048e-05 0 4.058e-05 3.3 4.0499999999999995e-05 3.3 4.06e-05 0 4.052e-05 0 4.062e-05 3.3 4.0539999999999995e-05 3.3 4.064e-05 0 4.056e-05 0 4.066e-05 3.3 4.0579999999999994e-05 3.3 4.068e-05 0 4.06e-05 0 4.07e-05 3.3 4.0619999999999994e-05 3.3 4.0719999999999996e-05 0 4.064e-05 0 4.074e-05 3.3 4.0659999999999994e-05 3.3 4.0759999999999996e-05 0 4.068e-05 0 4.078e-05 3.3 4.07e-05 3.3 4.08e-05 0 4.0719999999999996e-05 0 4.082e-05 3.3 4.074e-05 3.3 4.084e-05 0 4.0759999999999996e-05 0 4.086e-05 3.3 4.078e-05 3.3 4.088e-05 0 4.0799999999999996e-05 0 4.09e-05 3.3 4.082e-05 3.3 4.092e-05 0 4.0839999999999995e-05 0 4.094e-05 3.3 4.086e-05 3.3 4.096e-05 0 4.0879999999999995e-05 0 4.098e-05 3.3 4.09e-05 3.3 4.1e-05 0 4.0919999999999994e-05 0 4.102e-05 3.3 4.094e-05 3.3 4.104e-05 0 4.0959999999999994e-05 0 4.1059999999999997e-05 3.3 4.098e-05 3.3 4.108e-05 0 4.0999999999999994e-05 0 4.1099999999999996e-05 3.3 4.102e-05 3.3 4.112e-05 0 4.104e-05 0 4.114e-05 3.3 4.1059999999999997e-05 3.3 4.116e-05 0 4.108e-05 0 4.118e-05 3.3 4.1099999999999996e-05 3.3 4.12e-05 0 4.112e-05 0 4.122e-05 3.3 4.1139999999999996e-05 3.3 4.124e-05 0 4.116e-05 0 4.126e-05 3.3 4.1179999999999995e-05 3.3 4.128e-05 0 4.12e-05 0 4.13e-05 3.3 4.1219999999999995e-05 3.3 4.132e-05 0 4.124e-05 0 4.134e-05 3.3 4.1259999999999995e-05 3.3 4.136e-05 0 4.128e-05 0 4.138e-05 3.3 4.1299999999999994e-05 3.3 4.14e-05 0 4.132e-05 0 4.142e-05 3.3 4.1339999999999994e-05 3.3 4.1439999999999996e-05 0 4.136e-05 0 4.146e-05 3.3 4.1379999999999993e-05 3.3 4.1479999999999996e-05 0 4.14e-05 0 4.15e-05 3.3 4.142e-05 3.3 4.152e-05 0 4.1439999999999996e-05 0 4.154e-05 3.3 4.146e-05 3.3 4.156e-05 0 4.1479999999999996e-05 0 4.158e-05 3.3 4.15e-05 3.3 4.16e-05 0 4.1519999999999995e-05 0 4.162e-05 3.3 4.154e-05 3.3 4.164e-05 0 4.1559999999999995e-05 0 4.166e-05 3.3 4.158e-05 3.3 4.168e-05 0 4.1599999999999995e-05 0 4.17e-05 3.3 4.162e-05 3.3 4.172e-05 0 4.1639999999999994e-05 0 4.174e-05 3.3 4.166e-05 3.3 4.176e-05 0 4.1679999999999994e-05 0 4.1779999999999996e-05 3.3 4.17e-05 3.3 4.18e-05 0 4.1719999999999994e-05 0 4.1819999999999996e-05 3.3 4.174e-05 3.3 4.184e-05 0 4.176e-05 0 4.186e-05 3.3 4.1779999999999996e-05 3.3 4.188e-05 0 4.18e-05 0 4.19e-05 3.3 4.1819999999999996e-05 3.3 4.192e-05 0 4.184e-05 0 4.194e-05 3.3 4.1859999999999996e-05 3.3 4.196e-05 0 4.188e-05 0 4.198e-05 3.3 4.1899999999999995e-05 3.3 4.2e-05 0 4.192e-05 0 4.202e-05 3.3 4.1939999999999995e-05 3.3 4.204e-05 0 4.196e-05 0 4.206e-05 3.3 4.1979999999999994e-05 3.3 4.208e-05 0 4.2e-05 0 4.21e-05 3.3 4.2019999999999994e-05 3.3 4.2119999999999997e-05 0 4.204e-05 0 4.214e-05 3.3 4.2059999999999994e-05 3.3 4.2159999999999996e-05 0 4.208e-05 0 4.218e-05 3.3 4.21e-05 3.3 4.22e-05 0 4.2119999999999997e-05 0 4.222e-05 3.3 4.214e-05 3.3 4.224e-05 0 4.2159999999999996e-05 0 4.226e-05 3.3 4.218e-05 3.3 4.228e-05 0 4.2199999999999996e-05 0 4.23e-05 3.3 4.222e-05 3.3 4.232e-05 0 4.2239999999999995e-05 0 4.234e-05 3.3 4.226e-05 3.3 4.236e-05 0 4.2279999999999995e-05 0 4.238e-05 3.3 4.23e-05 3.3 4.24e-05 0 4.2319999999999995e-05 0 4.242e-05 3.3 4.234e-05 3.3 4.244e-05 0 4.2359999999999994e-05 0 4.246e-05 3.3 4.238e-05 3.3 4.248e-05 0 4.2399999999999994e-05 0 4.2499999999999996e-05 3.3 4.242e-05 3.3 4.252e-05 0 4.2439999999999993e-05 0 4.2539999999999996e-05 3.3 4.246e-05 3.3 4.256e-05 0 4.248e-05 0 4.258e-05 3.3 4.2499999999999996e-05 3.3 4.26e-05 0 4.252e-05 0 4.262e-05 3.3 4.2539999999999996e-05 3.3 4.264e-05 0 4.256e-05 0 4.266e-05 3.3 4.2579999999999996e-05 3.3 4.268e-05 0 4.26e-05 0 4.27e-05 3.3 4.2619999999999995e-05 3.3 4.272e-05 0 4.264e-05 0 4.274e-05 3.3 4.2659999999999995e-05 3.3 4.276e-05 0 4.268e-05 0 4.278e-05 3.3 4.2699999999999994e-05 3.3 4.28e-05 0 4.272e-05 0 4.282e-05 3.3 4.2739999999999994e-05 3.3 4.2839999999999996e-05 0 4.276e-05 0 4.286e-05 3.3 4.2779999999999994e-05 3.3 4.2879999999999996e-05 0 4.28e-05 0 4.29e-05 3.3 4.282e-05 3.3 4.292e-05 0 4.2839999999999996e-05 0 4.294e-05 3.3 4.286e-05 3.3 4.296e-05 0 4.2879999999999996e-05 0 4.298e-05 3.3 4.29e-05 3.3 4.3e-05 0 4.2919999999999996e-05 0 4.302e-05 3.3 4.294e-05 3.3 4.304e-05 0 4.2959999999999995e-05 0 4.306e-05 3.3 4.298e-05 3.3 4.308e-05 0 4.2999999999999995e-05 0 4.31e-05 3.3 4.302e-05 3.3 4.312e-05 0 4.3039999999999994e-05 0 4.314e-05 3.3 4.306e-05 3.3 4.316e-05 0 4.3079999999999994e-05 0 4.3179999999999997e-05 3.3 4.31e-05 3.3 4.32e-05 0 4.3119999999999994e-05 0 4.3219999999999996e-05 3.3 4.314e-05 3.3 4.324e-05 0 4.315999999999999e-05 0 4.3259999999999996e-05 3.3 4.3179999999999997e-05 3.3 4.328e-05 0 4.32e-05 0 4.33e-05 3.3 4.3219999999999996e-05 3.3 4.332e-05 0 4.324e-05 0 4.334e-05 3.3 4.3259999999999996e-05 3.3 4.336e-05 0 4.328e-05 0 4.338e-05 3.3 4.3299999999999995e-05 3.3 4.34e-05 0 4.332e-05 0 4.342e-05 3.3 4.3339999999999995e-05 3.3 4.344e-05 0 4.336e-05 0 4.346e-05 3.3 4.3379999999999995e-05 3.3 4.348e-05 0 4.34e-05 0 4.35e-05 3.3 4.3419999999999994e-05 3.3 4.352e-05 0 4.344e-05 0 4.354e-05 3.3 4.3459999999999994e-05 3.3 4.3559999999999996e-05 0 4.348e-05 0 4.358e-05 3.3 4.3499999999999993e-05 3.3 4.3599999999999996e-05 0 4.352e-05 0 4.362e-05 3.3 4.354e-05 3.3 4.364e-05 0 4.3559999999999996e-05 0 4.366e-05 3.3 4.358e-05 3.3 4.368e-05 0 4.3599999999999996e-05 0 4.37e-05 3.3 4.362e-05 3.3 4.372e-05 0 4.3639999999999996e-05 0 4.374e-05 3.3 4.366e-05 3.3 4.376e-05 0 4.3679999999999995e-05 0 4.378e-05 3.3 4.37e-05 3.3 4.38e-05 0 4.3719999999999995e-05 0 4.382e-05 3.3 4.374e-05 3.3 4.384e-05 0 4.3759999999999994e-05 0 4.386e-05 3.3 4.378e-05 3.3 4.388e-05 0 4.3799999999999994e-05 0 4.3899999999999996e-05 3.3 4.382e-05 3.3 4.392e-05 0 4.3839999999999994e-05 0 4.3939999999999996e-05 3.3 4.386e-05 3.3 4.396e-05 0 4.388e-05 0 4.398e-05 3.3 4.3899999999999996e-05 3.3 4.4e-05 0 4.392e-05 0 4.402e-05 3.3 4.3939999999999996e-05 3.3 4.404e-05 0 4.396e-05 0 4.406e-05 3.3 4.3979999999999996e-05 3.3 4.408e-05 0 4.4e-05 0 4.41e-05 3.3 4.4019999999999995e-05 3.3 4.412e-05 0 4.404e-05 0 4.414e-05 3.3 4.4059999999999995e-05 3.3 4.416e-05 0 4.408e-05 0 4.418e-05 3.3 4.4099999999999995e-05 3.3 4.42e-05 0 4.412e-05 0 4.422e-05 3.3 4.4139999999999994e-05 3.3 4.4239999999999997e-05 0 4.416e-05 0 4.426e-05 3.3 4.4179999999999994e-05 3.3 4.4279999999999996e-05 0 4.42e-05 0 4.43e-05 3.3 4.421999999999999e-05 3.3 4.4319999999999996e-05 0 4.4239999999999997e-05 0 4.434e-05 3.3 4.426e-05 3.3 4.436e-05 0 4.4279999999999996e-05 0 4.438e-05 3.3 4.43e-05 3.3 4.44e-05 0 4.4319999999999996e-05 0 4.442e-05 3.3 4.434e-05 3.3 4.444e-05 0 4.4359999999999995e-05 0 4.446e-05 3.3 4.438e-05 3.3 4.448e-05 0 4.4399999999999995e-05 0 4.45e-05 3.3 4.442e-05 3.3 4.452e-05 0 4.4439999999999995e-05 0 4.454e-05 3.3 4.446e-05 3.3 4.456e-05 0 4.4479999999999994e-05 0 4.458e-05 3.3 4.45e-05 3.3 4.46e-05 0 4.4519999999999994e-05 0 4.4619999999999996e-05 3.3 4.454e-05 3.3 4.464e-05 0 4.4559999999999993e-05 0 4.4659999999999996e-05 3.3 4.458e-05 3.3 4.468e-05 0 4.46e-05 0 4.47e-05 3.3 4.4619999999999996e-05 3.3 4.472e-05 0 4.464e-05 0 4.474e-05 3.3 4.4659999999999996e-05 3.3 4.476e-05 0 4.468e-05 0 4.478e-05 3.3 4.4699999999999996e-05 3.3 4.48e-05 0 4.472e-05 0 4.482e-05 3.3 4.4739999999999995e-05 3.3 4.484e-05 0 4.476e-05 0 4.486e-05 3.3 4.4779999999999995e-05 3.3 4.488e-05 0 4.48e-05 0 4.49e-05 3.3 4.4819999999999994e-05 3.3 4.492e-05 0 4.484e-05 0 4.494e-05 3.3 4.4859999999999994e-05 3.3 4.4959999999999996e-05 0 4.488e-05 0 4.498e-05 3.3 4.4899999999999994e-05 3.3 4.4999999999999996e-05 0 4.492e-05 0 4.502e-05 3.3 4.494e-05 3.3 4.504e-05 0 4.4959999999999996e-05 0 4.506e-05 3.3 4.498e-05 3.3 4.508e-05 0 4.4999999999999996e-05 0 4.51e-05 3.3 4.502e-05 3.3 4.512e-05 0 4.5039999999999996e-05 0 4.514e-05 3.3 4.506e-05 3.3 4.516e-05 0 4.5079999999999995e-05 0 4.518e-05 3.3 4.51e-05 3.3 4.52e-05 0 4.5119999999999995e-05 0 4.522e-05 3.3 4.514e-05 3.3 4.524e-05 0 4.5159999999999995e-05 0 4.526e-05 3.3 4.518e-05 3.3 4.528e-05 0 4.5199999999999994e-05 0 4.5299999999999997e-05 3.3 4.522e-05 3.3 4.532e-05 0 4.5239999999999994e-05 0 4.5339999999999996e-05 3.3 4.526e-05 3.3 4.536e-05 0 4.527999999999999e-05 0 4.5379999999999996e-05 3.3 4.5299999999999997e-05 3.3 4.54e-05 0 4.532e-05 0 4.542e-05 3.3 4.5339999999999996e-05 3.3 4.544e-05 0 4.536e-05 0 4.546e-05 3.3 4.5379999999999996e-05 3.3 4.548e-05 0 4.54e-05 0 4.55e-05 3.3 4.5419999999999995e-05 3.3 4.552e-05 0 4.544e-05 0 4.554e-05 3.3 4.5459999999999995e-05 3.3 4.556e-05 0 4.548e-05 0 4.558e-05 3.3 4.5499999999999995e-05 3.3 4.56e-05 0 4.552e-05 0 4.562e-05 3.3 4.5539999999999994e-05 3.3 4.564e-05 0 4.556e-05 0 4.566e-05 3.3 4.5579999999999994e-05 3.3 4.5679999999999996e-05 0 4.56e-05 0 4.57e-05 3.3 4.5619999999999994e-05 3.3 4.5719999999999996e-05 0 4.564e-05 0 4.574e-05 3.3 4.566e-05 3.3 4.576e-05 0 4.5679999999999996e-05 0 4.578e-05 3.3 4.57e-05 3.3 4.58e-05 0 4.5719999999999996e-05 0 4.582e-05 3.3 4.574e-05 3.3 4.584e-05 0 4.5759999999999996e-05 0 4.586e-05 3.3 4.578e-05 3.3 4.588e-05 0 4.5799999999999995e-05 0 4.59e-05 3.3 4.582e-05 3.3 4.592e-05 0 4.5839999999999995e-05 0 4.594e-05 3.3 4.586e-05 3.3 4.596e-05 0 4.5879999999999994e-05 0 4.598e-05 3.3 4.59e-05 3.3 4.6e-05 0 4.5919999999999994e-05 0 4.6019999999999996e-05 3.3 4.594e-05 3.3 4.604e-05 0 4.5959999999999994e-05 0 4.6059999999999996e-05 3.3 4.598e-05 3.3 4.608e-05 0 4.599999999999999e-05 0 4.6099999999999996e-05 3.3 4.6019999999999996e-05 3.3 4.612e-05 0 4.604e-05 0 4.614e-05 3.3 4.6059999999999996e-05 3.3 4.616e-05 0 4.608e-05 0 4.618e-05 3.3 4.6099999999999996e-05 3.3 4.62e-05 0 4.612e-05 0 4.622e-05 3.3 4.6139999999999995e-05 3.3 4.624e-05 0 4.616e-05 0 4.626e-05 3.3 4.6179999999999995e-05 3.3 4.628e-05 0 4.62e-05 0 4.63e-05 3.3 4.6219999999999995e-05 3.3 4.632e-05 0 4.624e-05 0 4.634e-05 3.3 4.6259999999999994e-05 3.3 4.6359999999999997e-05 0 4.628e-05 0 4.638e-05 3.3 4.6299999999999994e-05 3.3 4.6399999999999996e-05 0 4.632e-05 0 4.642e-05 3.3 4.6339999999999993e-05 3.3 4.6439999999999996e-05 0 4.6359999999999997e-05 0 4.646e-05 3.3 4.638e-05 3.3 4.648e-05 0 4.6399999999999996e-05 0 4.65e-05 3.3 4.642e-05 3.3 4.652e-05 0 4.6439999999999996e-05 0 4.654e-05 3.3 4.646e-05 3.3 4.656e-05 0 4.6479999999999995e-05 0 4.658e-05 3.3 4.65e-05 3.3 4.66e-05 0 4.6519999999999995e-05 0 4.662e-05 3.3 4.654e-05 3.3 4.664e-05 0 4.6559999999999995e-05 0 4.666e-05 3.3 4.658e-05 3.3 4.668e-05 0 4.6599999999999994e-05 0 4.67e-05 3.3 4.662e-05 3.3 4.672e-05 0 4.6639999999999994e-05 0 4.6739999999999996e-05 3.3 4.666e-05 3.3 4.676e-05 0 4.6679999999999994e-05 0 4.6779999999999996e-05 3.3 4.67e-05 3.3 4.68e-05 0 4.672e-05 0 4.682e-05 3.3 4.6739999999999996e-05 3.3 4.684e-05 0 4.676e-05 0 4.686e-05 3.3 4.6779999999999996e-05 3.3 4.688e-05 0 4.68e-05 0 4.69e-05 3.3 4.6819999999999996e-05 3.3 4.692e-05 0 4.684e-05 0 4.694e-05 3.3 4.6859999999999995e-05 3.3 4.696e-05 0 4.688e-05 0 4.698e-05 3.3 4.6899999999999995e-05 3.3 4.7e-05 0 4.692e-05 0 4.702e-05 3.3 4.6939999999999994e-05 3.3 4.704e-05 0 4.696e-05 0 4.706e-05 3.3 4.6979999999999994e-05 3.3 4.7079999999999996e-05 0 4.7e-05 0 4.71e-05 3.3 4.7019999999999994e-05 3.3 4.7119999999999996e-05 0 4.704e-05 0 4.714e-05 3.3 4.705999999999999e-05 3.3 4.7159999999999996e-05 0 4.7079999999999996e-05 0 4.718e-05 3.3 4.71e-05 3.3 4.72e-05 0 4.7119999999999996e-05 0 4.722e-05 3.3 4.714e-05 3.3 4.724e-05 0 4.7159999999999996e-05 0 4.726e-05 3.3 4.718e-05 3.3 4.728e-05 0 4.7199999999999995e-05 0 4.73e-05 3.3 4.722e-05 3.3 4.732e-05 0 4.7239999999999995e-05 0 4.734e-05 3.3 4.726e-05 3.3 4.736e-05 0 4.7279999999999995e-05 0 4.738e-05 3.3 4.73e-05 3.3 4.74e-05 0 4.7319999999999994e-05 0 4.7419999999999997e-05 3.3 4.734e-05 3.3 4.744e-05 0 4.7359999999999994e-05 0 4.7459999999999996e-05 3.3 4.738e-05 3.3 4.748e-05 0 4.7399999999999993e-05 0 4.7499999999999996e-05 3.3 4.7419999999999997e-05 3.3 4.752e-05 0 4.744e-05 0 4.754e-05 3.3 4.7459999999999996e-05 3.3 4.756e-05 0 4.748e-05 0 4.758e-05 3.3 4.7499999999999996e-05 3.3 4.76e-05 0 4.752e-05 0 4.762e-05 3.3 4.7539999999999995e-05 3.3 4.764e-05 0 4.756e-05 0 4.766e-05 3.3 4.7579999999999995e-05 3.3 4.768e-05 0 4.76e-05 0 4.77e-05 3.3 4.7619999999999995e-05 3.3 4.772e-05 0 4.764e-05 0 4.774e-05 3.3 4.7659999999999994e-05 3.3 4.776e-05 0 4.768e-05 0 4.778e-05 3.3 4.7699999999999994e-05 3.3 4.7799999999999996e-05 0 4.772e-05 0 4.782e-05 3.3 4.7739999999999994e-05 3.3 4.7839999999999996e-05 0 4.776e-05 0 4.786e-05 3.3 4.778e-05 3.3 4.788e-05 0 4.7799999999999996e-05 0 4.79e-05 3.3 4.782e-05 3.3 4.792e-05 0 4.7839999999999996e-05 0 4.794e-05 3.3 4.786e-05 3.3 4.796e-05 0 4.7879999999999996e-05 0 4.798e-05 3.3 4.79e-05 3.3 4.8e-05 0 4.7919999999999995e-05 0 4.802e-05 3.3 4.794e-05 3.3 4.804e-05 0 4.7959999999999995e-05 0 4.806e-05 3.3 4.798e-05 3.3 4.808e-05 0 4.7999999999999994e-05 0 4.81e-05 3.3 4.802e-05 3.3 4.812e-05 0 4.8039999999999994e-05 0 4.8139999999999996e-05 3.3 4.806e-05 3.3 4.816e-05 0 4.8079999999999994e-05 0 4.8179999999999996e-05 3.3 4.81e-05 3.3 4.82e-05 0 4.811999999999999e-05 0 4.8219999999999996e-05 3.3 4.8139999999999996e-05 3.3 4.824e-05 0 4.816e-05 0 4.826e-05 3.3 4.8179999999999996e-05 3.3 4.828e-05 0 4.82e-05 0 4.83e-05 3.3 4.8219999999999996e-05 3.3 4.832e-05 0 4.824e-05 0 4.834e-05 3.3 4.8259999999999995e-05 3.3 4.836e-05 0 4.828e-05 0 4.838e-05 3.3 4.8299999999999995e-05 3.3 4.84e-05 0 4.832e-05 0 4.842e-05 3.3 4.8339999999999995e-05 3.3 4.844e-05 0 4.836e-05 0 4.846e-05 3.3 4.8379999999999994e-05 3.3 4.848e-05 0 4.84e-05 0 4.85e-05 3.3 4.8419999999999994e-05 3.3 4.8519999999999996e-05 0 4.844e-05 0 4.854e-05 3.3 4.8459999999999993e-05 3.3 4.8559999999999996e-05 0 4.848e-05 0 4.858e-05 3.3 4.85e-05 3.3 4.86e-05 0 4.8519999999999996e-05 0 4.862e-05 3.3 4.854e-05 3.3 4.864e-05 0 4.8559999999999996e-05 0 4.866e-05 3.3 4.858e-05 3.3 4.868e-05 0 4.8599999999999995e-05 0 4.87e-05 3.3 4.862e-05 3.3 4.872e-05 0 4.8639999999999995e-05 0 4.874e-05 3.3 4.866e-05 3.3 4.876e-05 0 4.8679999999999995e-05 0 4.878e-05 3.3 4.87e-05 3.3 4.88e-05 0 4.8719999999999994e-05 0 4.882e-05 3.3 4.874e-05 3.3 4.884e-05 0 4.8759999999999994e-05 0 4.8859999999999996e-05 3.3 4.878e-05 3.3 4.888e-05 0 4.8799999999999994e-05 0 4.8899999999999996e-05 3.3 4.882e-05 3.3 4.892e-05 0 4.884e-05 0 4.894e-05 3.3 4.8859999999999996e-05 3.3 4.896e-05 0 4.888e-05 0 4.898e-05 3.3 4.8899999999999996e-05 3.3 4.9e-05 0 4.892e-05 0 4.902e-05 3.3 4.8939999999999996e-05 3.3 4.904e-05 0 4.896e-05 0 4.906e-05 3.3 4.8979999999999995e-05 3.3 4.908e-05 0 4.9e-05 0 4.91e-05 3.3 4.9019999999999995e-05 3.3 4.912e-05 0 4.904e-05 0 4.914e-05 3.3 4.9059999999999994e-05 3.3 4.916e-05 0 4.908e-05 0 4.918e-05 3.3 4.9099999999999994e-05 3.3 4.9199999999999997e-05 0 4.912e-05 0 4.922e-05 3.3 4.9139999999999994e-05 3.3 4.9239999999999996e-05 0 4.916e-05 0 4.926e-05 3.3 4.917999999999999e-05 3.3 4.9279999999999996e-05 0 4.9199999999999997e-05 0 4.93e-05 3.3 4.922e-05 3.3 4.932e-05 0 4.9239999999999996e-05 0 4.934e-05 3.3 4.926e-05 3.3 4.936e-05 0 4.9279999999999996e-05 0 4.938e-05 3.3 4.93e-05 3.3 4.94e-05 0 4.9319999999999995e-05 0 4.942e-05 3.3 4.934e-05 3.3 4.944e-05 0 4.9359999999999995e-05 0 4.946e-05 3.3 4.938e-05 3.3 4.948e-05 0 4.9399999999999995e-05 0 4.95e-05 3.3 4.942e-05 3.3 4.952e-05 0 4.9439999999999994e-05 0 4.954e-05 3.3 4.946e-05 3.3 4.956e-05 0 4.9479999999999994e-05 0 4.9579999999999996e-05 3.3 4.95e-05 3.3 4.96e-05 0 4.9519999999999993e-05 0 4.9619999999999996e-05 3.3 4.954e-05 3.3 4.964e-05 0 4.956e-05 0 4.966e-05 3.3 4.9579999999999996e-05 3.3 4.968e-05 0 4.96e-05 0 4.97e-05 3.3 4.9619999999999996e-05 3.3 4.972e-05 0 4.964e-05 0 4.974e-05 3.3 4.9659999999999995e-05 3.3 4.976e-05 0 4.968e-05 0 4.978e-05 3.3 4.9699999999999995e-05 3.3 4.98e-05 0 4.972e-05 0 4.982e-05 3.3 4.9739999999999995e-05 3.3 4.984e-05 0 4.976e-05 0 4.986e-05 3.3 4.9779999999999994e-05 3.3 4.988e-05 0 4.98e-05 0 4.99e-05 3.3 4.9819999999999994e-05 3.3 4.9919999999999996e-05 0 4.984e-05 0 4.994e-05 3.3 4.9859999999999994e-05 3.3 4.9959999999999996e-05 0 4.988e-05 0 4.998e-05 3.3 4.989999999999999e-05 3.3 4.9999999999999996e-05 0 4.9919999999999996e-05 0 5.002e-05 3.3 4.994e-05 3.3 5.004e-05 0 4.9959999999999996e-05 0 5.006e-05 3.3 4.998e-05 3.3 5.008e-05 0 4.9999999999999996e-05 0 5.01e-05 3.3 5.002e-05 3.3 5.012e-05 0 5.0039999999999995e-05 0 5.014e-05 3.3 5.006e-05 3.3 5.016e-05 0 5.0079999999999995e-05 0 5.018e-05 3.3 5.01e-05 3.3 5.02e-05 0 5.0119999999999994e-05 0 5.022e-05 3.3 5.014e-05 3.3 5.024e-05 0 5.0159999999999994e-05 0 5.0259999999999997e-05 3.3 5.018e-05 3.3 5.028e-05 0 5.0199999999999994e-05 0 5.0299999999999996e-05 3.3 5.022e-05 3.3 5.032e-05 0 5.023999999999999e-05 0 5.0339999999999996e-05 3.3 5.0259999999999997e-05 3.3 5.036e-05 0 5.028e-05 0 5.038e-05 3.3 5.0299999999999996e-05 3.3 5.04e-05 0 5.032e-05 0 5.042e-05 3.3 5.0339999999999996e-05 3.3 5.044e-05 0 5.036e-05 0 5.046e-05 3.3 5.0379999999999995e-05 3.3 5.048e-05 0 5.04e-05 0 5.05e-05 3.3 5.0419999999999995e-05 3.3 5.052e-05 0 5.044e-05 0 5.054e-05 3.3 5.0459999999999995e-05 3.3 5.056e-05 0 5.048e-05 0 5.058e-05 3.3 5.0499999999999994e-05 3.3 5.06e-05 0 5.052e-05 0 5.062e-05 3.3 5.0539999999999994e-05 3.3 5.0639999999999996e-05 0 5.056e-05 0 5.066e-05 3.3 5.0579999999999993e-05 3.3 5.0679999999999996e-05 0 5.06e-05 0 5.07e-05 3.3 5.062e-05 3.3 5.072e-05 0 5.0639999999999996e-05 0 5.074e-05 3.3 5.066e-05 3.3 5.076e-05 0 5.0679999999999996e-05 0 5.078e-05 3.3 5.07e-05 3.3 5.08e-05 0 5.0719999999999996e-05 0 5.082e-05 3.3 5.074e-05 3.3 5.084e-05 0 5.0759999999999995e-05 0 5.086e-05 3.3 5.078e-05 3.3 5.088e-05 0 5.0799999999999995e-05 0 5.09e-05 3.3 5.082e-05 3.3 5.092e-05 0 5.0839999999999994e-05 0 5.094e-05 3.3 5.086e-05 3.3 5.096e-05 0 5.0879999999999994e-05 0 5.0979999999999996e-05 3.3 5.09e-05 3.3 5.1e-05 0 5.0919999999999994e-05 0 5.1019999999999996e-05 3.3 5.094e-05 3.3 5.104e-05 0 5.095999999999999e-05 0 5.1059999999999996e-05 3.3 5.0979999999999996e-05 3.3 5.108e-05 0 5.1e-05 0 5.11e-05 3.3 5.1019999999999996e-05 3.3 5.112e-05 0 5.104e-05 0 5.114e-05 3.3 5.1059999999999996e-05 3.3 5.116e-05 0 5.108e-05 0 5.118e-05 3.3 5.1099999999999995e-05 3.3 5.12e-05 0 5.112e-05 0 5.122e-05 3.3 5.1139999999999995e-05 3.3 5.124e-05 0 5.116e-05 0 5.126e-05 3.3 5.1179999999999994e-05 3.3 5.128e-05 0 5.12e-05 0 5.13e-05 3.3 5.1219999999999994e-05 3.3 5.1319999999999997e-05 0 5.124e-05 0 5.134e-05 3.3 5.1259999999999994e-05 3.3 5.1359999999999996e-05 0 5.128e-05 0 5.138e-05 3.3 5.129999999999999e-05 3.3 5.1399999999999996e-05 0 5.1319999999999997e-05 0 5.142e-05 3.3 5.134e-05 3.3 5.144e-05 0 5.1359999999999996e-05 0 5.146e-05 3.3 5.138e-05 3.3 5.148e-05 0 5.1399999999999996e-05 0 5.15e-05 3.3 5.142e-05 3.3 5.152e-05 0 5.1439999999999995e-05 0 5.154e-05 3.3 5.146e-05 3.3 5.156e-05 0 5.1479999999999995e-05 0 5.158e-05 3.3 5.15e-05 3.3 5.16e-05 0 5.1519999999999995e-05 0 5.162e-05 3.3 5.154e-05 3.3 5.164e-05 0 5.1559999999999994e-05 0 5.166e-05 3.3 5.158e-05 3.3 5.168e-05 0 5.1599999999999994e-05 0 5.1699999999999996e-05 3.3 5.162e-05 3.3 5.172e-05 0 5.1639999999999993e-05 0 5.1739999999999996e-05 3.3 5.166e-05 3.3 5.176e-05 0 5.168e-05 0 5.178e-05 3.3 5.1699999999999996e-05 3.3 5.18e-05 0 5.172e-05 0 5.182e-05 3.3 5.1739999999999996e-05 3.3 5.184e-05 0 5.176e-05 0 5.186e-05 3.3 5.1779999999999996e-05 3.3 5.188e-05 0 5.18e-05 0 5.19e-05 3.3 5.1819999999999995e-05 3.3 5.192e-05 0 5.184e-05 0 5.194e-05 3.3 5.1859999999999995e-05 3.3 5.196e-05 0 5.188e-05 0 5.198e-05 3.3 5.1899999999999994e-05 3.3 5.2e-05 0 5.192e-05 0 5.202e-05 3.3 5.1939999999999994e-05 3.3 5.2039999999999996e-05 0 5.196e-05 0 5.206e-05 3.3 5.1979999999999994e-05 3.3 5.2079999999999996e-05 0 5.2e-05 0 5.21e-05 3.3 5.201999999999999e-05 3.3 5.2119999999999996e-05 0 5.2039999999999996e-05 0 5.214e-05 3.3 5.206e-05 3.3 5.216e-05 0 5.2079999999999996e-05 0 5.218e-05 3.3 5.21e-05 3.3 5.22e-05 0 5.2119999999999996e-05 0 5.222e-05 3.3 5.214e-05 3.3 5.224e-05 0 5.2159999999999995e-05 0 5.226e-05 3.3 5.218e-05 3.3 5.228e-05 0 5.2199999999999995e-05 0 5.23e-05 3.3 5.222e-05 3.3 5.232e-05 0 5.2239999999999995e-05 0 5.234e-05 3.3 5.226e-05 3.3 5.236e-05 0 5.2279999999999994e-05 0 5.2379999999999997e-05 3.3 5.23e-05 3.3 5.24e-05 0 5.2319999999999994e-05 0 5.2419999999999996e-05 3.3 5.234e-05 3.3 5.244e-05 0 5.235999999999999e-05 0 5.2459999999999996e-05 3.3 5.2379999999999997e-05 3.3 5.248e-05 0 5.24e-05 0 5.25e-05 3.3 5.2419999999999996e-05 3.3 5.252e-05 0 5.244e-05 0 5.254e-05 3.3 5.2459999999999996e-05 3.3 5.256e-05 0 5.248e-05 0 5.258e-05 3.3 5.2499999999999995e-05 3.3 5.26e-05 0 5.252e-05 0 5.262e-05 3.3 5.2539999999999995e-05 3.3 5.264e-05 0 5.256e-05 0 5.266e-05 3.3 5.2579999999999995e-05 3.3 5.268e-05 0 5.26e-05 0 5.27e-05 3.3 5.2619999999999994e-05 3.3 5.272e-05 0 5.264e-05 0 5.274e-05 3.3 5.2659999999999994e-05 3.3 5.2759999999999996e-05 0 5.268e-05 0 5.278e-05 3.3 5.2699999999999993e-05 3.3 5.2799999999999996e-05 0 5.272e-05 0 5.282e-05 3.3 5.274e-05 3.3 5.284e-05 0 5.2759999999999996e-05 0 5.286e-05 3.3 5.278e-05 3.3 5.288e-05 0 5.2799999999999996e-05 0 5.29e-05 3.3 5.282e-05 3.3 5.292e-05 0 5.2839999999999996e-05 0 5.294e-05 3.3 5.286e-05 3.3 5.296e-05 0 5.2879999999999995e-05 0 5.298e-05 3.3 5.29e-05 3.3 5.3e-05 0 5.2919999999999995e-05 0 5.302e-05 3.3 5.294e-05 3.3 5.304e-05 0 5.2959999999999994e-05 0 5.306e-05 3.3 5.298e-05 3.3 5.308e-05 0 5.2999999999999994e-05 0 5.3099999999999996e-05 3.3 5.302e-05 3.3 5.312e-05 0 5.3039999999999994e-05 0 5.3139999999999996e-05 3.3 5.306e-05 3.3 5.316e-05 0 5.307999999999999e-05 0 5.3179999999999996e-05 3.3 5.3099999999999996e-05 3.3 5.32e-05 0 5.312e-05 0 5.322e-05 3.3 5.3139999999999996e-05 3.3 5.324e-05 0 5.316e-05 0 5.326e-05 3.3 5.3179999999999996e-05 3.3 5.328e-05 0 5.32e-05 0 5.33e-05 3.3 5.3219999999999995e-05 3.3 5.332e-05 0 5.324e-05 0 5.334e-05 3.3 5.3259999999999995e-05 3.3 5.336e-05 0 5.328e-05 0 5.338e-05 3.3 5.3299999999999995e-05 3.3 5.34e-05 0 5.332e-05 0 5.342e-05 3.3 5.3339999999999994e-05 3.3 5.3439999999999997e-05 0 5.336e-05 0 5.346e-05 3.3 5.3379999999999994e-05 3.3 5.3479999999999996e-05 0 5.34e-05 0 5.35e-05 3.3 5.341999999999999e-05 3.3 5.3519999999999996e-05 0 5.3439999999999997e-05 0 5.354e-05 3.3 5.346e-05 3.3 5.356e-05 0 5.3479999999999996e-05 0 5.358e-05 3.3 5.35e-05 3.3 5.36e-05 0 5.3519999999999996e-05 0 5.362e-05 3.3 5.354e-05 3.3 5.364e-05 0 5.3559999999999995e-05 0 5.366e-05 3.3 5.358e-05 3.3 5.368e-05 0 5.3599999999999995e-05 0 5.37e-05 3.3 5.362e-05 3.3 5.372e-05 0 5.3639999999999995e-05 0 5.374e-05 3.3 5.366e-05 3.3 5.376e-05 0 5.3679999999999994e-05 0 5.378e-05 3.3 5.37e-05 3.3 5.38e-05 0 5.3719999999999994e-05 0 5.3819999999999996e-05 3.3 5.374e-05 3.3 5.384e-05 0 5.3759999999999994e-05 0 5.3859999999999996e-05 3.3 5.378e-05 3.3 5.388e-05 0 5.379999999999999e-05 0 5.3899999999999996e-05 3.3 5.3819999999999996e-05 3.3 5.392e-05 0 5.384e-05 0 5.394e-05 3.3 5.3859999999999996e-05 3.3 5.396e-05 0 5.388e-05 0 5.398e-05 3.3 5.3899999999999996e-05 3.3 5.4e-05 0 5.392e-05 0 5.402e-05 3.3 5.3939999999999995e-05 3.3 5.404e-05 0 5.396e-05 0 5.406e-05 3.3 5.3979999999999995e-05 3.3 5.408e-05 0 5.4e-05 0 5.41e-05 3.3 5.4019999999999994e-05 3.3 5.412e-05 0 5.404e-05 0 5.414e-05 3.3 5.4059999999999994e-05 3.3 5.4159999999999996e-05 0 5.408e-05 0 5.418e-05 3.3 5.4099999999999994e-05 3.3 5.4199999999999996e-05 0 5.412e-05 0 5.422e-05 3.3 5.413999999999999e-05 3.3 5.4239999999999996e-05 0 5.4159999999999996e-05 0 5.426e-05 3.3 5.418e-05 3.3 5.428e-05 0 5.4199999999999996e-05 0 5.43e-05 3.3 5.422e-05 3.3 5.432e-05 0 5.4239999999999996e-05 0 5.434e-05 3.3 5.426e-05 3.3 5.436e-05 0 5.4279999999999995e-05 0 5.438e-05 3.3 5.43e-05 3.3 5.44e-05 0 5.4319999999999995e-05 0 5.442e-05 3.3 5.434e-05 3.3 5.444e-05 0 5.4359999999999995e-05 0 5.446e-05 3.3 5.438e-05 3.3 5.448e-05 0 5.4399999999999994e-05 0 5.4499999999999997e-05 3.3 5.442e-05 3.3 5.452e-05 0 5.4439999999999994e-05 0 5.4539999999999996e-05 3.3 5.446e-05 3.3 5.456e-05 0 5.447999999999999e-05 0 5.4579999999999996e-05 3.3 5.4499999999999997e-05 3.3 5.46e-05 0 5.452e-05 0 5.462e-05 3.3 5.4539999999999996e-05 3.3 5.464e-05 0 5.456e-05 0 5.466e-05 3.3 5.4579999999999996e-05 3.3 5.468e-05 0 5.46e-05 0 5.47e-05 3.3 5.4619999999999995e-05 3.3 5.472e-05 0 5.464e-05 0 5.474e-05 3.3 5.4659999999999995e-05 3.3 5.476e-05 0 5.468e-05 0 5.478e-05 3.3 5.4699999999999995e-05 3.3 5.48e-05 0 5.472e-05 0 5.482e-05 3.3 5.4739999999999994e-05 3.3 5.484e-05 0 5.476e-05 0 5.486e-05 3.3 5.4779999999999994e-05 3.3 5.4879999999999996e-05 0 5.48e-05 0 5.49e-05 3.3 5.4819999999999994e-05 3.3 5.4919999999999996e-05 0 5.484e-05 0 5.494e-05 3.3 5.485999999999999e-05 3.3 5.4959999999999996e-05 0 5.4879999999999996e-05 0 5.498e-05 3.3 5.49e-05 3.3 5.5e-05 0 5.4919999999999996e-05 0 5.502e-05 3.3 5.494e-05 3.3 5.504e-05 0 5.4959999999999996e-05 0 5.506e-05 3.3 5.498e-05 3.3 5.508e-05 0 5.4999999999999995e-05 0 5.51e-05 3.3 5.502e-05 3.3 5.512e-05 0 5.5039999999999995e-05 0 5.514e-05 3.3 5.506e-05 3.3 5.516e-05 0 5.5079999999999994e-05 0 5.518e-05 3.3 5.51e-05 3.3 5.52e-05 0 5.5119999999999994e-05 0 5.5219999999999996e-05 3.3 5.514e-05 3.3 5.524e-05 0 5.5159999999999994e-05 0 5.5259999999999996e-05 3.3 5.518e-05 3.3 5.528e-05 0 5.519999999999999e-05 0 5.5299999999999996e-05 3.3 5.5219999999999996e-05 3.3 5.532e-05 0 5.524e-05 0 5.534e-05 3.3 5.5259999999999996e-05 3.3 5.536e-05 0 5.528e-05 0 5.538e-05 3.3 5.5299999999999996e-05 3.3 5.54e-05 0 5.532e-05 0 5.542e-05 3.3 5.5339999999999995e-05 3.3 5.544e-05 0 5.536e-05 0 5.546e-05 3.3 5.5379999999999995e-05 3.3 5.548e-05 0 5.54e-05 0 5.55e-05 3.3 5.5419999999999995e-05 3.3 5.552e-05 0 5.544e-05 0 5.554e-05 3.3 5.5459999999999994e-05 3.3 5.5559999999999997e-05 0 5.548e-05 0 5.558e-05 3.3 5.5499999999999994e-05 3.3 5.5599999999999996e-05 0 5.552e-05 0 5.562e-05 3.3 5.5539999999999993e-05 3.3 5.5639999999999996e-05 0 5.5559999999999997e-05 0 5.566e-05 3.3 5.558e-05 3.3 5.568e-05 0 5.5599999999999996e-05 0 5.57e-05 3.3 5.562e-05 3.3 5.572e-05 0 5.5639999999999996e-05 0 5.574e-05 3.3 5.566e-05 3.3 5.576e-05 0 5.5679999999999995e-05 0 5.578e-05 3.3 5.57e-05 3.3 5.58e-05 0 5.5719999999999995e-05 0 5.582e-05 3.3 5.574e-05 3.3 5.584e-05 0 5.5759999999999995e-05 0 5.586e-05 3.3 5.578e-05 3.3 5.588e-05 0 5.5799999999999994e-05 0 5.59e-05 3.3 5.582e-05 3.3 5.592e-05 0 5.5839999999999994e-05 0 5.5939999999999996e-05 3.3 5.586e-05 3.3 5.596e-05 0 5.5879999999999994e-05 0 5.5979999999999996e-05 3.3 5.59e-05 3.3 5.6e-05 0 5.591999999999999e-05 0 5.6019999999999996e-05 3.3 5.5939999999999996e-05 3.3 5.604e-05 0 5.596e-05 0 5.606e-05 3.3 5.5979999999999996e-05 3.3 5.608e-05 0 5.6e-05 0 5.61e-05 3.3 5.6019999999999996e-05 3.3 5.612e-05 0 5.604e-05 0 5.614e-05 3.3 5.6059999999999995e-05 3.3 5.616e-05 0 5.608e-05 0 5.618e-05 3.3 5.6099999999999995e-05 3.3 5.62e-05 0 5.612e-05 0 5.622e-05 3.3 5.6139999999999994e-05 3.3 5.624e-05 0 5.616e-05 0 5.626e-05 3.3 5.6179999999999994e-05 3.3 5.6279999999999996e-05 0 5.62e-05 0 5.63e-05 3.3 5.6219999999999994e-05 3.3 5.6319999999999996e-05 0 5.624e-05 0 5.634e-05 3.3 5.625999999999999e-05 3.3 5.6359999999999996e-05 0 5.6279999999999996e-05 0 5.638e-05 3.3 5.63e-05 3.3 5.64e-05 0 5.6319999999999996e-05 0 5.642e-05 3.3 5.634e-05 3.3 5.644e-05 0 5.6359999999999996e-05 0 5.646e-05 3.3 5.638e-05 3.3 5.648e-05 0 5.6399999999999995e-05 0 5.65e-05 3.3 5.642e-05 3.3 5.652e-05 0 5.6439999999999995e-05 0 5.654e-05 3.3 5.646e-05 3.3 5.656e-05 0 5.6479999999999995e-05 0 5.658e-05 3.3 5.65e-05 3.3 5.66e-05 0 5.6519999999999994e-05 0 5.662e-05 3.3 5.654e-05 3.3 5.664e-05 0 5.6559999999999994e-05 0 5.6659999999999996e-05 3.3 5.658e-05 3.3 5.668e-05 0 5.6599999999999993e-05 0 5.6699999999999996e-05 3.3 5.662e-05 3.3 5.672e-05 0 5.664e-05 0 5.674e-05 3.3 5.6659999999999996e-05 3.3 5.676e-05 0 5.668e-05 0 5.678e-05 3.3 5.6699999999999996e-05 3.3 5.68e-05 0 5.672e-05 0 5.682e-05 3.3 5.6739999999999995e-05 3.3 5.684e-05 0 5.676e-05 0 5.686e-05 3.3 5.6779999999999995e-05 3.3 5.688e-05 0 5.68e-05 0 5.69e-05 3.3 5.6819999999999995e-05 3.3 5.692e-05 0 5.684e-05 0 5.694e-05 3.3 5.6859999999999994e-05 3.3 5.696e-05 0 5.688e-05 0 5.698e-05 3.3 5.6899999999999994e-05 3.3 5.6999999999999996e-05 0 5.692e-05 0 5.702e-05 3.3 5.6939999999999994e-05 3.3 5.7039999999999996e-05 0 5.696e-05 0 5.706e-05 3.3 5.697999999999999e-05 3.3 5.7079999999999996e-05 0 5.6999999999999996e-05 0 5.71e-05 3.3 5.702e-05 3.3 5.712e-05 0 5.7039999999999996e-05 0 5.714e-05 3.3 5.706e-05 3.3 5.716e-05 0 5.7079999999999996e-05 0 5.718e-05 3.3 5.71e-05 3.3 5.72e-05 0 5.7119999999999995e-05 0 5.722e-05 3.3 5.714e-05 3.3 5.724e-05 0 5.7159999999999995e-05 0 5.726e-05 3.3 5.718e-05 3.3 5.728e-05 0 5.7199999999999994e-05 0 5.73e-05 3.3 5.722e-05 3.3 5.732e-05 0 5.7239999999999994e-05 0 5.7339999999999996e-05 3.3 5.726e-05 3.3 5.736e-05 0 5.7279999999999994e-05 0 5.7379999999999996e-05 3.3 5.73e-05 3.3 5.74e-05 0 5.731999999999999e-05 0 5.7419999999999996e-05 3.3 5.7339999999999996e-05 3.3 5.744e-05 0 5.736e-05 0 5.746e-05 3.3 5.7379999999999996e-05 3.3 5.748e-05 0 5.74e-05 0 5.75e-05 3.3 5.7419999999999996e-05 3.3 5.752e-05 0 5.744e-05 0 5.754e-05 3.3 5.7459999999999995e-05 3.3 5.756e-05 0 5.748e-05 0 5.758e-05 3.3 5.7499999999999995e-05 3.3 5.76e-05 0 5.752e-05 0 5.762e-05 3.3 5.7539999999999995e-05 3.3 5.764e-05 0 5.756e-05 0 5.766e-05 3.3 5.7579999999999994e-05 3.3 5.768e-05 0 5.76e-05 0 5.77e-05 3.3 5.7619999999999994e-05 3.3 5.7719999999999996e-05 0 5.764e-05 0 5.774e-05 3.3 5.7659999999999993e-05 3.3 5.7759999999999996e-05 0 5.768e-05 0 5.778e-05 3.3 5.769999999999999e-05 3.3 5.7799999999999995e-05 0 5.7719999999999996e-05 0 5.782e-05 3.3 5.774e-05 3.3 5.784e-05 0 5.7759999999999996e-05 0 5.786e-05 3.3 5.778e-05 3.3 5.788e-05 0 5.7799999999999995e-05 0 5.79e-05 3.3 5.782e-05 3.3 5.792e-05 0 5.7839999999999995e-05 0 5.794e-05 3.3 5.786e-05 3.3 5.796e-05 0 5.7879999999999995e-05 0 5.798e-05 3.3 5.79e-05 3.3 5.8e-05 0 5.7919999999999994e-05 0 5.802e-05 3.3 5.794e-05 3.3 5.804e-05 0 5.7959999999999994e-05 0 5.8059999999999996e-05 3.3 5.798e-05 3.3 5.808e-05 0 5.7999999999999994e-05 0 5.8099999999999996e-05 3.3 5.802e-05 3.3 5.812e-05 0 5.803999999999999e-05 0 5.8139999999999996e-05 3.3 5.8059999999999996e-05 3.3 5.816e-05 0 5.808e-05 0 5.818e-05 3.3 5.8099999999999996e-05 3.3 5.82e-05 0 5.812e-05 0 5.822e-05 3.3 5.8139999999999996e-05 3.3 5.824e-05 0 5.816e-05 0 5.826e-05 3.3 5.8179999999999995e-05 3.3 5.828e-05 0 5.82e-05 0 5.83e-05 3.3 5.8219999999999995e-05 3.3 5.832e-05 0 5.824e-05 0 5.834e-05 3.3 5.8259999999999994e-05 3.3 5.836e-05 0 5.828e-05 0 5.838e-05 3.3 5.8299999999999994e-05 3.3 5.8399999999999997e-05 0 5.832e-05 0 5.842e-05 3.3 5.8339999999999994e-05 3.3 5.8439999999999996e-05 0 5.836e-05 0 5.846e-05 3.3 5.837999999999999e-05 3.3 5.8479999999999996e-05 0 5.8399999999999997e-05 0 5.85e-05 3.3 5.842e-05 3.3 5.852e-05 0 5.8439999999999996e-05 0 5.854e-05 3.3 5.846e-05 3.3 5.856e-05 0 5.8479999999999996e-05 0 5.858e-05 3.3 5.85e-05 3.3 5.86e-05 0 5.8519999999999995e-05 0 5.862e-05 3.3 5.854e-05 3.3 5.864e-05 0 5.8559999999999995e-05 0 5.866e-05 3.3 5.858e-05 3.3 5.868e-05 0 5.8599999999999995e-05 0 5.87e-05 3.3 5.862e-05 3.3 5.872e-05 0 5.8639999999999994e-05 0 5.874e-05 3.3 5.866e-05 3.3 5.876e-05 0 5.8679999999999994e-05 0 5.8779999999999996e-05 3.3 5.87e-05 3.3 5.88e-05 0 5.8719999999999993e-05 0 5.8819999999999996e-05 3.3 5.874e-05 3.3 5.884e-05 0 5.875999999999999e-05 0 5.8859999999999995e-05 3.3 5.8779999999999996e-05 3.3 5.888e-05 0 5.88e-05 0 5.89e-05 3.3 5.8819999999999996e-05 3.3 5.892e-05 0 5.884e-05 0 5.894e-05 3.3 5.8859999999999995e-05 3.3 5.896e-05 0 5.888e-05 0 5.898e-05 3.3 5.8899999999999995e-05 3.3 5.9e-05 0 5.892e-05 0 5.902e-05 3.3 5.8939999999999995e-05 3.3 5.904e-05 0 5.896e-05 0 5.906e-05 3.3 5.8979999999999994e-05 3.3 5.908e-05 0 5.9e-05 0 5.91e-05 3.3 5.9019999999999994e-05 3.3 5.9119999999999996e-05 0 5.904e-05 0 5.914e-05 3.3 5.9059999999999994e-05 3.3 5.9159999999999996e-05 0 5.908e-05 0 5.918e-05 3.3 5.909999999999999e-05 3.3 5.9199999999999996e-05 0 5.9119999999999996e-05 0 5.922e-05 3.3 5.914e-05 3.3 5.924e-05 0 5.9159999999999996e-05 0 5.926e-05 3.3 5.918e-05 3.3 5.928e-05 0 5.9199999999999996e-05 0 5.93e-05 3.3 5.922e-05 3.3 5.932e-05 0 5.9239999999999995e-05 0 5.934e-05 3.3 5.926e-05 3.3 5.936e-05 0 5.9279999999999995e-05 0 5.938e-05 3.3 5.93e-05 3.3 5.94e-05 0 5.9319999999999994e-05 0 5.942e-05 3.3 5.934e-05 3.3 5.944e-05 0 5.9359999999999994e-05 0 5.9459999999999997e-05 3.3 5.938e-05 3.3 5.948e-05 0 5.9399999999999994e-05 0 5.9499999999999996e-05 3.3 5.942e-05 3.3 5.952e-05 0 5.943999999999999e-05 0 5.9539999999999996e-05 3.3 5.9459999999999997e-05 3.3 5.956e-05 0 5.948e-05 0 5.958e-05 3.3 5.9499999999999996e-05 3.3 5.96e-05 0 5.952e-05 0 5.962e-05 3.3 5.9539999999999996e-05 3.3 5.964e-05 0 5.956e-05 0 5.966e-05 3.3 5.9579999999999995e-05 3.3 5.968e-05 0 5.96e-05 0 5.97e-05 3.3 5.9619999999999995e-05 3.3 5.972e-05 0 5.964e-05 0 5.974e-05 3.3 5.9659999999999995e-05 3.3 5.976e-05 0 5.968e-05 0 5.978e-05 3.3 5.9699999999999994e-05 3.3 5.98e-05 0 5.972e-05 0 5.982e-05 3.3 5.9739999999999994e-05 3.3 5.9839999999999996e-05 0 5.976e-05 0 5.986e-05 3.3 5.9779999999999993e-05 3.3 5.9879999999999996e-05 0 5.98e-05 0 5.99e-05 3.3 5.981999999999999e-05 3.3 5.9919999999999996e-05 0 5.9839999999999996e-05 0 5.994e-05 3.3 5.986e-05 3.3 5.996e-05 0 5.9879999999999996e-05 0 5.998e-05 3.3 5.99e-05 3.3 6e-05 0 5.9919999999999996e-05 0 6.002e-05 3.3 5.994e-05 3.3 6.004e-05 0 5.9959999999999995e-05 0 6.006e-05 3.3 5.998e-05 3.3 6.008e-05 0 5.9999999999999995e-05 0 6.01e-05 3.3 6.002e-05 3.3 6.012e-05 0 6.0039999999999994e-05 0 6.014e-05 3.3 6.006e-05 3.3 6.016e-05 0 6.0079999999999994e-05 0 6.0179999999999996e-05 3.3 6.01e-05 3.3 6.02e-05 0 6.0119999999999994e-05 0 6.0219999999999996e-05 3.3 6.014e-05 3.3 6.024e-05 0 6.015999999999999e-05 0 6.0259999999999996e-05 3.3 6.0179999999999996e-05 3.3 6.028e-05 0 6.02e-05 0 6.03e-05 3.3 6.0219999999999996e-05 3.3 6.032e-05 0 6.024e-05 0 6.034e-05 3.3 6.0259999999999996e-05 3.3 6.036e-05 0 6.028e-05 0 6.038e-05 3.3 6.0299999999999995e-05 3.3 6.04e-05 0 6.032e-05 0 6.042e-05 3.3 6.0339999999999995e-05 3.3 6.044e-05 0 6.036e-05 0 6.046e-05 3.3 6.0379999999999994e-05 3.3 6.048e-05 0 6.04e-05 0 6.05e-05 3.3 6.0419999999999994e-05 3.3 6.0519999999999997e-05 0 6.044e-05 0 6.054e-05 3.3 6.0459999999999994e-05 3.3 6.0559999999999996e-05 0 6.048e-05 0 6.058e-05 3.3 6.049999999999999e-05 3.3 6.0599999999999996e-05 0 6.0519999999999997e-05 0 6.062e-05 3.3 6.053999999999999e-05 3.3 6.0639999999999995e-05 0 6.0559999999999996e-05 0 6.066e-05 3.3 6.058e-05 3.3 6.068e-05 0 6.0599999999999996e-05 0 6.07e-05 3.3 6.062e-05 3.3 6.072e-05 0 6.0639999999999995e-05 0 6.074e-05 3.3 6.066e-05 3.3 6.076e-05 0 6.0679999999999995e-05 0 6.078e-05 3.3 6.07e-05 3.3 6.08e-05 0 6.0719999999999995e-05 0 6.082e-05 3.3 6.074e-05 3.3 6.084e-05 0 6.0759999999999994e-05 0 6.086e-05 3.3 6.078e-05 3.3 6.088e-05 0 6.0799999999999994e-05 0 6.0899999999999996e-05 3.3 6.082e-05 3.3 6.092e-05 0 6.0839999999999993e-05 0 6.0939999999999996e-05 3.3 6.086e-05 3.3 6.096e-05 0 6.087999999999999e-05 0 6.0979999999999996e-05 3.3 6.0899999999999996e-05 3.3 6.1e-05 0 6.092e-05 0 6.102e-05 3.3 6.0939999999999996e-05 3.3 6.104e-05 0 6.096e-05 0 6.106e-05 3.3 6.098e-05 3.3 6.108e-05 0 6.099999999999999e-05 0 6.11e-05 3.3 6.1019999999999995e-05 3.3 6.112e-05 0 6.104e-05 0 6.114e-05 3.3 6.106e-05 3.3 6.116e-05 0 6.107999999999999e-05 0 6.118e-05 3.3 6.11e-05 3.3 6.12e-05 0 6.112e-05 0 6.122e-05 3.3 6.114e-05 3.3 6.124e-05 0 6.115999999999999e-05 0 6.125999999999999e-05 3.3 6.118e-05 3.3 6.128e-05 0 6.12e-05 0 6.13e-05 3.3 6.122e-05 3.3 6.132e-05 0 6.123999999999999e-05 0 6.133999999999999e-05 3.3 6.125999999999999e-05 3.3 6.136e-05 0 6.128e-05 0 6.138e-05 3.3 6.13e-05 3.3 6.14e-05 0 6.132e-05 0 6.142e-05 3.3 6.133999999999999e-05 3.3 6.144e-05 0 6.136e-05 0 6.146e-05 3.3 6.138e-05 3.3 6.148e-05 0 6.14e-05 0 6.15e-05 3.3 6.141999999999999e-05 3.3 6.152e-05 0 6.144e-05 0 6.154e-05 3.3 6.146e-05 3.3 6.156e-05 0 6.148e-05 0 6.158e-05 3.3 6.149999999999999e-05 3.3 6.159999999999999e-05 0 6.152e-05 0 6.162e-05 3.3 6.154e-05 3.3 6.164e-05 0 6.156e-05 0 6.166e-05 3.3 6.157999999999999e-05 3.3 6.167999999999999e-05 0 6.159999999999999e-05 0 6.17e-05 3.3 6.162e-05 3.3 6.172e-05 0 6.164e-05 0 6.174e-05 3.3 6.166e-05 3.3 6.176e-05 0 6.167999999999999e-05 0 6.178e-05 3.3 6.17e-05 3.3 6.18e-05 0 6.172e-05 0 6.182e-05 3.3 6.174e-05 3.3 6.184e-05 0 6.175999999999999e-05 0 6.186e-05 3.3 6.178e-05 3.3 6.188e-05 0 6.18e-05 0 6.19e-05 3.3 6.182e-05 3.3 6.192e-05 0 6.183999999999999e-05 0 6.193999999999999e-05 3.3 6.186e-05 3.3 6.196e-05 0 6.188e-05 0 6.198e-05 3.3 6.19e-05 3.3 6.2e-05 0 6.191999999999999e-05 0 6.201999999999999e-05 3.3 6.193999999999999e-05 3.3 6.204e-05 0 6.196e-05 0 6.206e-05 3.3 6.198e-05 3.3 6.208e-05 0 6.2e-05 0 6.21e-05 3.3 6.201999999999999e-05 3.3 6.212e-05 0 6.204e-05 0 6.214e-05 3.3 6.206e-05 3.3 6.216e-05 0 6.208e-05 0 6.218e-05 3.3 6.209999999999999e-05 3.3 6.22e-05 0 6.212e-05 0 6.222e-05 3.3 6.214e-05 3.3 6.224e-05 0 6.216e-05 0 6.226e-05 3.3 6.217999999999999e-05 3.3 6.228e-05 0 6.22e-05 0 6.23e-05 3.3 6.222e-05 3.3 6.232e-05 0 6.224e-05 0 6.234e-05 3.3 6.225999999999999e-05 3.3 6.235999999999999e-05 0 6.228e-05 0 6.238e-05 3.3 6.23e-05 3.3 6.24e-05 0 6.232e-05 0 6.242e-05 3.3 6.234e-05 3.3 6.244e-05 0 6.235999999999999e-05 0 6.246e-05 3.3 6.238e-05 3.3 6.248e-05 0 6.24e-05 0 6.25e-05 3.3 6.242e-05 3.3 6.252e-05 0 6.243999999999999e-05 0 6.254e-05 3.3 6.246e-05 3.3 6.256e-05 0 6.248e-05 0 6.258e-05 3.3 6.25e-05 3.3 6.26e-05 0 6.251999999999999e-05 0 6.262e-05 3.3 6.254e-05 3.3 6.264e-05 0 6.256e-05 0 6.266e-05 3.3 6.258e-05 3.3 6.268e-05 0 6.259999999999999e-05 0 6.269999999999999e-05 3.3 6.262e-05 3.3 6.272e-05 0 6.264e-05 0 6.274e-05 3.3 6.266e-05 3.3 6.276e-05 0 6.268e-05 0 6.278e-05 3.3 6.269999999999999e-05 3.3 6.28e-05 0 6.272e-05 0 6.282e-05 3.3 6.274e-05 3.3 6.284e-05 0 6.276e-05 0 6.286e-05 3.3 6.277999999999999e-05 3.3 6.288e-05 0 6.28e-05 0 6.29e-05 3.3 6.282e-05 3.3 6.292e-05 0 6.284e-05 0 6.294e-05 3.3 6.285999999999999e-05 3.3 6.296e-05 0 6.288e-05 0 6.298e-05 3.3 6.29e-05 3.3 6.3e-05 0 6.292e-05 0 6.302e-05 3.3 6.293999999999999e-05 3.3 6.303999999999999e-05 0 6.296e-05 0 6.306e-05 3.3 6.298e-05 3.3 6.308e-05 0 6.3e-05 0 6.31e-05 3.3 6.301999999999999e-05 3.3 6.311999999999999e-05 0 6.303999999999999e-05 0 6.314e-05 3.3 6.306e-05 3.3 6.316e-05 0 6.308e-05 0 6.318e-05 3.3 6.31e-05 3.3 6.32e-05 0 6.311999999999999e-05 0 6.322e-05 3.3 6.314e-05 3.3 6.324e-05 0 6.316e-05 0 6.326e-05 3.3 6.318e-05 3.3 6.328e-05 0 6.319999999999999e-05 0 6.33e-05 3.3 6.322e-05 3.3 6.332e-05 0 6.324e-05 0 6.334e-05 3.3 6.326e-05 3.3 6.336e-05 0 6.327999999999999e-05 0 6.337999999999999e-05 3.3 6.33e-05 3.3 6.34e-05 0 6.332e-05 0 6.342e-05 3.3 6.334e-05 3.3 6.344e-05 0 6.335999999999999e-05 0 6.345999999999999e-05 3.3 6.337999999999999e-05 3.3 6.348e-05 0 6.34e-05 0 6.35e-05 3.3 6.342e-05 3.3 6.352e-05 0 6.344e-05 0 6.354e-05 3.3 6.345999999999999e-05 3.3 6.356e-05 0 6.348e-05 0 6.358e-05 3.3 6.35e-05 3.3 6.36e-05 0 6.352e-05 0 6.362e-05 3.3 6.353999999999999e-05 3.3 6.364e-05 0 6.356e-05 0 6.366e-05 3.3 6.358e-05 3.3 6.368e-05 0 6.36e-05 0 6.37e-05 3.3 6.361999999999999e-05 3.3 6.371999999999999e-05 0 6.364e-05 0 6.374e-05 3.3 6.366e-05 3.3 6.376e-05 0 6.368e-05 0 6.378e-05 3.3 6.369999999999999e-05 3.3 6.379999999999999e-05 0 6.371999999999999e-05 0 6.382e-05 3.3 6.374e-05 3.3 6.384e-05 0 6.376e-05 0 6.386e-05 3.3 6.378e-05 3.3 6.388e-05 0 6.379999999999999e-05 0 6.39e-05 3.3 6.382e-05 3.3 6.392e-05 0 6.384e-05 0 6.394e-05 3.3 6.386e-05 3.3 6.396e-05 0 6.387999999999999e-05 0 6.398e-05 3.3 6.39e-05 3.3 6.4e-05 0 6.392e-05 0 6.402e-05 3.3 6.394e-05 3.3 6.404e-05 0 6.395999999999999e-05 0 6.405999999999999e-05 3.3 6.398e-05 3.3 6.408e-05 0 6.4e-05 0 6.41e-05 3.3 6.402e-05 3.3 6.412e-05 0 6.403999999999999e-05 0 6.413999999999999e-05 3.3 6.405999999999999e-05 3.3 6.416e-05 0 6.408e-05 0 6.418e-05 3.3 6.41e-05 3.3 6.42e-05 0 6.412e-05 0 6.422e-05 3.3 6.413999999999999e-05 3.3 6.424e-05 0 6.416e-05 0 6.426e-05 3.3 6.418e-05 3.3 6.428e-05 0 6.42e-05 0 6.43e-05 3.3 6.421999999999999e-05 3.3 6.432e-05 0 6.424e-05 0 6.434e-05 3.3 6.426e-05 3.3 6.436e-05 0 6.428e-05 0 6.438e-05 3.3 6.429999999999999e-05 3.3 6.44e-05 0 6.432e-05 0 6.442e-05 3.3 6.434e-05 3.3 6.444e-05 0 6.436e-05 0 6.446e-05 3.3 6.437999999999999e-05 3.3 6.447999999999999e-05 0 6.44e-05 0 6.45e-05 3.3 6.442e-05 3.3 6.452e-05 0 6.444e-05 0 6.454e-05 3.3 6.446e-05 3.3 6.456e-05 0 6.447999999999999e-05 0 6.458e-05 3.3 6.45e-05 3.3 6.46e-05 0 6.452e-05 0 6.462e-05 3.3 6.454e-05 3.3 6.464e-05 0 6.455999999999999e-05 0 6.466e-05 3.3 6.458e-05 3.3 6.468e-05 0 6.46e-05 0 6.47e-05 3.3 6.462e-05 3.3 6.472e-05 0 6.463999999999999e-05 0 6.474e-05 3.3 6.466e-05 3.3 6.476e-05 0 6.468e-05 0 6.478e-05 3.3 6.47e-05 3.3 6.48e-05 0 6.471999999999999e-05 0 6.481999999999999e-05 3.3 6.474e-05 3.3 6.484e-05 0 6.476e-05 0 6.486e-05 3.3 6.478e-05 3.3 6.488e-05 0 6.48e-05 0 6.49e-05 3.3 6.481999999999999e-05 3.3 6.492e-05 0 6.484e-05 0 6.494e-05 3.3 6.486e-05 3.3 6.496e-05 0 6.488e-05 0 6.498e-05 3.3 6.489999999999999e-05 3.3 6.5e-05 0 6.492e-05 0 6.502e-05 3.3 6.494e-05 3.3 6.504e-05 0 6.496e-05 0 6.506e-05 3.3 6.497999999999999e-05 3.3 6.508e-05 0 6.5e-05 0 6.51e-05 3.3 6.502e-05 3.3 6.512e-05 0 6.504e-05 0 6.514e-05 3.3 6.505999999999999e-05 3.3 6.515999999999999e-05 0 6.508e-05 0 6.518e-05 3.3 6.51e-05 3.3 6.52e-05 0 6.512e-05 0 6.522e-05 3.3 6.513999999999999e-05 3.3 6.523999999999999e-05 0 6.515999999999999e-05 0 6.526e-05 3.3 6.518e-05 3.3 6.528e-05 0 6.52e-05 0 6.53e-05 3.3 6.522e-05 3.3 6.532e-05 0 6.523999999999999e-05 0 6.534e-05 3.3 6.526e-05 3.3 6.536e-05 0 6.528e-05 0 6.538e-05 3.3 6.53e-05 3.3 6.54e-05 0 6.531999999999999e-05 0 6.542e-05 3.3 6.534e-05 3.3 6.544e-05 0 6.536e-05 0 6.546e-05 3.3 6.538e-05 3.3 6.548e-05 0 6.539999999999999e-05 0 6.549999999999999e-05 3.3 6.542e-05 3.3 6.552e-05 0 6.544e-05 0 6.554e-05 3.3 6.546e-05 3.3 6.556e-05 0 6.547999999999999e-05 0 6.557999999999999e-05 3.3 6.549999999999999e-05 3.3 6.56e-05 0 6.552e-05 0 6.562e-05 3.3 6.554e-05 3.3 6.564e-05 0 6.556e-05 0 6.566e-05 3.3 6.557999999999999e-05 3.3 6.568e-05 0 6.56e-05 0 6.57e-05 3.3 6.562e-05 3.3 6.572e-05 0 6.564e-05 0 6.574e-05 3.3 6.565999999999999e-05 3.3 6.576e-05 0 6.568e-05 0 6.578e-05 3.3 6.57e-05 3.3 6.58e-05 0 6.572e-05 0 6.582e-05 3.3 6.573999999999999e-05 3.3 6.583999999999999e-05 0 6.576e-05 0 6.586e-05 3.3 6.578e-05 3.3 6.588e-05 0 6.58e-05 0 6.59e-05 3.3 6.581999999999999e-05 3.3 6.591999999999999e-05 0 6.583999999999999e-05 0 6.594e-05 3.3 6.586e-05 3.3 6.596e-05 0 6.588e-05 0 6.598e-05 3.3 6.59e-05 3.3 6.6e-05 0 6.591999999999999e-05 0 6.602e-05 3.3 6.594e-05 3.3 6.604e-05 0 6.596e-05 0 6.606e-05 3.3 6.598e-05 3.3 6.608e-05 0 6.599999999999999e-05 0 6.61e-05 3.3 6.602e-05 3.3 6.612e-05 0 6.604e-05 0 6.614e-05 3.3 6.606e-05 3.3 6.616e-05 0 6.607999999999999e-05 0 6.617999999999999e-05 3.3 6.61e-05 3.3 6.62e-05 0 6.612e-05 0 6.622e-05 3.3 6.614e-05 3.3 6.624e-05 0 6.615999999999999e-05 0 6.625999999999999e-05 3.3 6.617999999999999e-05 3.3 6.628e-05 0 6.62e-05 0 6.63e-05 3.3 6.622e-05 3.3 6.632e-05 0 6.624e-05 0 6.634e-05 3.3 6.625999999999999e-05 3.3 6.636e-05 0 6.628e-05 0 6.638e-05 3.3 6.63e-05 3.3 6.64e-05 0 6.632e-05 0 6.642e-05 3.3 6.633999999999999e-05 3.3 6.644e-05 0 6.636e-05 0 6.646e-05 3.3 6.638e-05 3.3 6.648e-05 0 6.64e-05 0 6.65e-05 3.3 6.641999999999999e-05 3.3 6.652e-05 0 6.644e-05 0 6.654e-05 3.3 6.646e-05 3.3 6.656e-05 0 6.648e-05 0 6.658e-05 3.3 6.649999999999999e-05 3.3 6.659999999999999e-05 0 6.652e-05 0 6.662e-05 3.3 6.654e-05 3.3 6.664e-05 0 6.656e-05 0 6.666e-05 3.3 6.658e-05 3.3 6.668e-05 0 6.659999999999999e-05 0 6.67e-05 3.3 6.662e-05 3.3 6.672e-05 0 6.664e-05 0 6.674e-05 3.3 6.666e-05 3.3 6.676e-05 0 6.667999999999999e-05 0 6.678e-05 3.3 6.67e-05 3.3 6.68e-05 0 6.672e-05 0 6.682e-05 3.3 6.674e-05 3.3 6.684e-05 0 6.675999999999999e-05 0 6.686e-05 3.3 6.678e-05 3.3 6.688e-05 0 6.68e-05 0 6.69e-05 3.3 6.682e-05 3.3 6.692e-05 0 6.683999999999999e-05 0 6.693999999999999e-05 3.3 6.686e-05 3.3 6.696e-05 0 6.688e-05 0 6.698e-05 3.3 6.69e-05 3.3 6.7e-05 0 6.691999999999999e-05 0 6.701999999999999e-05 3.3 6.693999999999999e-05 3.3 6.704e-05 0 6.696e-05 0 6.706e-05 3.3 6.698e-05 3.3 6.708e-05 0 6.7e-05 0 6.71e-05 3.3 6.701999999999999e-05 3.3 6.712e-05 0 6.704e-05 0 6.714e-05 3.3 6.706e-05 3.3 6.716e-05 0 6.708e-05 0 6.718e-05 3.3 6.709999999999999e-05 3.3 6.72e-05 0 6.712e-05 0 6.722e-05 3.3 6.714e-05 3.3 6.724e-05 0 6.716e-05 0 6.726e-05 3.3 6.717999999999999e-05 3.3 6.727999999999999e-05 0 6.72e-05 0 6.73e-05 3.3 6.722e-05 3.3 6.732e-05 0 6.724e-05 0 6.734e-05 3.3 6.725999999999999e-05 3.3 6.735999999999999e-05 0 6.727999999999999e-05 0 6.738e-05 3.3 6.73e-05 3.3 6.74e-05 0 6.732e-05 0 6.742e-05 3.3 6.734e-05 3.3 6.744e-05 0 6.735999999999999e-05 0 6.746e-05 3.3 6.738e-05 3.3 6.748e-05 0 6.74e-05 0 6.75e-05 3.3 6.742e-05 3.3 6.752e-05 0 6.743999999999999e-05 0 6.754e-05 3.3 6.746e-05 3.3 6.756e-05 0 6.748e-05 0 6.758e-05 3.3 6.75e-05 3.3 6.76e-05 0 6.751999999999999e-05 0 6.761999999999999e-05 3.3 6.754e-05 3.3 6.764e-05 0 6.756e-05 0 6.766e-05 3.3 6.758e-05 3.3 6.768e-05 0 6.759999999999999e-05 0 6.769999999999999e-05 3.3 6.761999999999999e-05 3.3 6.772e-05 0 6.764e-05 0 6.774e-05 3.3 6.766e-05 3.3 6.776e-05 0 6.768e-05 0 6.778e-05 3.3 6.769999999999999e-05 3.3 6.78e-05 0 6.772e-05 0 6.782e-05 3.3 6.774e-05 3.3 6.784e-05 0 6.776e-05 0 6.786e-05 3.3 6.777999999999999e-05 3.3 6.788e-05 0 6.78e-05 0 6.79e-05 3.3 6.782e-05 3.3 6.792e-05 0 6.784e-05 0 6.794e-05 3.3 6.785999999999999e-05 3.3 6.795999999999999e-05 0 6.788e-05 0 6.798e-05 3.3 6.79e-05 3.3 6.8e-05 0 6.792e-05 0 6.802e-05 3.3 6.793999999999999e-05 3.3 6.803999999999999e-05 0 6.795999999999999e-05 0 6.806e-05 3.3 6.798e-05 3.3 6.808e-05 0 6.8e-05 0 6.81e-05 3.3 6.802e-05 3.3 6.812e-05 0 6.803999999999999e-05 0 6.814e-05 3.3 6.806e-05 3.3 6.816e-05 0 6.808e-05 0 6.818e-05 3.3 6.81e-05 3.3 6.82e-05 0 6.811999999999999e-05 0 6.822e-05 3.3 6.814e-05 3.3 6.824e-05 0 6.816e-05 0 6.826e-05 3.3 6.818e-05 3.3 6.828e-05 0 6.819999999999999e-05 0 6.829999999999999e-05 3.3 6.822e-05 3.3 6.832e-05 0 6.824e-05 0 6.834e-05 3.3 6.826e-05 3.3 6.836e-05 0 6.827999999999999e-05 0 6.837999999999999e-05 3.3 6.829999999999999e-05 3.3 6.84e-05 0 6.832e-05 0 6.842e-05 3.3 6.834e-05 3.3 6.844e-05 0 6.836e-05 0 6.846e-05 3.3 6.837999999999999e-05 3.3 6.848e-05 0 6.84e-05 0 6.85e-05 3.3 6.842e-05 3.3 6.852e-05 0 6.844e-05 0 6.854e-05 3.3 6.845999999999999e-05 3.3 6.856e-05 0 6.848e-05 0 6.858e-05 3.3 6.85e-05 3.3 6.86e-05 0 6.852e-05 0 6.862e-05 3.3 6.853999999999999e-05 3.3 6.864e-05 0 6.856e-05 0 6.866e-05 3.3 6.858e-05 3.3 6.868e-05 0 6.86e-05 0 6.87e-05 3.3 6.861999999999999e-05 3.3 6.871999999999999e-05 0 6.864e-05 0 6.874e-05 3.3 6.866e-05 3.3 6.876e-05 0 6.868e-05 0 6.878e-05 3.3 6.87e-05 3.3 6.88e-05 0 6.871999999999999e-05 0 6.882e-05 3.3 6.874e-05 3.3 6.884e-05 0 6.876e-05 0 6.886e-05 3.3 6.878e-05 3.3 6.888e-05 0 6.879999999999999e-05 0 6.89e-05 3.3 6.882e-05 3.3 6.892e-05 0 6.884e-05 0 6.894e-05 3.3 6.886e-05 3.3 6.896e-05 0 6.887999999999999e-05 0 6.898e-05 3.3 6.89e-05 3.3 6.9e-05 0 6.892e-05 0 6.902e-05 3.3 6.894e-05 3.3 6.904e-05 0 6.895999999999999e-05 0 6.905999999999999e-05 3.3 6.898e-05 3.3 6.908e-05 0 6.9e-05 0 6.91e-05 3.3 6.902e-05 3.3 6.912e-05 0 6.903999999999999e-05 0 6.913999999999999e-05 3.3 6.905999999999999e-05 3.3 6.916e-05 0 6.908e-05 0 6.918e-05 3.3 6.91e-05 3.3 6.92e-05 0 6.912e-05 0 6.922e-05 3.3 6.913999999999999e-05 3.3 6.924e-05 0 6.916e-05 0 6.926e-05 3.3 6.918e-05 3.3 6.928e-05 0 6.92e-05 0 6.93e-05 3.3 6.921999999999999e-05 3.3 6.932e-05 0 6.924e-05 0 6.934e-05 3.3 6.926e-05 3.3 6.936e-05 0 6.928e-05 0 6.938e-05 3.3 6.929999999999999e-05 3.3 6.939999999999999e-05 0 6.932e-05 0 6.942e-05 3.3 6.934e-05 3.3 6.944e-05 0 6.936e-05 0 6.946e-05 3.3 6.937999999999999e-05 3.3 6.947999999999999e-05 0 6.939999999999999e-05 0 6.95e-05 3.3 6.942e-05 3.3 6.952e-05 0 6.944e-05 0 6.954e-05 3.3 6.946e-05 3.3 6.956e-05 0 6.947999999999999e-05 0 6.958e-05 3.3 6.95e-05 3.3 6.96e-05 0 6.952e-05 0 6.962e-05 3.3 6.954e-05 3.3 6.964e-05 0 6.955999999999999e-05 0 6.966e-05 3.3 6.958e-05 3.3 6.968e-05 0 6.96e-05 0 6.97e-05 3.3 6.962e-05 3.3 6.972e-05 0 6.963999999999999e-05 0 6.973999999999999e-05 3.3 6.966e-05 3.3 6.976e-05 0 6.968e-05 0 6.978e-05 3.3 6.97e-05 3.3 6.98e-05 0 6.971999999999999e-05 0 6.981999999999999e-05 3.3 6.973999999999999e-05 3.3 6.984e-05 0 6.976e-05 0 6.986e-05 3.3 6.978e-05 3.3 6.988e-05 0 6.98e-05 0 6.99e-05 3.3 6.981999999999999e-05 3.3 6.992e-05 0 6.984e-05 0 6.994e-05 3.3 6.986e-05 3.3 6.996e-05 0 6.988e-05 0 6.998e-05 3.3 6.989999999999999e-05 3.3 7e-05 0 6.992e-05 0 7.002e-05 3.3 6.994e-05 3.3 7.004e-05 0 6.996e-05 0 7.006e-05 3.3 6.997999999999999e-05 3.3 7.007999999999999e-05 0 7e-05 0 7.01e-05 3.3 7.002e-05 3.3 7.012e-05 0 7.004e-05 0 7.014e-05 3.3 7.005999999999999e-05 3.3 7.015999999999999e-05 0 7.007999999999999e-05 0 7.018e-05 3.3 7.01e-05 3.3 7.02e-05 0 7.012e-05 0 7.022e-05 3.3 7.014e-05 3.3 7.024e-05 0 7.015999999999999e-05 0 7.026e-05 3.3 7.018e-05 3.3 7.028e-05 0 7.02e-05 0 7.03e-05 3.3 7.022e-05 3.3 7.032e-05 0 7.023999999999999e-05 0 7.034e-05 3.3 7.026e-05 3.3 7.036e-05 0 7.028e-05 0 7.038e-05 3.3 7.03e-05 3.3 7.04e-05 0 7.031999999999999e-05 0 7.042e-05 3.3 7.034e-05 3.3 7.044e-05 0 7.036e-05 0 7.046e-05 3.3 7.038e-05 3.3 7.048e-05 0 7.039999999999999e-05 0 7.049999999999999e-05 3.3 7.042e-05 3.3 7.052e-05 0 7.044e-05 0 7.054e-05 3.3 7.046e-05 3.3 7.056e-05 0 7.048e-05 0 7.058e-05 3.3 7.049999999999999e-05 3.3 7.06e-05 0 7.052e-05 0 7.062e-05 3.3 7.054e-05 3.3 7.064e-05 0 7.056e-05 0 7.066e-05 3.3 7.057999999999999e-05 3.3 7.068e-05 0 7.06e-05 0 7.07e-05 3.3 7.062e-05 3.3 7.072e-05 0 7.064e-05 0 7.074e-05 3.3 7.065999999999999e-05 3.3 7.076e-05 0 7.068e-05 0 7.078e-05 3.3 7.07e-05 3.3 7.08e-05 0 7.072e-05 0 7.082e-05 3.3 7.073999999999999e-05 3.3 7.083999999999999e-05 0 7.076e-05 0 7.086e-05 3.3 7.078e-05 3.3 7.088e-05 0 7.08e-05 0 7.09e-05 3.3 7.081999999999999e-05 3.3 7.091999999999999e-05 0 7.083999999999999e-05 0 7.094e-05 3.3 7.086e-05 3.3 7.096e-05 0 7.088e-05 0 7.098e-05 3.3 7.09e-05 3.3 7.1e-05 0 7.091999999999999e-05 0 7.102e-05 3.3 7.094e-05 3.3 7.104e-05 0 7.096e-05 0 7.106e-05 3.3 7.098e-05 3.3 7.108e-05 0 7.099999999999999e-05 0 7.11e-05 3.3 7.102e-05 3.3 7.112e-05 0 7.104e-05 0 7.114e-05 3.3 7.106e-05 3.3 7.116e-05 0 7.107999999999999e-05 0 7.117999999999999e-05 3.3 7.11e-05 3.3 7.12e-05 0 7.112e-05 0 7.122e-05 3.3 7.114e-05 3.3 7.124e-05 0 7.115999999999999e-05 0 7.125999999999999e-05 3.3 7.117999999999999e-05 3.3 7.128e-05 0 7.12e-05 0 7.13e-05 3.3 7.122e-05 3.3 7.132e-05 0 7.124e-05 0 7.134e-05 3.3 7.125999999999999e-05 3.3 7.136e-05 0 7.128e-05 0 7.138e-05 3.3 7.13e-05 3.3 7.14e-05 0 7.132e-05 0 7.142e-05 3.3 7.133999999999999e-05 3.3 7.144e-05 0 7.136e-05 0 7.146e-05 3.3 7.138e-05 3.3 7.148e-05 0 7.14e-05 0 7.15e-05 3.3 7.141999999999999e-05 3.3 7.151999999999999e-05 0 7.144e-05 0 7.154e-05 3.3 7.146e-05 3.3 7.156e-05 0 7.148e-05 0 7.158e-05 3.3 7.149999999999999e-05 3.3 7.159999999999999e-05 0 7.151999999999999e-05 0 7.162e-05 3.3 7.154e-05 3.3 7.164e-05 0 7.156e-05 0 7.166e-05 3.3 7.158e-05 3.3 7.168e-05 0 7.159999999999999e-05 0 7.17e-05 3.3 7.162e-05 3.3 7.172e-05 0 7.164e-05 0 7.174e-05 3.3 7.166e-05 3.3 7.176e-05 0 7.167999999999999e-05 0 7.178e-05 3.3 7.17e-05 3.3 7.18e-05 0 7.172e-05 0 7.182e-05 3.3 7.174e-05 3.3 7.184e-05 0 7.175999999999999e-05 0 7.185999999999999e-05 3.3 7.178e-05 3.3 7.188e-05 0 7.18e-05 0 7.19e-05 3.3 7.182e-05 3.3 7.192e-05 0 7.183999999999999e-05 0 7.193999999999999e-05 3.3 7.185999999999999e-05 3.3 7.196e-05 0 7.188e-05 0 7.198e-05 3.3 7.19e-05 3.3 7.2e-05 0 7.192e-05 0 7.202e-05 3.3 7.193999999999999e-05 3.3 7.204e-05 0 7.196e-05 0 7.206e-05 3.3 7.198e-05 3.3 7.208e-05 0 7.2e-05 0 7.21e-05 3.3 7.201999999999999e-05 3.3 7.212e-05 0 7.204e-05 0 7.214e-05 3.3 7.206e-05 3.3 7.216e-05 0 7.208e-05 0 7.218e-05 3.3 7.209999999999999e-05 3.3 7.219999999999999e-05 0 7.212e-05 0 7.222e-05 3.3 7.214e-05 3.3 7.224e-05 0 7.216e-05 0 7.226e-05 3.3 7.217999999999999e-05 3.3 7.227999999999999e-05 0 7.219999999999999e-05 0 7.23e-05 3.3 7.222e-05 3.3 7.232e-05 0 7.224e-05 0 7.234e-05 3.3 7.226e-05 3.3 7.236e-05 0 7.227999999999999e-05 0 7.238e-05 3.3 7.23e-05 3.3 7.24e-05 0 7.232e-05 0 7.242e-05 3.3 7.234e-05 3.3 7.244e-05 0 7.235999999999999e-05 0 7.246e-05 3.3 7.238e-05 3.3 7.248e-05 0 7.24e-05 0 7.25e-05 3.3 7.242e-05 3.3 7.252e-05 0 7.243999999999999e-05 0 7.254e-05 3.3 7.246e-05 3.3 7.256e-05 0 7.248e-05 0 7.258e-05 3.3 7.25e-05 3.3 7.26e-05 0 7.251999999999999e-05 0 7.261999999999999e-05 3.3 7.254e-05 3.3 7.264e-05 0 7.256e-05 0 7.266e-05 3.3 7.258e-05 3.3 7.268e-05 0 7.26e-05 0 7.27e-05 3.3 7.261999999999999e-05 3.3 7.272e-05 0 7.264e-05 0 7.274e-05 3.3 7.266e-05 3.3 7.276e-05 0 7.268e-05 0 7.278e-05 3.3 7.269999999999999e-05 3.3 7.28e-05 0 7.272e-05 0 7.282e-05 3.3 7.274e-05 3.3 7.284e-05 0 7.276e-05 0 7.286e-05 3.3 7.277999999999999e-05 3.3 7.288e-05 0 7.28e-05 0 7.29e-05 3.3 7.282e-05 3.3 7.292e-05 0 7.284e-05 0 7.294e-05 3.3 7.285999999999999e-05 3.3 7.295999999999999e-05 0 7.288e-05 0 7.298e-05 3.3 7.29e-05 3.3 7.3e-05 0 7.292e-05 0 7.302e-05 3.3 7.293999999999999e-05 3.3 7.303999999999999e-05 0 7.295999999999999e-05 0 7.306e-05 3.3 7.298e-05 3.3 7.308e-05 0 7.3e-05 0 7.31e-05 3.3 7.302e-05 3.3 7.312e-05 0 7.303999999999999e-05 0 7.314e-05 3.3 7.306e-05 3.3 7.316e-05 0 7.308e-05 0 7.318e-05 3.3 7.31e-05 3.3 7.32e-05 0 7.311999999999999e-05 0 7.322e-05 3.3 7.314e-05 3.3 7.324e-05 0 7.316e-05 0 7.326e-05 3.3 7.318e-05 3.3 7.328e-05 0 7.319999999999999e-05 0 7.329999999999999e-05 3.3 7.322e-05 3.3 7.332e-05 0 7.324e-05 0 7.334e-05 3.3 7.326e-05 3.3 7.336e-05 0 7.327999999999999e-05 0 7.337999999999999e-05 3.3 7.329999999999999e-05 3.3 7.34e-05 0 7.332e-05 0 7.342e-05 3.3 7.334e-05 3.3 7.344e-05 0 7.336e-05 0 7.346e-05 3.3 7.337999999999999e-05 3.3 7.348e-05 0 7.34e-05 0 7.35e-05 3.3 7.342e-05 3.3 7.352e-05 0 7.344e-05 0 7.354e-05 3.3 7.345999999999999e-05 3.3 7.356e-05 0 7.348e-05 0 7.358e-05 3.3 7.35e-05 3.3 7.36e-05 0 7.352e-05 0 7.362e-05 3.3 7.353999999999999e-05 3.3 7.363999999999999e-05 0 7.356e-05 0 7.366e-05 3.3 7.358e-05 3.3 7.368e-05 0 7.36e-05 0 7.37e-05 3.3 7.361999999999999e-05 3.3 7.371999999999999e-05 0 7.363999999999999e-05 0 7.374e-05 3.3 7.366e-05 3.3 7.376e-05 0 7.368e-05 0 7.378e-05 3.3 7.37e-05 3.3 7.38e-05 0 7.371999999999999e-05 0 7.382e-05 3.3 7.374e-05 3.3 7.384e-05 0 7.376e-05 0 7.386e-05 3.3 7.378e-05 3.3 7.388e-05 0 7.379999999999999e-05 0 7.39e-05 3.3 7.382e-05 3.3 7.392e-05 0 7.384e-05 0 7.394e-05 3.3 7.386e-05 3.3 7.396e-05 0 7.387999999999999e-05 0 7.397999999999999e-05 3.3 7.39e-05 3.3 7.4e-05 0 7.392e-05 0 7.402e-05 3.3 7.394e-05 3.3 7.404e-05 0 7.395999999999999e-05 0 7.405999999999999e-05 3.3 7.397999999999999e-05 3.3 7.408e-05 0 7.4e-05 0 7.41e-05 3.3 7.402e-05 3.3 7.412e-05 0 7.404e-05 0 7.414e-05 3.3 7.405999999999999e-05 3.3 7.416e-05 0 7.408e-05 0 7.418e-05 3.3 7.41e-05 3.3 7.42e-05 0 7.412e-05 0 7.422e-05 3.3 7.413999999999999e-05 3.3 7.424e-05 0 7.416e-05 0 7.426e-05 3.3 7.418e-05 3.3 7.428e-05 0 7.42e-05 0 7.43e-05 3.3 7.421999999999999e-05 3.3 7.431999999999999e-05 0 7.424e-05 0 7.434e-05 3.3 7.426e-05 3.3 7.436e-05 0 7.428e-05 0 7.438e-05 3.3 7.429999999999999e-05 3.3 7.439999999999999e-05 0 7.431999999999999e-05 0 7.442e-05 3.3 7.434e-05 3.3 7.444e-05 0 7.436e-05 0 7.446e-05 3.3 7.438e-05 3.3 7.448e-05 0 7.439999999999999e-05 0 7.45e-05 3.3 7.442e-05 3.3 7.452e-05 0 7.444e-05 0 7.454e-05 3.3 7.446e-05 3.3 7.456e-05 0 7.447999999999999e-05 0 7.458e-05 3.3 7.45e-05 3.3 7.46e-05 0 7.452e-05 0 7.462e-05 3.3 7.454e-05 3.3 7.464e-05 0 7.455999999999999e-05 0 7.466e-05 3.3 7.458e-05 3.3 7.468e-05 0 7.46e-05 0 7.47e-05 3.3 7.462e-05 3.3 7.472e-05 0 7.463999999999999e-05 0 7.473999999999999e-05 3.3 7.466e-05 3.3 7.476e-05 0 7.468e-05 0 7.478e-05 3.3 7.47e-05 3.3 7.48e-05 0 7.471999999999999e-05 0 7.481999999999999e-05 3.3 7.473999999999999e-05 3.3 7.484e-05 0 7.476e-05 0 7.486e-05 3.3 7.478e-05 3.3 7.488e-05 0 7.48e-05 0 7.49e-05 3.3 7.481999999999999e-05 3.3 7.492e-05 0 7.484e-05 0 7.494e-05 3.3 7.486e-05 3.3 7.496e-05 0 7.488e-05 0 7.498e-05 3.3 7.489999999999999e-05 3.3 7.5e-05 0 7.492e-05 0 7.502e-05 3.3 7.494e-05 3.3 7.504e-05 0 7.496e-05 0 7.506e-05 3.3 7.497999999999999e-05 3.3 7.507999999999999e-05 0 7.5e-05 0 7.51e-05 3.3 7.502e-05 3.3 7.512e-05 0 7.504e-05 0 7.514e-05 3.3 7.505999999999999e-05 3.3 7.515999999999999e-05 0 7.507999999999999e-05 0 7.518e-05 3.3 7.51e-05 3.3 7.52e-05 0 7.512e-05 0 7.522e-05 3.3 7.514e-05 3.3 7.524e-05 0 7.515999999999999e-05 0 7.526e-05 3.3 7.518e-05 3.3 7.528e-05 0 7.52e-05 0 7.53e-05 3.3 7.522e-05 3.3 7.532e-05 0 7.523999999999999e-05 0 7.534e-05 3.3 7.526e-05 3.3 7.536e-05 0 7.528e-05 0 7.538e-05 3.3 7.53e-05 3.3 7.54e-05 0 7.531999999999999e-05 0 7.541999999999999e-05 3.3 7.534e-05 3.3 7.544e-05 0 7.536e-05 0 7.546e-05 3.3 7.538e-05 3.3 7.548e-05 0 7.539999999999999e-05 0 7.549999999999999e-05 3.3 7.541999999999999e-05 3.3 7.552e-05 0 7.544e-05 0 7.554e-05 3.3 7.546e-05 3.3 7.556e-05 0 7.548e-05 0 7.558e-05 3.3 7.549999999999999e-05 3.3 7.56e-05 0 7.552e-05 0 7.562e-05 3.3 7.554e-05 3.3 7.564e-05 0 7.556e-05 0 7.566e-05 3.3 7.557999999999999e-05 3.3 7.568e-05 0 7.56e-05 0 7.57e-05 3.3 7.562e-05 3.3 7.572e-05 0 7.564e-05 0 7.574e-05 3.3 7.565999999999999e-05 3.3 7.575999999999999e-05 0 7.568e-05 0 7.578e-05 3.3 7.57e-05 3.3 7.58e-05 0 7.572e-05 0 7.582e-05 3.3 7.573999999999999e-05 3.3 7.583999999999999e-05 0 7.575999999999999e-05 0 7.586e-05 3.3 7.578e-05 3.3 7.588e-05 0 7.58e-05 0 7.59e-05 3.3 7.582e-05 3.3 7.592e-05 0 7.583999999999999e-05 0 7.594e-05 3.3 7.586e-05 3.3 7.596e-05 0 7.588e-05 0 7.598e-05 3.3 7.59e-05 3.3 7.6e-05 0 7.591999999999999e-05 0 7.602e-05 3.3 7.594e-05 3.3 7.604e-05 0 7.596e-05 0 7.606e-05 3.3 7.598e-05 3.3 7.608e-05 0 7.599999999999999e-05 0 7.609999999999999e-05 3.3 7.602e-05 3.3 7.612e-05 0 7.604e-05 0 7.614e-05 3.3 7.606e-05 3.3 7.616e-05 0 7.607999999999999e-05 0 7.617999999999999e-05 3.3 7.609999999999999e-05 3.3 7.62e-05 0 7.612e-05 0 7.622e-05 3.3 7.614e-05 3.3 7.624e-05 0 7.616e-05 0 7.626e-05 3.3 7.617999999999999e-05 3.3 7.628e-05 0 7.62e-05 0 7.63e-05 3.3 7.622e-05 3.3 7.632e-05 0 7.624e-05 0 7.634e-05 3.3 7.625999999999999e-05 3.3 7.636e-05 0 7.628e-05 0 7.638e-05 3.3 7.63e-05 3.3 7.64e-05 0 7.632e-05 0 7.642e-05 3.3 7.633999999999999e-05 3.3 7.643999999999999e-05 0 7.636e-05 0 7.646e-05 3.3 7.638e-05 3.3 7.648e-05 0 7.64e-05 0 7.65e-05 3.3 7.641999999999999e-05 3.3 7.651999999999999e-05 0 7.643999999999999e-05 0 7.654e-05 3.3 7.646e-05 3.3 7.656e-05 0 7.648e-05 0 7.658e-05 3.3 7.65e-05 3.3 7.66e-05 0 7.651999999999999e-05 0 7.662e-05 3.3 7.654e-05 3.3 7.664e-05 0 7.656e-05 0 7.666e-05 3.3 7.658e-05 3.3 7.668e-05 0 7.659999999999999e-05 0 7.67e-05 3.3 7.662e-05 3.3 7.672e-05 0 7.664e-05 0 7.674e-05 3.3 7.666e-05 3.3 7.676e-05 0 7.667999999999999e-05 0 7.678e-05 3.3 7.67e-05 3.3 7.68e-05 0 7.672e-05 0 7.682e-05 3.3 7.674e-05 3.3 7.684e-05 0 7.675999999999999e-05 0 7.685999999999999e-05 3.3 7.678e-05 3.3 7.688e-05 0 7.68e-05 0 7.69e-05 3.3 7.682e-05 3.3 7.692e-05 0 7.683999999999999e-05 0 7.693999999999999e-05 3.3 7.685999999999999e-05 3.3 7.696e-05 0 7.688e-05 0 7.698e-05 3.3 7.69e-05 3.3 7.7e-05 0 7.692e-05 0 7.702e-05 3.3 7.693999999999999e-05 3.3 7.704e-05 0 7.696e-05 0 7.706e-05 3.3 7.698e-05 3.3 7.708e-05 0 7.7e-05 0 7.71e-05 3.3 7.701999999999999e-05 3.3 7.712e-05 0 7.704e-05 0 7.714e-05 3.3 7.706e-05 3.3 7.716e-05 0 7.708e-05 0 7.718e-05 3.3 7.709999999999999e-05 3.3 7.719999999999999e-05 0 7.712e-05 0 7.722e-05 3.3 7.714e-05 3.3 7.724e-05 0 7.716e-05 0 7.726e-05 3.3 7.717999999999999e-05 3.3 7.727999999999999e-05 0 7.719999999999999e-05 0 7.73e-05 3.3 7.722e-05 3.3 7.732e-05 0 7.724e-05 0 7.734e-05 3.3 7.726e-05 3.3 7.736e-05 0 7.727999999999999e-05 0 7.738e-05 3.3 7.73e-05 3.3 7.74e-05 0 7.732e-05 0 7.742e-05 3.3 7.734e-05 3.3 7.744e-05 0 7.735999999999999e-05 0 7.746e-05 3.3 7.738e-05 3.3 7.748e-05 0 7.74e-05 0 7.75e-05 3.3 7.742e-05 3.3 7.752e-05 0 7.743999999999999e-05 0 7.753999999999999e-05 3.3 7.746e-05 3.3 7.756e-05 0 7.748e-05 0 7.758e-05 3.3 7.75e-05 3.3 7.76e-05 0 7.751999999999999e-05 0 7.761999999999999e-05 3.3 7.753999999999999e-05 3.3 7.764e-05 0 7.756e-05 0 7.766e-05 3.3 7.758e-05 3.3 7.768e-05 0 7.76e-05 0 7.77e-05 3.3 7.761999999999999e-05 3.3 7.772e-05 0 7.764e-05 0 7.774e-05 3.3 7.766e-05 3.3 7.776e-05 0 7.768e-05 0 7.778e-05 3.3 7.769999999999999e-05 3.3 7.78e-05 0 7.772e-05 0 7.782e-05 3.3 7.774e-05 3.3 7.784e-05 0 7.776e-05 0 7.786e-05 3.3 7.777999999999999e-05 3.3 7.787999999999999e-05 0 7.78e-05 0 7.79e-05 3.3 7.782e-05 3.3 7.792e-05 0 7.784e-05 0 7.794e-05 3.3 7.785999999999999e-05 3.3 7.795999999999999e-05 0 7.787999999999999e-05 0 7.798e-05 3.3 7.79e-05 3.3 7.8e-05 0 7.792e-05 0 7.802e-05 3.3 7.794e-05 3.3 7.804e-05 0 7.795999999999999e-05 0 7.806e-05 3.3 7.798e-05 3.3 7.808e-05 0 7.8e-05 0 7.81e-05 3.3 7.802e-05 3.3 7.812e-05 0 7.803999999999999e-05 0 7.814e-05 3.3 7.806e-05 3.3 7.816e-05 0 7.808e-05 0 7.818e-05 3.3 7.81e-05 3.3 7.82e-05 0 7.811999999999999e-05 0 7.821999999999999e-05 3.3 7.814e-05 3.3 7.824e-05 0 7.816e-05 0 7.826e-05 3.3 7.818e-05 3.3 7.828e-05 0 7.819999999999999e-05 0 7.829999999999999e-05 3.3 7.821999999999999e-05 3.3 7.832e-05 0 7.824e-05 0 7.834e-05 3.3 7.826e-05 3.3 7.836e-05 0 7.828e-05 0 7.838e-05 3.3 7.829999999999999e-05 3.3 7.84e-05 0 7.832e-05 0 7.842e-05 3.3 7.834e-05 3.3 7.844e-05 0 7.836e-05 0 7.846e-05 3.3 7.837999999999999e-05 3.3 7.848e-05 0 7.84e-05 0 7.85e-05 3.3 7.842e-05 3.3 7.852e-05 0 7.844e-05 0 7.854e-05 3.3 7.845999999999999e-05 3.3 7.856e-05 0 7.848e-05 0 7.858e-05 3.3 7.85e-05 3.3 7.86e-05 0 7.852e-05 0 7.862e-05 3.3 7.853999999999999e-05 3.3 7.863999999999999e-05 0 7.856e-05 0 7.866e-05 3.3 7.858e-05 3.3 7.868e-05 0 7.86e-05 0 7.87e-05 3.3 7.861999999999999e-05 3.3 7.871999999999999e-05 0 7.863999999999999e-05 0 7.874e-05 3.3 7.866e-05 3.3 7.876e-05 0 7.868e-05 0 7.878e-05 3.3 7.87e-05 3.3 7.88e-05 0 7.871999999999999e-05 0 7.882e-05 3.3 7.874e-05 3.3 7.884e-05 0 7.876e-05 0 7.886e-05 3.3 7.878e-05 3.3 7.888e-05 0 7.879999999999999e-05 0 7.89e-05 3.3 7.882e-05 3.3 7.892e-05 0 7.884e-05 0 7.894e-05 3.3 7.886e-05 3.3 7.896e-05 0 7.887999999999999e-05 0 7.897999999999999e-05 3.3 7.89e-05 3.3 7.9e-05 0 7.892e-05 0 7.902e-05 3.3 7.894e-05 3.3 7.904e-05 0 7.895999999999999e-05 0 7.905999999999999e-05 3.3 7.897999999999999e-05 3.3 7.908e-05 0 7.9e-05 0 7.91e-05 3.3 7.902e-05 3.3 7.912e-05 0 7.904e-05 0 7.914e-05 3.3 7.905999999999999e-05 3.3 7.916e-05 0 7.908e-05 0 7.918e-05 3.3 7.91e-05 3.3 7.92e-05 0 7.912e-05 0 7.922e-05 3.3 7.913999999999999e-05 3.3 7.924e-05 0 7.916e-05 0 7.926e-05 3.3 7.918e-05 3.3 7.928e-05 0 7.92e-05 0 7.93e-05 3.3 7.921999999999999e-05 3.3 7.931999999999999e-05 0 7.924e-05 0 7.934e-05 3.3 7.926e-05 3.3 7.936e-05 0 7.928e-05 0 7.938e-05 3.3 7.929999999999999e-05 3.3 7.939999999999999e-05 0 7.931999999999999e-05 0 7.942e-05 3.3 7.934e-05 3.3 7.944e-05 0 7.936e-05 0 7.946e-05 3.3 7.938e-05 3.3 7.948e-05 0 7.939999999999999e-05 0 7.95e-05 3.3 7.942e-05 3.3 7.952e-05 0 7.944e-05 0 7.954e-05 3.3 7.946e-05 3.3 7.956e-05 0 7.947999999999999e-05 0 7.958e-05 3.3 7.95e-05 3.3 7.96e-05 0 7.952e-05 0 7.962e-05 3.3 7.954e-05 3.3 7.964e-05 0 7.955999999999999e-05 0 7.965999999999999e-05 3.3 7.958e-05 3.3 7.968e-05 0 7.96e-05 0 7.97e-05 3.3 7.962e-05 3.3 7.972e-05 0 7.963999999999999e-05 0 7.973999999999999e-05 3.3 7.965999999999999e-05 3.3 7.976e-05 0 7.968e-05 0 7.978e-05 3.3 7.97e-05 3.3 7.98e-05 0 7.972e-05 0 7.982e-05 3.3 7.973999999999999e-05 3.3 7.984e-05 0 7.976e-05 0 7.986e-05 3.3 7.978e-05 3.3 7.988e-05 0 7.98e-05 0 7.99e-05 3.3 7.981999999999999e-05 3.3 7.992e-05 0 7.984e-05 0 7.994e-05 3.3 7.986e-05 3.3 7.996e-05 0 7.988e-05 0 7.998e-05 3.3 7.989999999999999e-05 3.3 7.999999999999999e-05 0 7.992e-05 0 8.002e-05 3.3 7.994e-05 3.3 8.004e-05 0 7.996e-05 0 8.006e-05 3.3 7.997999999999999e-05 3.3 8.007999999999999e-05 0 7.999999999999999e-05 0 8.01e-05 3.3 8.002e-05 3.3 8.012e-05 0 8.004e-05 0 8.014e-05 3.3 8.006e-05 3.3 8.016e-05 0 8.007999999999999e-05 0 8.018e-05 3.3 8.01e-05 3.3 8.02e-05 0 8.012e-05 0 8.022e-05 3.3 8.014e-05 3.3 8.024e-05 0 8.015999999999999e-05 0 8.026e-05 3.3 8.018e-05 3.3 8.028e-05 0 8.02e-05 0 8.03e-05 3.3 8.022e-05 3.3 8.032e-05 0 8.023999999999999e-05 0 8.033999999999999e-05 3.3 8.026e-05 3.3 8.036e-05 0 8.028e-05 0 8.038e-05 3.3 8.03e-05 3.3 8.04e-05 0 8.031999999999999e-05 0 8.041999999999999e-05 3.3 8.033999999999999e-05 3.3 8.044e-05 0 8.036e-05 0 8.046e-05 3.3 8.038e-05 3.3 8.048e-05 0 8.04e-05 0 8.05e-05 3.3 8.041999999999999e-05 3.3 8.052e-05 0 8.044e-05 0 8.054e-05 3.3 8.046e-05 3.3 8.056e-05 0 8.048e-05 0 8.058e-05 3.3 8.049999999999999e-05 3.3 8.06e-05 0 8.052e-05 0 8.062e-05 3.3 8.054e-05 3.3 8.064e-05 0 8.056e-05 0 8.066e-05 3.3 8.057999999999999e-05 3.3 8.068e-05 0 8.06e-05 0 8.07e-05 3.3 8.062e-05 3.3 8.072e-05 0 8.064e-05 0 8.074e-05 3.3 8.065999999999999e-05 3.3 8.075999999999999e-05 0 8.068e-05 0 8.078e-05 3.3 8.07e-05 3.3 8.08e-05 0 8.072e-05 0 8.082e-05 3.3 8.073999999999999e-05 3.3 8.083999999999999e-05 0 8.075999999999999e-05 0 8.086e-05 3.3 8.078e-05 3.3 8.088e-05 0 8.08e-05 0 8.09e-05 3.3 8.082e-05 3.3 8.092e-05 0 8.083999999999999e-05 0 8.094e-05 3.3 8.086e-05 3.3 8.096e-05 0 8.088e-05 0 8.098e-05 3.3 8.09e-05 3.3 8.1e-05 0 8.091999999999999e-05 0 8.102e-05 3.3 8.094e-05 3.3 8.104e-05 0 8.096e-05 0 8.106e-05 3.3 8.098e-05 3.3 8.108e-05 0 8.099999999999999e-05 0 8.109999999999999e-05 3.3 8.102e-05 3.3 8.112e-05 0 8.104e-05 0 8.114e-05 3.3 8.106e-05 3.3 8.116e-05 0 8.107999999999999e-05 0 8.117999999999999e-05 3.3 8.109999999999999e-05 3.3 8.12e-05 0 8.112e-05 0 8.122e-05 3.3 8.114e-05 3.3 8.124e-05 0 8.116e-05 0 8.126e-05 3.3 8.117999999999999e-05 3.3 8.128e-05 0 8.12e-05 0 8.13e-05 3.3 8.122e-05 3.3 8.132e-05 0 8.124e-05 0 8.134e-05 3.3 8.125999999999999e-05 3.3 8.136e-05 0 8.128e-05 0 8.138e-05 3.3 8.13e-05 3.3 8.14e-05 0 8.132e-05 0 8.142e-05 3.3 8.133999999999999e-05 3.3 8.143999999999999e-05 0 8.136e-05 0 8.146e-05 3.3 8.138e-05 3.3 8.148e-05 0 8.14e-05 0 8.15e-05 3.3 8.141999999999999e-05 3.3 8.151999999999999e-05 0 8.143999999999999e-05 0 8.154e-05 3.3 8.146e-05 3.3 8.156e-05 0 8.148e-05 0 8.158e-05 3.3 8.15e-05 3.3 8.16e-05 0 8.151999999999999e-05 0 8.162e-05 3.3 8.154e-05 3.3 8.164e-05 0 8.156e-05 0 8.166e-05 3.3 8.158e-05 3.3 8.168e-05 0 8.159999999999999e-05 0 8.17e-05 3.3 8.162e-05 3.3 8.172e-05 0 8.164e-05 0 8.174e-05 3.3 8.166e-05 3.3 8.176e-05 0 8.167999999999999e-05 0 8.177999999999999e-05 3.3 8.17e-05 3.3 8.18e-05 0 8.172e-05 0 8.182e-05 3.3 8.174e-05 3.3 8.184e-05 0 8.175999999999999e-05 0 8.185999999999999e-05 3.3 8.177999999999999e-05 3.3 8.188e-05 0 8.18e-05 0 8.19e-05 3.3 8.182e-05 3.3 8.192e-05 0 8.184e-05 0 8.194e-05 3.3 8.185999999999999e-05 3.3 8.196e-05 0 8.188e-05 0 8.198e-05 3.3 8.19e-05 3.3 8.2e-05 0 8.192e-05 0 8.202e-05 3.3 8.193999999999999e-05 3.3 8.204e-05 0 8.196e-05 0 8.206e-05 3.3 8.198e-05 3.3 8.208e-05 0 8.2e-05 0 8.21e-05 3.3 8.201999999999999e-05 3.3 8.211999999999999e-05 0 8.204e-05 0 8.214e-05 3.3 8.206e-05 3.3 8.216e-05 0 8.208e-05 0 8.218e-05 3.3 8.209999999999999e-05 3.3 8.219999999999999e-05 0 8.211999999999999e-05 0 8.222e-05 3.3 8.214e-05 3.3 8.224e-05 0 8.216e-05 0 8.226e-05 3.3 8.218e-05 3.3 8.228e-05 0 8.219999999999999e-05 0 8.23e-05 3.3 8.222e-05 3.3 8.232e-05 0 8.224e-05 0 8.234e-05 3.3 8.226e-05 3.3 8.236e-05 0 8.227999999999999e-05 0 8.238e-05 3.3 8.23e-05 3.3 8.24e-05 0 8.232e-05 0 8.242e-05 3.3 8.234e-05 3.3 8.244e-05 0 8.235999999999999e-05 0 8.245999999999999e-05 3.3 8.238e-05 3.3 8.248e-05 0 8.24e-05 0 8.25e-05 3.3 8.242e-05 3.3 8.252e-05 0 8.243999999999999e-05 0 8.253999999999999e-05 3.3 8.245999999999999e-05 3.3 8.256e-05 0 8.248e-05 0 8.258e-05 3.3 8.25e-05 3.3 8.26e-05 0 8.251999999999999e-05 0 8.261999999999999e-05 3.3 8.253999999999999e-05 3.3 8.264e-05 0 8.256e-05 0 8.266e-05 3.3 8.258e-05 3.3 8.268e-05 0 8.26e-05 0 8.27e-05 3.3 8.261999999999999e-05 3.3 8.272e-05 0 8.264e-05 0 8.274e-05 3.3 8.266e-05 3.3 8.276e-05 0 8.268e-05 0 8.278e-05 3.3 8.269999999999999e-05 3.3 8.28e-05 0 8.272e-05 0 8.282e-05 3.3 8.274e-05 3.3 8.284e-05 0 8.276e-05 0 8.286e-05 3.3 8.277999999999999e-05 3.3 8.287999999999999e-05 0 8.28e-05 0 8.29e-05 3.3 8.282e-05 3.3 8.292e-05 0 8.284e-05 0 8.294e-05 3.3 8.285999999999999e-05 3.3 8.295999999999999e-05 0 8.287999999999999e-05 0 8.298e-05 3.3 8.29e-05 3.3 8.3e-05 0 8.292e-05 0 8.302e-05 3.3 8.294e-05 3.3 8.304e-05 0 8.295999999999999e-05 0 8.306e-05 3.3 8.298e-05 3.3 8.308e-05 0 8.3e-05 0 8.31e-05 3.3 8.302e-05 3.3 8.312e-05 0 8.303999999999999e-05 0 8.314e-05 3.3 8.306e-05 3.3 8.316e-05 0 8.308e-05 0 8.318e-05 3.3 8.31e-05 3.3 8.32e-05 0 8.311999999999999e-05 0 8.321999999999999e-05 3.3 8.314e-05 3.3 8.324e-05 0 8.316e-05 0 8.326e-05 3.3 8.318e-05 3.3 8.328e-05 0 8.319999999999999e-05 0 8.329999999999999e-05 3.3 8.321999999999999e-05 3.3 8.332e-05 0 8.324e-05 0 8.334e-05 3.3 8.326e-05 3.3 8.336e-05 0 8.328e-05 0 8.338e-05 3.3 8.329999999999999e-05 3.3 8.34e-05 0 8.332e-05 0 8.342e-05 3.3 8.334e-05 3.3 8.344e-05 0 8.336e-05 0 8.346e-05 3.3 8.337999999999999e-05 3.3 8.348e-05 0 8.34e-05 0 8.35e-05 3.3 8.342e-05 3.3 8.352e-05 0 8.344e-05 0 8.354e-05 3.3 8.345999999999999e-05 3.3 8.355999999999999e-05 0 8.348e-05 0 8.358e-05 3.3 8.35e-05 3.3 8.36e-05 0 8.352e-05 0 8.362e-05 3.3 8.353999999999999e-05 3.3 8.363999999999999e-05 0 8.355999999999999e-05 0 8.366e-05 3.3 8.358e-05 3.3 8.368e-05 0 8.36e-05 0 8.37e-05 3.3 8.362e-05 3.3 8.372e-05 0 8.363999999999999e-05 0 8.374e-05 3.3 8.366e-05 3.3 8.376e-05 0 8.368e-05 0 8.378e-05 3.3 8.37e-05 3.3 8.38e-05 0 8.371999999999999e-05 0 8.382e-05 3.3 8.374e-05 3.3 8.384e-05 0 8.376e-05 0 8.386e-05 3.3 8.378e-05 3.3 8.388e-05 0 8.379999999999999e-05 0 8.389999999999999e-05 3.3 8.382e-05 3.3 8.392e-05 0 8.384e-05 0 8.394e-05 3.3 8.386e-05 3.3 8.396e-05 0 8.387999999999999e-05 0 8.397999999999999e-05 3.3 8.389999999999999e-05 3.3 8.4e-05 0 8.392e-05 0 8.402e-05 3.3 8.394e-05 3.3 8.404e-05 0 8.396e-05 0 8.406e-05 3.3 8.397999999999999e-05 3.3 8.408e-05 0 8.4e-05 0 8.41e-05 3.3 8.402e-05 3.3 8.412e-05 0 8.404e-05 0 8.414e-05 3.3 8.405999999999999e-05 3.3 8.416e-05 0 8.408e-05 0 8.418e-05 3.3 8.41e-05 3.3 8.42e-05 0 8.412e-05 0 8.422e-05 3.3 8.413999999999999e-05 3.3 8.423999999999999e-05 0 8.416e-05 0 8.426e-05 3.3 8.418e-05 3.3 8.428e-05 0 8.42e-05 0 8.43e-05 3.3 8.421999999999999e-05 3.3 8.431999999999999e-05 0 8.423999999999999e-05 0 8.434e-05 3.3 8.426e-05 3.3 8.436e-05 0 8.428e-05 0 8.438e-05 3.3 8.43e-05 3.3 8.44e-05 0 8.431999999999999e-05 0 8.442e-05 3.3 8.434e-05 3.3 8.444e-05 0 8.436e-05 0 8.446e-05 3.3 8.438e-05 3.3 8.448e-05 0 8.439999999999999e-05 0 8.45e-05 3.3 8.442e-05 3.3 8.452e-05 0 8.444e-05 0 8.454e-05 3.3 8.446e-05 3.3 8.456e-05 0 8.447999999999999e-05 0 8.457999999999999e-05 3.3 8.45e-05 3.3 8.46e-05 0 8.452e-05 0 8.462e-05 3.3 8.454e-05 3.3 8.464e-05 0 8.455999999999999e-05 0 8.465999999999999e-05 3.3 8.457999999999999e-05 3.3 8.468e-05 0 8.46e-05 0 8.47e-05 3.3 8.462e-05 3.3 8.472e-05 0 8.463999999999999e-05 0 8.473999999999999e-05 3.3 8.465999999999999e-05 3.3 8.476e-05 0 8.468e-05 0 8.478e-05 3.3 8.47e-05 3.3 8.48e-05 0 8.472e-05 0 8.482e-05 3.3 8.473999999999999e-05 3.3 8.484e-05 0 8.476e-05 0 8.486e-05 3.3 8.478e-05 3.3 8.488e-05 0 8.48e-05 0 8.49e-05 3.3 8.481999999999999e-05 3.3 8.492e-05 0 8.484e-05 0 8.494e-05 3.3 8.486e-05 3.3 8.496e-05 0 8.488e-05 0 8.498e-05 3.3 8.489999999999999e-05 3.3 8.499999999999999e-05 0 8.492e-05 0 8.502e-05 3.3 8.494e-05 3.3 8.504e-05 0 8.496e-05 0 8.506e-05 3.3 8.497999999999999e-05 3.3 8.507999999999999e-05 0 8.499999999999999e-05 0 8.51e-05 3.3 8.502e-05 3.3 8.512e-05 0 8.504e-05 0 8.514e-05 3.3 8.506e-05 3.3 8.516e-05 0 8.507999999999999e-05 0 8.518e-05 3.3 8.51e-05 3.3 8.52e-05 0 8.512e-05 0 8.522e-05 3.3 8.514e-05 3.3 8.524e-05 0 8.515999999999999e-05 0 8.526e-05 3.3 8.518e-05 3.3 8.528e-05 0 8.52e-05 0 8.53e-05 3.3 8.522e-05 3.3 8.532e-05 0 8.523999999999999e-05 0 8.533999999999999e-05 3.3 8.526e-05 3.3 8.536e-05 0 8.528e-05 0 8.538e-05 3.3 8.53e-05 3.3 8.54e-05 0 8.531999999999999e-05 0 8.541999999999999e-05 3.3 8.533999999999999e-05 3.3 8.544e-05 0 8.536e-05 0 8.546e-05 3.3 8.538e-05 3.3 8.548e-05 0 8.54e-05 0 8.55e-05 3.3 8.541999999999999e-05 3.3 8.552e-05 0 8.544e-05 0 8.554e-05 3.3 8.546e-05 3.3 8.556e-05 0 8.548e-05 0 8.558e-05 3.3 8.549999999999999e-05 3.3 8.56e-05 0 8.552e-05 0 8.562e-05 3.3 8.554e-05 3.3 8.564e-05 0 8.556e-05 0 8.566e-05 3.3 8.557999999999999e-05 3.3 8.567999999999999e-05 0 8.56e-05 0 8.57e-05 3.3 8.562e-05 3.3 8.572e-05 0 8.564e-05 0 8.574e-05 3.3 8.565999999999999e-05 3.3 8.575999999999999e-05 0 8.567999999999999e-05 0 8.578e-05 3.3 8.57e-05 3.3 8.58e-05 0 8.572e-05 0 8.582e-05 3.3 8.574e-05 3.3 8.584e-05 0 8.575999999999999e-05 0 8.586e-05 3.3 8.578e-05 3.3 8.588e-05 0 8.58e-05 0 8.59e-05 3.3 8.582e-05 3.3 8.592e-05 0 8.583999999999999e-05 0 8.594e-05 3.3 8.586e-05 3.3 8.596e-05 0 8.588e-05 0 8.598e-05 3.3 8.59e-05 3.3 8.6e-05 0 8.591999999999999e-05 0 8.601999999999999e-05 3.3 8.594e-05 3.3 8.604e-05 0 8.596e-05 0 8.606e-05 3.3 8.598e-05 3.3 8.608e-05 0 8.599999999999999e-05 0 8.609999999999999e-05 3.3 8.601999999999999e-05 3.3 8.612e-05 0 8.604e-05 0 8.614e-05 3.3 8.606e-05 3.3 8.616e-05 0 8.608e-05 0 8.618e-05 3.3 8.609999999999999e-05 3.3 8.62e-05 0 8.612e-05 0 8.622e-05 3.3 8.614e-05 3.3 8.624e-05 0 8.616e-05 0 8.626e-05 3.3 8.617999999999999e-05 3.3 8.628e-05 0 8.62e-05 0 8.63e-05 3.3 8.622e-05 3.3 8.632e-05 0 8.624e-05 0 8.634e-05 3.3 8.625999999999999e-05 3.3 8.635999999999999e-05 0 8.628e-05 0 8.638e-05 3.3 8.63e-05 3.3 8.64e-05 0 8.632e-05 0 8.642e-05 3.3 8.633999999999999e-05 3.3 8.643999999999999e-05 0 8.635999999999999e-05 0 8.646e-05 3.3 8.638e-05 3.3 8.648e-05 0 8.64e-05 0 8.65e-05 3.3 8.641999999999999e-05 3.3 8.651999999999999e-05 0 8.643999999999999e-05 0 8.654e-05 3.3 8.646e-05 3.3 8.656e-05 0 8.648e-05 0 8.658e-05 3.3 8.65e-05 3.3 8.66e-05 0 8.651999999999999e-05 0 8.662e-05 3.3 8.654e-05 3.3 8.664e-05 0 8.656e-05 0 8.666e-05 3.3 8.658e-05 3.3 8.668e-05 0 8.659999999999999e-05 0 8.669999999999999e-05 3.3 8.662e-05 3.3 8.672e-05 0 8.664e-05 0 8.674e-05 3.3 8.666e-05 3.3 8.676e-05 0 8.667999999999999e-05 0 8.677999999999999e-05 3.3 8.669999999999999e-05 3.3 8.68e-05 0 8.672e-05 0 8.682e-05 3.3 8.674e-05 3.3 8.684e-05 0 8.675999999999999e-05 0 8.685999999999999e-05 3.3 8.677999999999999e-05 3.3 8.688e-05 0 8.68e-05 0 8.69e-05 3.3 8.682e-05 3.3 8.692e-05 0 8.684e-05 0 8.694e-05 3.3 8.685999999999999e-05 3.3 8.696e-05 0 8.688e-05 0 8.698e-05 3.3 8.69e-05 3.3 8.7e-05 0 8.692e-05 0 8.702e-05 3.3 8.693999999999999e-05 3.3 8.704e-05 0 8.696e-05 0 8.706e-05 3.3 8.698e-05 3.3 8.708e-05 0 8.7e-05 0 8.71e-05 3.3 8.701999999999999e-05 3.3 8.711999999999999e-05 0 8.704e-05 0 8.714e-05 3.3 8.706e-05 3.3 8.716e-05 0 8.708e-05 0 8.718e-05 3.3 8.709999999999999e-05 3.3 8.719999999999999e-05 0 8.711999999999999e-05 0 8.722e-05 3.3 8.714e-05 3.3 8.724e-05 0 8.716e-05 0 8.726e-05 3.3 8.718e-05 3.3 8.728e-05 0 8.719999999999999e-05 0 8.73e-05 3.3 8.722e-05 3.3 8.732e-05 0 8.724e-05 0 8.734e-05 3.3 8.726e-05 3.3 8.736e-05 0 8.727999999999999e-05 0 8.738e-05 3.3 8.73e-05 3.3 8.74e-05 0 8.732e-05 0 8.742e-05 3.3 8.734e-05 3.3 8.744e-05 0 8.735999999999999e-05 0 8.745999999999999e-05 3.3 8.738e-05 3.3 8.748e-05 0 8.74e-05 0 8.75e-05 3.3 8.742e-05 3.3 8.752e-05 0 8.743999999999999e-05 0 8.753999999999999e-05 3.3 8.745999999999999e-05 3.3 8.756e-05 0 8.748e-05 0 8.758e-05 3.3 8.75e-05 3.3 8.76e-05 0 8.752e-05 0 8.762e-05 3.3 8.753999999999999e-05 3.3 8.764e-05 0 8.756e-05 0 8.766e-05 3.3 8.758e-05 3.3 8.768e-05 0 8.76e-05 0 8.77e-05 3.3 8.761999999999999e-05 3.3 8.772e-05 0 8.764e-05 0 8.774e-05 3.3 8.766e-05 3.3 8.776e-05 0 8.768e-05 0 8.778e-05 3.3 8.769999999999999e-05 3.3 8.779999999999999e-05 0 8.772e-05 0 8.782e-05 3.3 8.774e-05 3.3 8.784e-05 0 8.776e-05 0 8.786e-05 3.3 8.777999999999999e-05 3.3 8.787999999999999e-05 0 8.779999999999999e-05 0 8.79e-05 3.3 8.782e-05 3.3 8.792e-05 0 8.784e-05 0 8.794e-05 3.3 8.786e-05 3.3 8.796e-05 0 8.787999999999999e-05 0 8.798e-05 3.3 8.79e-05 3.3 8.8e-05 0 8.792e-05 0 8.802e-05 3.3 8.794e-05 3.3 8.804e-05 0 8.795999999999999e-05 0 8.806e-05 3.3 8.798e-05 3.3 8.808e-05 0 8.8e-05 0 8.81e-05 3.3 8.802e-05 3.3 8.812e-05 0 8.803999999999999e-05 0 8.813999999999999e-05 3.3 8.806e-05 3.3 8.816e-05 0 8.808e-05 0 8.818e-05 3.3 8.81e-05 3.3 8.82e-05 0 8.811999999999999e-05 0 8.821999999999999e-05 3.3 8.813999999999999e-05 3.3 8.824e-05 0 8.816e-05 0 8.826e-05 3.3 8.818e-05 3.3 8.828e-05 0 8.819999999999999e-05 0 8.829999999999999e-05 3.3 8.821999999999999e-05 3.3 8.832e-05 0 8.824e-05 0 8.834e-05 3.3 8.826e-05 3.3 8.836e-05 0 8.828e-05 0 8.838e-05 3.3 8.829999999999999e-05 3.3 8.84e-05 0 8.832e-05 0 8.842e-05 3.3 8.834e-05 3.3 8.844e-05 0 8.836e-05 0 8.846e-05 3.3 8.837999999999999e-05 3.3 8.847999999999999e-05 0 8.84e-05 0 8.85e-05 3.3 8.842e-05 3.3 8.852e-05 0 8.844e-05 0 8.854e-05 3.3 8.845999999999999e-05 3.3 8.855999999999999e-05 0 8.847999999999999e-05 0 8.858e-05 3.3 8.85e-05 3.3 8.86e-05 0 8.852e-05 0 8.862e-05 3.3 8.853999999999999e-05 3.3 8.863999999999999e-05 0 8.855999999999999e-05 0 8.866e-05 3.3 8.858e-05 3.3 8.868e-05 0 8.86e-05 0 8.87e-05 3.3 8.862e-05 3.3 8.872e-05 0 8.863999999999999e-05 0 8.874e-05 3.3 8.866e-05 3.3 8.876e-05 0 8.868e-05 0 8.878e-05 3.3 8.87e-05 3.3 8.88e-05 0 8.871999999999999e-05 0 8.882e-05 3.3 8.874e-05 3.3 8.884e-05 0 8.876e-05 0 8.886e-05 3.3 8.878e-05 3.3 8.888e-05 0 8.879999999999999e-05 0 8.889999999999999e-05 3.3 8.882e-05 3.3 8.892e-05 0 8.884e-05 0 8.894e-05 3.3 8.886e-05 3.3 8.896e-05 0 8.887999999999999e-05 0 8.897999999999999e-05 3.3 8.889999999999999e-05 3.3 8.9e-05 0 8.892e-05 0 8.902e-05 3.3 8.894e-05 3.3 8.904e-05 0 8.896e-05 0 8.906e-05 3.3 8.897999999999999e-05 3.3 8.908e-05 0 8.9e-05 0 8.91e-05 3.3 8.902e-05 3.3 8.912e-05 0 8.904e-05 0 8.914e-05 3.3 8.905999999999999e-05 3.3 8.916e-05 0 8.908e-05 0 8.918e-05 3.3 8.91e-05 3.3 8.92e-05 0 8.912e-05 0 8.922e-05 3.3 8.913999999999999e-05 3.3 8.923999999999999e-05 0 8.916e-05 0 8.926e-05 3.3 8.918e-05 3.3 8.928e-05 0 8.92e-05 0 8.93e-05 3.3 8.921999999999999e-05 3.3 8.931999999999999e-05 0 8.923999999999999e-05 0 8.934e-05 3.3 8.926e-05 3.3 8.936e-05 0 8.928e-05 0 8.938e-05 3.3 8.93e-05 3.3 8.94e-05 0 8.931999999999999e-05 0 8.942e-05 3.3 8.934e-05 3.3 8.944e-05 0 8.936e-05 0 8.946e-05 3.3 8.938e-05 3.3 8.948e-05 0 8.939999999999999e-05 0 8.95e-05 3.3 8.942e-05 3.3 8.952e-05 0 8.944e-05 0 8.954e-05 3.3 8.946e-05 3.3 8.956e-05 0 8.947999999999999e-05 0 8.957999999999999e-05 3.3 8.95e-05 3.3 8.96e-05 0 8.952e-05 0 8.962e-05 3.3 8.954e-05 3.3 8.964e-05 0 8.955999999999999e-05 0 8.965999999999999e-05 3.3 8.957999999999999e-05 3.3 8.968e-05 0 8.96e-05 0 8.97e-05 3.3 8.962e-05 3.3 8.972e-05 0 8.964e-05 0 8.974e-05 3.3 8.965999999999999e-05 3.3 8.976e-05 0 8.968e-05 0 8.978e-05 3.3 8.97e-05 3.3 8.98e-05 0 8.972e-05 0 8.982e-05 3.3 8.973999999999999e-05 3.3 8.984e-05 0 8.976e-05 0 8.986e-05 3.3 8.978e-05 3.3 8.988e-05 0 8.98e-05 0 8.99e-05 3.3 8.981999999999999e-05 3.3 8.991999999999999e-05 0 8.984e-05 0 8.994e-05 3.3 8.986e-05 3.3 8.996e-05 0 8.988e-05 0 8.998e-05 3.3 8.989999999999999e-05 3.3 8.999999999999999e-05 0 8.991999999999999e-05 0 9.002e-05 3.3 8.994e-05 3.3 9.004e-05 0 8.996e-05 0 9.006e-05 3.3 8.998e-05 3.3 9.008e-05 0 8.999999999999999e-05 0 9.01e-05 3.3 9.002e-05 3.3 9.012e-05 0 9.004e-05 0 9.014e-05 3.3 9.006e-05 3.3 9.016e-05 0 9.007999999999999e-05 0 9.018e-05 3.3 9.01e-05 3.3 9.02e-05 0 9.012e-05 0 9.022e-05 3.3 9.014e-05 3.3 9.024e-05 0 9.015999999999999e-05 0 9.025999999999999e-05 3.3 9.018e-05 3.3 9.028e-05 0 9.02e-05 0 9.03e-05 3.3 9.022e-05 3.3 9.032e-05 0 9.023999999999999e-05 0 9.033999999999999e-05 3.3 9.025999999999999e-05 3.3 9.036e-05 0 9.028e-05 0 9.038e-05 3.3 9.03e-05 3.3 9.04e-05 0 9.031999999999999e-05 0 9.041999999999999e-05 3.3 9.033999999999999e-05 3.3 9.044e-05 0 9.036e-05 0 9.046e-05 3.3 9.038e-05 3.3 9.048e-05 0 9.04e-05 0 9.05e-05 3.3 9.041999999999999e-05 3.3 9.052e-05 0 9.044e-05 0 9.054e-05 3.3 9.046e-05 3.3 9.056e-05 0 9.048e-05 0 9.058e-05 3.3 9.049999999999999e-05 3.3 9.059999999999999e-05 0 9.052e-05 0 9.062e-05 3.3 9.054e-05 3.3 9.064e-05 0 9.056e-05 0 9.066e-05 3.3 9.057999999999999e-05 3.3 9.067999999999999e-05 0 9.059999999999999e-05 0 9.07e-05 3.3 9.062e-05 3.3 9.072e-05 0 9.064e-05 0 9.074e-05 3.3 9.065999999999999e-05 3.3 9.075999999999999e-05 0 9.067999999999999e-05 0 9.078e-05 3.3 9.07e-05 3.3 9.08e-05 0 9.072e-05 0 9.082e-05 3.3 9.074e-05 3.3 9.084e-05 0 9.075999999999999e-05 0 9.086e-05 3.3 9.078e-05 3.3 9.088e-05 0 9.08e-05 0 9.09e-05 3.3 9.082e-05 3.3 9.092e-05 0 9.083999999999999e-05 0 9.094e-05 3.3 9.086e-05 3.3 9.096e-05 0 9.088e-05 0 9.098e-05 3.3 9.09e-05 3.3 9.1e-05 0 9.091999999999999e-05 0 9.101999999999999e-05 3.3 9.094e-05 3.3 9.104e-05 0 9.096e-05 0 9.106e-05 3.3 9.098e-05 3.3 9.108e-05 0 9.099999999999999e-05 0 9.109999999999999e-05 3.3 9.101999999999999e-05 3.3 9.112e-05 0 9.104e-05 0 9.114e-05 3.3 9.106e-05 3.3 9.116e-05 0 9.108e-05 0 9.118e-05 3.3 9.109999999999999e-05 3.3 9.12e-05 0 9.112e-05 0 9.122e-05 3.3 9.114e-05 3.3 9.124e-05 0 9.116e-05 0 9.126e-05 3.3 9.117999999999999e-05 3.3 9.128e-05 0 9.12e-05 0 9.13e-05 3.3 9.122e-05 3.3 9.132e-05 0 9.124e-05 0 9.134e-05 3.3 9.125999999999999e-05 3.3 9.135999999999999e-05 0 9.128e-05 0 9.138e-05 3.3 9.13e-05 3.3 9.14e-05 0 9.132e-05 0 9.142e-05 3.3 9.133999999999999e-05 3.3 9.143999999999999e-05 0 9.135999999999999e-05 0 9.146e-05 3.3 9.138e-05 3.3 9.148e-05 0 9.14e-05 0 9.15e-05 3.3 9.142e-05 3.3 9.152e-05 0 9.143999999999999e-05 0 9.154e-05 3.3 9.146e-05 3.3 9.156e-05 0 9.148e-05 0 9.158e-05 3.3 9.15e-05 3.3 9.16e-05 0 9.151999999999999e-05 0 9.162e-05 3.3 9.154e-05 3.3 9.164e-05 0 9.156e-05 0 9.166e-05 3.3 9.158e-05 3.3 9.168e-05 0 9.159999999999999e-05 0 9.169999999999999e-05 3.3 9.162e-05 3.3 9.172e-05 0 9.164e-05 0 9.174e-05 3.3 9.166e-05 3.3 9.176e-05 0 9.167999999999999e-05 0 9.177999999999999e-05 3.3 9.169999999999999e-05 3.3 9.18e-05 0 9.172e-05 0 9.182e-05 3.3 9.174e-05 3.3 9.184e-05 0 9.176e-05 0 9.186e-05 3.3 9.177999999999999e-05 3.3 9.188e-05 0 9.18e-05 0 9.19e-05 3.3 9.182e-05 3.3 9.192e-05 0 9.184e-05 0 9.194e-05 3.3 9.185999999999999e-05 3.3 9.196e-05 0 9.188e-05 0 9.198e-05 3.3 9.19e-05 3.3 9.2e-05 0 9.192e-05 0 9.202e-05 3.3 9.193999999999999e-05 3.3 9.203999999999999e-05 0 9.196e-05 0 9.206e-05 3.3 9.198e-05 3.3 9.208e-05 0 9.2e-05 0 9.21e-05 3.3 9.201999999999999e-05 3.3 9.211999999999999e-05 0 9.203999999999999e-05 0 9.214e-05 3.3 9.206e-05 3.3 9.216e-05 0 9.208e-05 0 9.218e-05 3.3 9.209999999999999e-05 3.3 9.219999999999999e-05 0 9.211999999999999e-05 0 9.222e-05 3.3 9.214e-05 3.3 9.224e-05 0 9.216e-05 0 9.226e-05 3.3 9.218e-05 3.3 9.228e-05 0 9.219999999999999e-05 0 9.23e-05 3.3 9.222e-05 3.3 9.232e-05 0 9.224e-05 0 9.234e-05 3.3 9.226e-05 3.3 9.236e-05 0 9.227999999999999e-05 0 9.237999999999999e-05 3.3 9.23e-05 3.3 9.24e-05 0 9.232e-05 0 9.242e-05 3.3 9.234e-05 3.3 9.244e-05 0 9.235999999999999e-05 0 9.245999999999999e-05 3.3 9.237999999999999e-05 3.3 9.248e-05 0 9.24e-05 0 9.25e-05 3.3 9.242e-05 3.3 9.252e-05 0 9.243999999999999e-05 0 9.253999999999999e-05 3.3 9.245999999999999e-05 3.3 9.256e-05 0 9.248e-05 0 9.258e-05 3.3 9.25e-05 3.3 9.26e-05 0 9.252e-05 0 9.262e-05 3.3 9.253999999999999e-05 3.3 9.264e-05 0 9.256e-05 0 9.266e-05 3.3 9.258e-05 3.3 9.268e-05 0 9.26e-05 0 9.27e-05 3.3 9.261999999999999e-05 3.3 9.271999999999999e-05 0 9.264e-05 0 9.274e-05 3.3 9.266e-05 3.3 9.276e-05 0 9.268e-05 0 9.278e-05 3.3 9.269999999999999e-05 3.3 9.279999999999999e-05 0 9.271999999999999e-05 0 9.282e-05 3.3 9.274e-05 3.3 9.284e-05 0 9.276e-05 0 9.286e-05 3.3 9.277999999999999e-05 3.3 9.287999999999999e-05 0 9.279999999999999e-05 0 9.29e-05 3.3 9.282e-05 3.3 9.292e-05 0 9.284e-05 0 9.294e-05 3.3 9.286e-05 3.3 9.296e-05 0 9.287999999999999e-05 0 9.298e-05 3.3 9.29e-05 3.3 9.3e-05 0 9.292e-05 0 9.302e-05 3.3 9.294e-05 3.3 9.304e-05 0 9.295999999999999e-05 0 9.306e-05 3.3 9.298e-05 3.3 9.308e-05 0 9.3e-05 0 9.31e-05 3.3 9.302e-05 3.3 9.312e-05 0 9.303999999999999e-05 0 9.313999999999999e-05 3.3 9.306e-05 3.3 9.316e-05 0 9.308e-05 0 9.318e-05 3.3 9.31e-05 3.3 9.32e-05 0 9.311999999999999e-05 0 9.321999999999999e-05 3.3 9.313999999999999e-05 3.3 9.324e-05 0 9.316e-05 0 9.326e-05 3.3 9.318e-05 3.3 9.328e-05 0 9.32e-05 0 9.33e-05 3.3 9.321999999999999e-05 3.3 9.332e-05 0 9.324e-05 0 9.334e-05 3.3 9.326e-05 3.3 9.336e-05 0 9.328e-05 0 9.338e-05 3.3 9.329999999999999e-05 3.3 9.34e-05 0 9.332e-05 0 9.342e-05 3.3 9.334e-05 3.3 9.344e-05 0 9.336e-05 0 9.346e-05 3.3 9.337999999999999e-05 3.3 9.347999999999999e-05 0 9.34e-05 0 9.35e-05 3.3 9.342e-05 3.3 9.352e-05 0 9.344e-05 0 9.354e-05 3.3 9.345999999999999e-05 3.3 9.355999999999999e-05 0 9.347999999999999e-05 0 9.358e-05 3.3 9.35e-05 3.3 9.36e-05 0 9.352e-05 0 9.362e-05 3.3 9.354e-05 3.3 9.364e-05 0 9.355999999999999e-05 0 9.366e-05 3.3 9.358e-05 3.3 9.368e-05 0 9.36e-05 0 9.37e-05 3.3 9.362e-05 3.3 9.372e-05 0 9.363999999999999e-05 0 9.374e-05 3.3 9.366e-05 3.3 9.376e-05 0 9.368e-05 0 9.378e-05 3.3 9.37e-05 3.3 9.38e-05 0 9.371999999999999e-05 0 9.381999999999999e-05 3.3 9.374e-05 3.3 9.384e-05 0 9.376e-05 0 9.386e-05 3.3 9.378e-05 3.3 9.388e-05 0 9.379999999999999e-05 0 9.389999999999999e-05 3.3 9.381999999999999e-05 3.3 9.392e-05 0 9.384e-05 0 9.394e-05 3.3 9.386e-05 3.3 9.396e-05 0 9.388e-05 0 9.398e-05 3.3 9.389999999999999e-05 3.3 9.4e-05 0 9.392e-05 0 9.402e-05 3.3 9.394e-05 3.3 9.404e-05 0 9.396e-05 0 9.406e-05 3.3 9.397999999999999e-05 3.3 9.408e-05 0 9.4e-05 0 9.41e-05 3.3 9.402e-05 3.3 9.412e-05 0 9.404e-05 0 9.414e-05 3.3 9.405999999999999e-05 3.3 9.415999999999999e-05 0 9.408e-05 0 9.418e-05 3.3 9.41e-05 3.3 9.42e-05 0 9.412e-05 0 9.422e-05 3.3 9.413999999999999e-05 3.3 9.423999999999999e-05 0 9.415999999999999e-05 0 9.426e-05 3.3 9.418e-05 3.3 9.428e-05 0 9.42e-05 0 9.43e-05 3.3 9.421999999999999e-05 3.3 9.431999999999999e-05 0 9.423999999999999e-05 0 9.434e-05 3.3 9.426e-05 3.3 9.436e-05 0 9.428e-05 0 9.438e-05 3.3 9.43e-05 3.3 9.44e-05 0 9.431999999999999e-05 0 9.442e-05 3.3 9.434e-05 3.3 9.444e-05 0 9.436e-05 0 9.446e-05 3.3 9.438e-05 3.3 9.448e-05 0 9.439999999999999e-05 0 9.449999999999999e-05 3.3 9.442e-05 3.3 9.452e-05 0 9.444e-05 0 9.454e-05 3.3 9.446e-05 3.3 9.456e-05 0 9.447999999999999e-05 0 9.457999999999999e-05 3.3 9.449999999999999e-05 3.3 9.46e-05 0 9.452e-05 0 9.462e-05 3.3 9.454e-05 3.3 9.464e-05 0 9.455999999999999e-05 0 9.465999999999999e-05 3.3 9.457999999999999e-05 3.3 9.468e-05 0 9.46e-05 0 9.47e-05 3.3 9.462e-05 3.3 9.472e-05 0 9.464e-05 0 9.474e-05 3.3 9.465999999999999e-05 3.3 9.476e-05 0 9.468e-05 0 9.478e-05 3.3 9.47e-05 3.3 9.48e-05 0 9.472e-05 0 9.482e-05 3.3 9.473999999999999e-05 3.3 9.483999999999999e-05 0 9.476e-05 0 9.486e-05 3.3 9.478e-05 3.3 9.488e-05 0 9.48e-05 0 9.49e-05 3.3 9.481999999999999e-05 3.3 9.491999999999999e-05 0 9.483999999999999e-05 0 9.494e-05 3.3 9.486e-05 3.3 9.496e-05 0 9.488e-05 0 9.498e-05 3.3 9.489999999999999e-05 3.3 9.499999999999999e-05 0 9.491999999999999e-05 0 9.502e-05 3.3 9.494e-05 3.3 9.504e-05 0 9.496e-05 0 9.506e-05 3.3 9.498e-05 3.3 9.508e-05 0 9.499999999999999e-05 0 9.51e-05 3.3 9.502e-05 3.3 9.512e-05 0 9.504e-05 0 9.514e-05 3.3 9.506e-05 3.3 9.516e-05 0 9.507999999999999e-05 0 9.518e-05 3.3 9.51e-05 3.3 9.52e-05 0 9.512e-05 0 9.522e-05 3.3 9.514e-05 3.3 9.524e-05 0 9.515999999999999e-05 0 9.525999999999999e-05 3.3 9.518e-05 3.3 9.528e-05 0 9.52e-05 0 9.53e-05 3.3 9.522e-05 3.3 9.532e-05 0 9.523999999999999e-05 0 9.533999999999999e-05 3.3 9.525999999999999e-05 3.3 9.536e-05 0 9.528e-05 0 9.538e-05 3.3 9.53e-05 3.3 9.54e-05 0 9.532e-05 0 9.542e-05 3.3 9.533999999999999e-05 3.3 9.544e-05 0 9.536e-05 0 9.546e-05 3.3 9.538e-05 3.3 9.548e-05 0 9.54e-05 0 9.55e-05 3.3 9.541999999999999e-05 3.3 9.552e-05 0 9.544e-05 0 9.554e-05 3.3 9.546e-05 3.3 9.556e-05 0 9.548e-05 0 9.558e-05 3.3 9.549999999999999e-05 3.3 9.559999999999999e-05 0 9.552e-05 0 9.562e-05 3.3 9.554e-05 3.3 9.564e-05 0 9.556e-05 0 9.566e-05 3.3 9.557999999999999e-05 3.3 9.567999999999999e-05 0 9.559999999999999e-05 0 9.57e-05 3.3 9.562e-05 3.3 9.572e-05 0 9.564e-05 0 9.574e-05 3.3 9.566e-05 3.3 9.576e-05 0 9.567999999999999e-05 0 9.578e-05 3.3 9.57e-05 3.3 9.58e-05 0 9.572e-05 0 9.582e-05 3.3 9.574e-05 3.3 9.584e-05 0 9.575999999999999e-05 0 9.586e-05 3.3 9.578e-05 3.3 9.588e-05 0 9.58e-05 0 9.59e-05 3.3 9.582e-05 3.3 9.592e-05 0 9.583999999999999e-05 0 9.593999999999999e-05 3.3 9.586e-05 3.3 9.596e-05 0 9.588e-05 0 9.598e-05 3.3 9.59e-05 3.3 9.6e-05 0 9.591999999999999e-05 0 9.601999999999999e-05 3.3 9.593999999999999e-05 3.3 9.604e-05 0 9.596e-05 0 9.606e-05 3.3 9.598e-05 3.3 9.608e-05 0 9.599999999999999e-05 0 9.609999999999999e-05 3.3 9.601999999999999e-05 3.3 9.612e-05 0 9.604e-05 0 9.614e-05 3.3 9.606e-05 3.3 9.616e-05 0 9.608e-05 0 9.618e-05 3.3 9.609999999999999e-05 3.3 9.62e-05 0 9.612e-05 0 9.622e-05 3.3 9.614e-05 3.3 9.624e-05 0 9.616e-05 0 9.626e-05 3.3 9.617999999999999e-05 3.3 9.627999999999999e-05 0 9.62e-05 0 9.63e-05 3.3 9.622e-05 3.3 9.632e-05 0 9.624e-05 0 9.634e-05 3.3 9.625999999999999e-05 3.3 9.635999999999999e-05 0 9.627999999999999e-05 0 9.638e-05 3.3 9.63e-05 3.3 9.64e-05 0 9.632e-05 0 9.642e-05 3.3 9.633999999999999e-05 3.3 9.643999999999999e-05 0 9.635999999999999e-05 0 9.646e-05 3.3 9.638e-05 3.3 9.648e-05 0 9.64e-05 0 9.65e-05 3.3 9.642e-05 3.3 9.652e-05 0 9.643999999999999e-05 0 9.654e-05 3.3 9.646e-05 3.3 9.656e-05 0 9.648e-05 0 9.658e-05 3.3 9.65e-05 3.3 9.66e-05 0 9.651999999999999e-05 0 9.661999999999999e-05 3.3 9.654e-05 3.3 9.664e-05 0 9.656e-05 0 9.666e-05 3.3 9.658e-05 3.3 9.668e-05 0 9.659999999999999e-05 0 9.669999999999999e-05 3.3 9.661999999999999e-05 3.3 9.672e-05 0 9.664e-05 0 9.674e-05 3.3 9.666e-05 3.3 9.676e-05 0 9.667999999999999e-05 0 9.677999999999999e-05 3.3 9.669999999999999e-05 3.3 9.68e-05 0 9.672e-05 0 9.682e-05 3.3 9.674e-05 3.3 9.684e-05 0 9.676e-05 0 9.686e-05 3.3 9.677999999999999e-05 3.3 9.688e-05 0 9.68e-05 0 9.69e-05 3.3 9.682e-05 3.3 9.692e-05 0 9.684e-05 0 9.694e-05 3.3 9.685999999999999e-05 3.3 9.696e-05 0 9.688e-05 0 9.698e-05 3.3 9.69e-05 3.3 9.7e-05 0 9.692e-05 0 9.702e-05 3.3 9.693999999999999e-05 3.3 9.703999999999999e-05 0 9.696e-05 0 9.706e-05 3.3 9.698e-05 3.3 9.708e-05 0 9.7e-05 0 9.71e-05 3.3 9.701999999999999e-05 3.3 9.711999999999999e-05 0 9.703999999999999e-05 0 9.714e-05 3.3 9.706e-05 3.3 9.716e-05 0 9.708e-05 0 9.718e-05 3.3 9.71e-05 3.3 9.72e-05 0 9.711999999999999e-05 0 9.722e-05 3.3 9.714e-05 3.3 9.724e-05 0 9.716e-05 0 9.726e-05 3.3 9.718e-05 3.3 9.728e-05 0 9.719999999999999e-05 0 9.73e-05 3.3 9.722e-05 3.3 9.732e-05 0 9.724e-05 0 9.734e-05 3.3 9.726e-05 3.3 9.736e-05 0 9.727999999999999e-05 0 9.737999999999999e-05 3.3 9.73e-05 3.3 9.74e-05 0 9.732e-05 0 9.742e-05 3.3 9.734e-05 3.3 9.744e-05 0 9.735999999999999e-05 0 9.745999999999999e-05 3.3 9.737999999999999e-05 3.3 9.748e-05 0 9.74e-05 0 9.75e-05 3.3 9.742e-05 3.3 9.752e-05 0 9.744e-05 0 9.754e-05 3.3 9.745999999999999e-05 3.3 9.756e-05 0 9.748e-05 0 9.758e-05 3.3 9.75e-05 3.3 9.76e-05 0 9.752e-05 0 9.762e-05 3.3 9.753999999999999e-05 3.3 9.764e-05 0 9.756e-05 0 9.766e-05 3.3 9.758e-05 3.3 9.768e-05 0 9.76e-05 0 9.77e-05 3.3 9.761999999999999e-05 3.3 9.771999999999999e-05 0 9.764e-05 0 9.774e-05 3.3 9.766e-05 3.3 9.776e-05 0 9.768e-05 0 9.778e-05 3.3 9.769999999999999e-05 3.3 9.779999999999999e-05 0 9.771999999999999e-05 0 9.782e-05 3.3 9.774e-05 3.3 9.784e-05 0 9.776e-05 0 9.786e-05 3.3 9.778e-05 3.3 9.788e-05 0 9.779999999999999e-05 0 9.79e-05 3.3 9.782e-05 3.3 9.792e-05 0 9.784e-05 0 9.794e-05 3.3 9.786e-05 3.3 9.796e-05 0 9.787999999999999e-05 0 9.798e-05 3.3 9.79e-05 3.3 9.8e-05 0 9.792e-05 0 9.802e-05 3.3 9.794e-05 3.3 9.804e-05 0 9.795999999999999e-05 0 9.805999999999999e-05 3.3 9.798e-05 3.3 9.808e-05 0 9.8e-05 0 9.81e-05 3.3 9.802e-05 3.3 9.812e-05 0 9.803999999999999e-05 0 9.813999999999999e-05 3.3 9.805999999999999e-05 3.3 9.816e-05 0 9.808e-05 0 9.818e-05 3.3 9.81e-05 3.3 9.82e-05 0 9.811999999999999e-05 0 9.821999999999999e-05 3.3 9.813999999999999e-05 3.3 9.824e-05 0 9.816e-05 0 9.826e-05 3.3 9.818e-05 3.3 9.828e-05 0 9.82e-05 0 9.83e-05 3.3 9.821999999999999e-05 3.3 9.832e-05 0 9.824e-05 0 9.834e-05 3.3 9.826e-05 3.3 9.836e-05 0 9.828e-05 0 9.838e-05 3.3 9.829999999999999e-05 3.3 9.839999999999999e-05 0 9.832e-05 0 9.842e-05 3.3 9.834e-05 3.3 9.844e-05 0 9.836e-05 0 9.846e-05 3.3 9.837999999999999e-05 3.3 9.847999999999999e-05 0 9.839999999999999e-05 0 9.85e-05 3.3 9.842e-05 3.3 9.852e-05 0 9.844e-05 0 9.854e-05 3.3 9.845999999999999e-05 3.3 9.855999999999999e-05 0 9.847999999999999e-05 0 9.858e-05 3.3 9.85e-05 3.3 9.86e-05 0 9.852e-05 0 9.862e-05 3.3 9.854e-05 3.3 9.864e-05 0 9.855999999999999e-05 0 9.866e-05 3.3 9.858e-05 3.3 9.868e-05 0 9.86e-05 0 9.87e-05 3.3 9.862e-05 3.3 9.872e-05 0 9.863999999999999e-05 0 9.873999999999999e-05 3.3 9.866e-05 3.3 9.876e-05 0 9.868e-05 0 9.878e-05 3.3 9.87e-05 3.3 9.88e-05 0 9.871999999999999e-05 0 9.881999999999999e-05 3.3 9.873999999999999e-05 3.3 9.884e-05 0 9.876e-05 0 9.886e-05 3.3 9.878e-05 3.3 9.888e-05 0 9.879999999999999e-05 0 9.889999999999999e-05 3.3 9.881999999999999e-05 3.3 9.892e-05 0 9.884e-05 0 9.894e-05 3.3 9.886e-05 3.3 9.896e-05 0 9.888e-05 0 9.898e-05 3.3 9.889999999999999e-05 3.3 9.9e-05 0 9.892e-05 0 9.902e-05 3.3 9.894e-05 3.3 9.904e-05 0 9.896e-05 0 9.906e-05 3.3 9.897999999999999e-05 3.3 9.908e-05 0 9.9e-05 0 9.91e-05 3.3 9.902e-05 3.3 9.912e-05 0 9.904e-05 0 9.914e-05 3.3 9.905999999999999e-05 3.3 9.915999999999999e-05 0 9.908e-05 0 9.918e-05 3.3 9.91e-05 3.3 9.92e-05 0 9.912e-05 0 9.922e-05 3.3 9.913999999999999e-05 3.3 9.923999999999999e-05 0 9.915999999999999e-05 0 9.926e-05 3.3 9.918e-05 3.3 9.928e-05 0 9.92e-05 0 9.93e-05 3.3 9.922e-05 3.3 9.932e-05 0 9.923999999999999e-05 0 9.934e-05 3.3 9.926e-05 3.3 9.936e-05 0 9.928e-05 0 9.938e-05 3.3 9.93e-05 3.3 9.94e-05 0 9.931999999999999e-05 0 9.942e-05 3.3 9.934e-05 3.3 9.944e-05 0 9.936e-05 0 9.946e-05 3.3 9.938e-05 3.3 9.948e-05 0 9.939999999999999e-05 0 9.949999999999999e-05 3.3 9.942e-05 3.3 9.952e-05 0 9.944e-05 0 9.954e-05 3.3 9.946e-05 3.3 9.956e-05 0 9.947999999999999e-05 0 9.957999999999999e-05 3.3 9.949999999999999e-05 3.3 9.96e-05 0 9.952e-05 0 9.962e-05 3.3 9.954e-05 3.3 9.964e-05 0 9.956e-05 0 9.966e-05 3.3 9.957999999999999e-05 3.3 9.968e-05 0 9.96e-05 0 9.97e-05 3.3 9.962e-05 3.3 9.972e-05 0 9.964e-05 0 9.974e-05 3.3 9.965999999999999e-05 3.3 9.976e-05 0 9.968e-05 0 9.978e-05 3.3 9.97e-05 3.3 9.98e-05 0 9.972e-05 0 9.982e-05 3.3 9.973999999999999e-05 3.3 9.983999999999999e-05 0 9.976e-05 0 9.986e-05 3.3 9.978e-05 3.3 9.988e-05 0 9.98e-05 0 9.99e-05 3.3 9.981999999999999e-05 3.3 9.991999999999999e-05 0 9.983999999999999e-05 0 9.994e-05 3.3 9.986e-05 3.3 9.996e-05 0 9.988e-05 0 9.998e-05 3.3 9.989999999999999e-05 3.3 9.999999999999999e-05 0 9.991999999999999e-05 0 0.00010002 3.3 9.994e-05 3.3 0.00010004 0 9.996e-05 0 0.00010006 3.3 9.998e-05 3.3 0.00010008 0 9.999999999999999e-05 0 0.0001001 3.3 0.00010002 3.3 0.00010012 0 0.00010004 0 0.00010014 3.3 0.00010006 3.3 0.00010016 0 0.00010007999999999999 0 0.00010017999999999999 3.3 0.0001001 3.3 0.0001002 0 0.00010012 0 0.00010022 3.3 0.00010014 3.3 0.00010024 0 0.00010015999999999999 0 0.00010025999999999999 3.3 0.00010017999999999999 3.3 0.00010028 0 0.0001002 0 0.0001003 3.3 0.00010022 3.3 0.00010032 0 0.00010023999999999999 0 0.00010033999999999999 3.3 0.00010025999999999999 3.3 0.00010036 0 0.00010028 0 0.00010038 3.3 0.0001003 3.3 0.0001004 0 0.00010032 0 0.00010042 3.3 0.00010033999999999999 3.3 0.00010044 0 0.00010036 0 0.00010046 3.3 0.00010038 3.3 0.00010048 0 0.0001004 0 0.0001005 3.3 0.00010041999999999999 3.3 0.00010051999999999999 0 0.00010044 0 0.00010054 3.3 0.00010046 3.3 0.00010056 0 0.00010048 0 0.00010058 3.3 0.00010049999999999999 3.3 0.00010059999999999999 0 0.00010051999999999999 0 0.00010062 3.3 0.00010054 3.3 0.00010064 0 0.00010056 0 0.00010066 3.3 0.00010057999999999999 3.3 0.00010067999999999999 0 0.00010059999999999999 0 0.0001007 3.3 0.00010062 3.3 0.00010072 0 0.00010064 0 0.00010074 3.3 0.00010066 3.3 0.00010076 0 0.00010067999999999999 0 0.00010078 3.3 0.0001007 3.3 0.0001008 0 0.00010072 0 0.00010082 3.3 0.00010074 3.3 0.00010084 0 0.00010075999999999999 0 0.00010085999999999999 3.3 0.00010078 3.3 0.00010088 0 0.0001008 0 0.0001009 3.3 0.00010082 3.3 0.00010092 0 0.00010083999999999999 0 0.00010093999999999999 3.3 0.00010085999999999999 3.3 0.00010096 0 0.00010088 0 0.00010098 3.3 0.0001009 3.3 0.000101 0 0.00010091999999999999 0 0.00010101999999999999 3.3 0.00010093999999999999 3.3 0.00010104 0 0.00010096 0 0.00010106 3.3 0.00010098 3.3 0.00010108 0 0.000101 0 0.0001011 3.3 0.00010101999999999999 3.3 0.00010112 0 0.00010104 0 0.00010114 3.3 0.00010106 3.3 0.00010116 0 0.00010108 0 0.00010118 3.3 0.00010109999999999999 3.3 0.0001012 0 0.00010112 0 0.00010122 3.3 0.00010114 3.3 0.00010124 0 0.00010116 0 0.00010126 3.3 0.00010117999999999999 3.3 0.00010127999999999999 0 0.0001012 0 0.0001013 3.3 0.00010122 3.3 0.00010132 0 0.00010124 0 0.00010134 3.3 0.00010125999999999999 3.3 0.00010135999999999999 0 0.00010127999999999999 0 0.00010138 3.3 0.0001013 3.3 0.0001014 0 0.00010132 0 0.00010142 3.3 0.00010134 3.3 0.00010144 0 0.00010135999999999999 0 0.00010146 3.3 0.00010138 3.3 0.00010148 0 0.0001014 0 0.0001015 3.3 0.00010142 3.3 0.00010152 0 0.00010143999999999999 0 0.00010154 3.3 0.00010146 3.3 0.00010156 0 0.00010148 0 0.00010158 3.3 0.0001015 3.3 0.0001016 0 0.00010151999999999999 0 0.00010161999999999999 3.3 0.00010154 3.3 0.00010164 0 0.00010156 0 0.00010166 3.3 0.00010158 3.3 0.00010168 0 0.00010159999999999999 0 0.00010169999999999999 3.3 0.00010161999999999999 3.3 0.00010172 0 0.00010164 0 0.00010174 3.3 0.00010166 3.3 0.00010176 0 0.00010168 0 0.00010178 3.3 0.00010169999999999999 3.3 0.0001018 0 0.00010172 0 0.00010182 3.3 0.00010174 3.3 0.00010184 0 0.00010176 0 0.00010186 3.3 0.00010177999999999999 3.3 0.00010188 0 0.0001018 0 0.0001019 3.3 0.00010182 3.3 0.00010192 0 0.00010184 0 0.00010194 3.3 0.00010185999999999999 3.3 0.00010195999999999999 0 0.00010188 0 0.00010198 3.3 0.0001019 3.3 0.000102 0 0.00010192 0 0.00010202 3.3 0.00010193999999999999 3.3 0.00010203999999999999 0 0.00010195999999999999 0 0.00010206 3.3 0.00010198 3.3 0.00010208 0 0.000102 0 0.0001021 3.3 0.00010201999999999999 3.3 0.00010211999999999999 0 0.00010203999999999999 0 0.00010214 3.3 0.00010206 3.3 0.00010216 0 0.00010208 0 0.00010218 3.3 0.0001021 3.3 0.0001022 0 0.00010211999999999999 0 0.00010222 3.3 0.00010214 3.3 0.00010224 0 0.00010216 0 0.00010226 3.3 0.00010218 3.3 0.00010228 0 0.00010219999999999999 0 0.00010229999999999999 3.3 0.00010222 3.3 0.00010232 0 0.00010224 0 0.00010234 3.3 0.00010226 3.3 0.00010236 0 0.00010227999999999999 0 0.00010237999999999999 3.3 0.00010229999999999999 3.3 0.0001024 0 0.00010232 0 0.00010242 3.3 0.00010234 3.3 0.00010244 0 0.00010235999999999999 0 0.00010245999999999999 3.3 0.00010237999999999999 3.3 0.00010248 0 0.0001024 0 0.0001025 3.3 0.00010242 3.3 0.00010252 0 0.00010244 0 0.00010254 3.3 0.00010245999999999999 3.3 0.00010256 0 0.00010248 0 0.00010258 3.3 0.0001025 3.3 0.0001026 0 0.00010252 0 0.00010262 3.3 0.00010253999999999999 3.3 0.00010263999999999999 0 0.00010256 0 0.00010266 3.3 0.00010258 3.3 0.00010268 0 0.0001026 0 0.0001027 3.3 0.00010261999999999999 3.3 0.00010271999999999999 0 0.00010263999999999999 0 0.00010274 3.3 0.00010266 3.3 0.00010276 0 0.00010268 0 0.00010278 3.3 0.00010269999999999999 3.3 0.00010279999999999999 0 0.00010271999999999999 0 0.00010282 3.3 0.00010274 3.3 0.00010284 0 0.00010276 0 0.00010286 3.3 0.00010278 3.3 0.00010288 0 0.00010279999999999999 0 0.0001029 3.3 0.00010282 3.3 0.00010292 0 0.00010284 0 0.00010294 3.3 0.00010286 3.3 0.00010296 0 0.00010287999999999999 0 0.00010297999999999999 3.3 0.0001029 3.3 0.000103 0 0.00010292 0 0.00010302 3.3 0.00010294 3.3 0.00010304 0 0.00010295999999999999 0 0.00010305999999999999 3.3 0.00010297999999999999 3.3 0.00010308 0 0.000103 0 0.0001031 3.3 0.00010302 3.3 0.00010312 0 0.00010303999999999999 0 0.00010313999999999999 3.3 0.00010305999999999999 3.3 0.00010316 0 0.00010308 0 0.00010318 3.3 0.0001031 3.3 0.0001032 0 0.00010312 0 0.00010322 3.3 0.00010313999999999999 3.3 0.00010324 0 0.00010316 0 0.00010326 3.3 0.00010318 3.3 0.00010328 0 0.0001032 0 0.0001033 3.3 0.00010321999999999999 3.3 0.00010332 0 0.00010324 0 0.00010334 3.3 0.00010326 3.3 0.00010336 0 0.00010328 0 0.00010338 3.3 0.00010329999999999999 3.3 0.00010339999999999999 0 0.00010332 0 0.00010342 3.3 0.00010334 3.3 0.00010344 0 0.00010336 0 0.00010346 3.3 0.00010337999999999999 3.3 0.00010347999999999999 0 0.00010339999999999999 0 0.0001035 3.3 0.00010342 3.3 0.00010352 0 0.00010344 0 0.00010354 3.3 0.00010346 3.3 0.00010356 0 0.00010347999999999999 0 0.00010358 3.3 0.0001035 3.3 0.0001036 0 0.00010352 0 0.00010362 3.3 0.00010354 3.3 0.00010364 0 0.00010355999999999999 0 0.00010366 3.3 0.00010358 3.3 0.00010368 0 0.0001036 0 0.0001037 3.3 0.00010362 3.3 0.00010372 0 0.00010363999999999999 0 0.00010373999999999999 3.3 0.00010366 3.3 0.00010376 0 0.00010368 0 0.00010378 3.3 0.0001037 3.3 0.0001038 0 0.00010371999999999999 0 0.00010381999999999999 3.3 0.00010373999999999999 3.3 0.00010384 0 0.00010376 0 0.00010386 3.3 0.00010378 3.3 0.00010388 0 0.00010379999999999999 0 0.00010389999999999999 3.3 0.00010381999999999999 3.3 0.00010392 0 0.00010384 0 0.00010394 3.3 0.00010386 3.3 0.00010396 0 0.00010388 0 0.00010398 3.3 0.00010389999999999999 3.3 0.000104 0 0.00010392 0 0.00010402 3.3 0.00010394 3.3 0.00010404 0 0.00010396 0 0.00010406 3.3 0.00010397999999999999 3.3 0.00010407999999999999 0 0.000104 0 0.0001041 3.3 0.00010402 3.3 0.00010412 0 0.00010404 0 0.00010414 3.3 0.00010405999999999999 3.3 0.00010415999999999999 0 0.00010407999999999999 0 0.00010418 3.3 0.0001041 3.3 0.0001042 0 0.00010412 0 0.00010422 3.3 0.00010413999999999999 3.3 0.00010423999999999999 0 0.00010415999999999999 0 0.00010426 3.3 0.00010418 3.3 0.00010428 0 0.0001042 0 0.0001043 3.3 0.00010422 3.3 0.00010432 0 0.00010423999999999999 0 0.00010434 3.3 0.00010426 3.3 0.00010436 0 0.00010428 0 0.00010438 3.3 0.0001043 3.3 0.0001044 0 0.00010431999999999999 0 0.00010441999999999999 3.3 0.00010434 3.3 0.00010444 0 0.00010436 0 0.00010446 3.3 0.00010438 3.3 0.00010448 0 0.00010439999999999999 0 0.00010449999999999999 3.3 0.00010441999999999999 3.3 0.00010452 0 0.00010444 0 0.00010454 3.3 0.00010446 3.3 0.00010456 0 0.00010447999999999999 0 0.00010457999999999999 3.3 0.00010449999999999999 3.3 0.0001046 0 0.00010452 0 0.00010462 3.3 0.00010454 3.3 0.00010464 0 0.00010456 0 0.00010466 3.3 0.00010457999999999999 3.3 0.00010468 0 0.0001046 0 0.0001047 3.3 0.00010462 3.3 0.00010472 0 0.00010464 0 0.00010474 3.3 0.00010465999999999999 3.3 0.00010475999999999999 0 0.00010468 0 0.00010478 3.3 0.0001047 3.3 0.0001048 0 0.00010472 0 0.00010482 3.3 0.00010473999999999999 3.3 0.00010483999999999999 0 0.00010475999999999999 0 0.00010486 3.3 0.00010478 3.3 0.00010488 0 0.0001048 0 0.0001049 3.3 0.00010481999999999999 3.3 0.00010491999999999999 0 0.00010483999999999999 0 0.00010494 3.3 0.00010486 3.3 0.00010496 0 0.00010488 0 0.00010498 3.3 0.0001049 3.3 0.000105 0 0.00010491999999999999 0 0.00010502 3.3 0.00010494 3.3 0.00010504 0 0.00010496 0 0.00010506 3.3 0.00010498 3.3 0.00010508 0 0.00010499999999999999 0 0.0001051 3.3 0.00010502 3.3 0.00010512 0 0.00010504 0 0.00010514 3.3 0.00010506 3.3 0.00010516 0 0.00010507999999999999 0 0.00010517999999999999 3.3 0.0001051 3.3 0.0001052 0 0.00010512 0 0.00010522 3.3 0.00010514 3.3 0.00010524 0 0.00010515999999999999 0 0.00010525999999999999 3.3 0.00010517999999999999 3.3 0.00010528 0 0.0001052 0 0.0001053 3.3 0.00010522 3.3 0.00010532 0 0.00010524 0 0.00010534 3.3 0.00010525999999999999 3.3 0.00010536 0 0.00010528 0 0.00010538 3.3 0.0001053 3.3 0.0001054 0 0.00010532 0 0.00010542 3.3 0.00010533999999999999 3.3 0.00010544 0 0.00010536 0 0.00010546 3.3 0.00010538 3.3 0.00010548 0 0.0001054 0 0.0001055 3.3 0.00010541999999999999 3.3 0.00010551999999999999 0 0.00010544 0 0.00010554 3.3 0.00010546 3.3 0.00010556 0 0.00010548 0 0.00010558 3.3 0.00010549999999999999 3.3 0.00010559999999999999 0 0.00010551999999999999 0 0.00010562 3.3 0.00010554 3.3 0.00010564 0 0.00010556 0 0.00010566 3.3 0.00010558 3.3 0.00010568 0 0.00010559999999999999 0 0.0001057 3.3 0.00010562 3.3 0.00010572 0 0.00010564 0 0.00010574 3.3 0.00010566 3.3 0.00010576 0 0.00010567999999999999 0 0.00010578 3.3 0.0001057 3.3 0.0001058 0 0.00010572 0 0.00010582 3.3 0.00010574 3.3 0.00010584 0 0.00010575999999999999 0 0.00010585999999999999 3.3 0.00010578 3.3 0.00010588 0 0.0001058 0 0.0001059 3.3 0.00010582 3.3 0.00010592 0 0.00010583999999999999 0 0.00010593999999999999 3.3 0.00010585999999999999 3.3 0.00010596 0 0.00010588 0 0.00010598 3.3 0.0001059 3.3 0.000106 0 0.00010591999999999999 0 0.00010601999999999999 3.3 0.00010593999999999999 3.3 0.00010604 0 0.00010596 0 0.00010606 3.3 0.00010598 3.3 0.00010608 0 0.000106 0 0.0001061 3.3 0.00010601999999999999 3.3 0.00010612 0 0.00010604 0 0.00010614 3.3 0.00010606 3.3 0.00010616 0 0.00010608 0 0.00010618 3.3 0.00010609999999999999 3.3 0.00010619999999999999 0 0.00010612 0 0.00010622 3.3 0.00010614 3.3 0.00010624 0 0.00010616 0 0.00010626 3.3 0.00010617999999999999 3.3 0.00010627999999999999 0 0.00010619999999999999 0 0.0001063 3.3 0.00010622 3.3 0.00010632 0 0.00010624 0 0.00010634 3.3 0.00010625999999999999 3.3 0.00010635999999999999 0 0.00010627999999999999 0 0.00010638 3.3 0.0001063 3.3 0.0001064 0 0.00010632 0 0.00010642 3.3 0.00010634 3.3 0.00010644 0 0.00010635999999999999 0 0.00010646 3.3 0.00010638 3.3 0.00010648 0 0.0001064 0 0.0001065 3.3 0.00010642 3.3 0.00010652 0 0.00010643999999999999 0 0.00010653999999999999 3.3 0.00010646 3.3 0.00010656 0 0.00010648 0 0.00010658 3.3 0.0001065 3.3 0.0001066 0 0.00010651999999999999 0 0.00010661999999999999 3.3 0.00010653999999999999 3.3 0.00010664 0 0.00010656 0 0.00010666 3.3 0.00010658 3.3 0.00010668 0 0.00010659999999999999 0 0.00010669999999999999 3.3 0.00010661999999999999 3.3 0.00010672 0 0.00010664 0 0.00010674 3.3 0.00010666 3.3 0.00010676 0 0.00010668 0 0.00010678 3.3 0.00010669999999999999 3.3 0.0001068 0 0.00010672 0 0.00010682 3.3 0.00010674 3.3 0.00010684 0 0.00010676 0 0.00010686 3.3 0.00010677999999999999 3.3 0.00010687999999999999 0 0.0001068 0 0.0001069 3.3 0.00010682 3.3 0.00010692 0 0.00010684 0 0.00010694 3.3 0.00010685999999999999 3.3 0.00010695999999999999 0 0.00010687999999999999 0 0.00010698 3.3 0.0001069 3.3 0.000107 0 0.00010692 0 0.00010702 3.3 0.00010693999999999999 3.3 0.00010703999999999999 0 0.00010695999999999999 0 0.00010706 3.3 0.00010698 3.3 0.00010708 0 0.000107 0 0.0001071 3.3 0.00010702 3.3 0.00010712 0 0.00010703999999999999 0 0.00010714 3.3 0.00010706 3.3 0.00010716 0 0.00010708 0 0.00010718 3.3 0.0001071 3.3 0.0001072 0 0.00010711999999999999 0 0.00010722 3.3 0.00010714 3.3 0.00010724 0 0.00010716 0 0.00010726 3.3 0.00010718 3.3 0.00010728 0 0.00010719999999999999 0 0.00010729999999999999 3.3 0.00010722 3.3 0.00010732 0 0.00010724 0 0.00010734 3.3 0.00010726 3.3 0.00010736 0 0.00010727999999999999 0 0.00010737999999999999 3.3 0.00010729999999999999 3.3 0.0001074 0 0.00010732 0 0.00010742 3.3 0.00010734 3.3 0.00010744 0 0.00010736 0 0.00010746 3.3 0.00010737999999999999 3.3 0.00010748 0 0.0001074 0 0.0001075 3.3 0.00010742 3.3 0.00010752 0 0.00010744 0 0.00010754 3.3 0.00010745999999999999 3.3 0.00010756 0 0.00010748 0 0.00010758 3.3 0.0001075 3.3 0.0001076 0 0.00010752 0 0.00010762 3.3 0.00010753999999999999 3.3 0.00010763999999999999 0 0.00010756 0 0.00010766 3.3 0.00010758 3.3 0.00010768 0 0.0001076 0 0.0001077 3.3 0.00010761999999999999 3.3 0.00010771999999999999 0 0.00010763999999999999 0 0.00010774 3.3 0.00010766 3.3 0.00010776 0 0.00010768 0 0.00010778 3.3 0.00010769999999999999 3.3 0.00010779999999999999 0 0.00010771999999999999 0 0.00010782 3.3 0.00010774 3.3 0.00010784 0 0.00010776 0 0.00010786 3.3 0.00010778 3.3 0.00010788 0 0.00010779999999999999 0 0.0001079 3.3 0.00010782 3.3 0.00010792 0 0.00010784 0 0.00010794 3.3 0.00010786 3.3 0.00010796 0 0.00010787999999999999 0 0.00010797999999999999 3.3 0.0001079 3.3 0.000108 0 0.00010792 0 0.00010802 3.3 0.00010794 3.3 0.00010804 0 0.00010795999999999999 0 0.00010805999999999999 3.3 0.00010797999999999999 3.3 0.00010808 0 0.000108 0 0.0001081 3.3 0.00010802 3.3 0.00010812 0 0.00010803999999999999 0 0.00010813999999999999 3.3 0.00010805999999999999 3.3 0.00010816 0 0.00010808 0 0.00010818 3.3 0.0001081 3.3 0.0001082 0 0.00010812 0 0.00010822 3.3 0.00010813999999999999 3.3 0.00010824 0 0.00010816 0 0.00010826 3.3 0.00010818 3.3 0.00010828 0 0.0001082 0 0.0001083 3.3 0.00010821999999999999 3.3 0.00010831999999999999 0 0.00010824 0 0.00010834 3.3 0.00010826 3.3 0.00010836 0 0.00010828 0 0.00010838 3.3 0.00010829999999999999 3.3 0.00010839999999999999 0 0.00010831999999999999 0 0.00010842 3.3 0.00010834 3.3 0.00010844 0 0.00010836 0 0.00010846 3.3 0.00010837999999999999 3.3 0.00010847999999999999 0 0.00010839999999999999 0 0.0001085 3.3 0.00010842 3.3 0.00010852 0 0.00010844 0 0.00010854 3.3 0.00010846 3.3 0.00010856 0 0.00010847999999999999 0 0.00010858 3.3 0.0001085 3.3 0.0001086 0 0.00010852 0 0.00010862 3.3 0.00010854 3.3 0.00010864 0 0.00010855999999999999 0 0.00010865999999999999 3.3 0.00010858 3.3 0.00010868 0 0.0001086 0 0.0001087 3.3 0.00010862 3.3 0.00010872 0 0.00010863999999999999 0 0.00010873999999999999 3.3 0.00010865999999999999 3.3 0.00010876 0 0.00010868 0 0.00010878 3.3 0.0001087 3.3 0.0001088 0 0.00010871999999999999 0 0.00010881999999999999 3.3 0.00010873999999999999 3.3 0.00010884 0 0.00010876 0 0.00010886 3.3 0.00010878 3.3 0.00010888 0 0.0001088 0 0.0001089 3.3 0.00010881999999999999 3.3 0.00010892 0 0.00010884 0 0.00010894 3.3 0.00010886 3.3 0.00010896 0 0.00010888 0 0.00010898 3.3 0.00010889999999999999 3.3 0.00010899999999999999 0 0.00010892 0 0.00010902 3.3 0.00010894 3.3 0.00010904 0 0.00010896 0 0.00010906 3.3 0.00010897999999999999 3.3 0.00010907999999999999 0 0.00010899999999999999 0 0.0001091 3.3 0.00010902 3.3 0.00010912 0 0.00010904 0 0.00010914 3.3 0.00010905999999999999 3.3 0.00010915999999999999 0 0.00010907999999999999 0 0.00010918 3.3 0.0001091 3.3 0.0001092 0 0.00010912 0 0.00010922 3.3 0.00010914 3.3 0.00010924 0 0.00010915999999999999 0 0.00010926 3.3 0.00010918 3.3 0.00010928 0 0.0001092 0 0.0001093 3.3 0.00010922 3.3 0.00010932 0 0.00010923999999999999 0 0.00010934 3.3 0.00010926 3.3 0.00010936 0 0.00010928 0 0.00010938 3.3 0.0001093 3.3 0.0001094 0 0.00010931999999999999 0 0.00010941999999999999 3.3 0.00010934 3.3 0.00010944 0 0.00010936 0 0.00010946 3.3 0.00010938 3.3 0.00010948 0 0.00010939999999999999 0 0.00010949999999999999 3.3 0.00010941999999999999 3.3 0.00010952 0 0.00010944 0 0.00010954 3.3 0.00010946 3.3 0.00010956 0 0.00010948 0 0.00010958 3.3 0.00010949999999999999 3.3 0.0001096 0 0.00010952 0 0.00010962 3.3 0.00010954 3.3 0.00010964 0 0.00010956 0 0.00010966 3.3 0.00010957999999999999 3.3 0.00010968 0 0.0001096 0 0.0001097 3.3 0.00010962 3.3 0.00010972 0 0.00010964 0 0.00010974 3.3 0.00010965999999999999 3.3 0.00010975999999999999 0 0.00010968 0 0.00010978 3.3 0.0001097 3.3 0.0001098 0 0.00010972 0 0.00010982 3.3 0.00010973999999999999 3.3 0.00010983999999999999 0 0.00010975999999999999 0 0.00010986 3.3 0.00010978 3.3 0.00010988 0 0.0001098 0 0.0001099 3.3 0.00010981999999999999 3.3 0.00010991999999999999 0 0.00010983999999999999 0 0.00010994 3.3 0.00010986 3.3 0.00010996 0 0.00010988 0 0.00010998 3.3 0.0001099 3.3 0.00011 0 0.00010991999999999999 0 0.00011002 3.3 0.00010994 3.3 0.00011004 0 0.00010996 0 0.00011006 3.3 0.00010998 3.3 0.00011008 0 0.00010999999999999999 0 0.00011009999999999999 3.3 0.00011002 3.3 0.00011012 0 0.00011004 0 0.00011014 3.3 0.00011006 3.3 0.00011016 0 0.00011007999999999999 0 0.00011017999999999999 3.3 0.00011009999999999999 3.3 0.0001102 0 0.00011012 0 0.00011022 3.3 0.00011014 3.3 0.00011024 0 0.00011015999999999999 0 0.00011025999999999999 3.3 0.00011017999999999999 3.3 0.00011028 0 0.0001102 0 0.0001103 3.3 0.00011022 3.3 0.00011032 0 0.00011024 0 0.00011034 3.3 0.00011025999999999999 3.3 0.00011036 0 0.00011028 0 0.00011038 3.3 0.0001103 3.3 0.0001104 0 0.00011032 0 0.00011042 3.3 0.00011033999999999999 3.3 0.00011043999999999999 0 0.00011036 0 0.00011046 3.3 0.00011038 3.3 0.00011048 0 0.0001104 0 0.0001105 3.3 0.00011041999999999999 3.3 0.00011051999999999999 0 0.00011043999999999999 0 0.00011054 3.3 0.00011046 3.3 0.00011056 0 0.00011048 0 0.00011058 3.3 0.00011049999999999999 3.3 0.00011059999999999999 0 0.00011051999999999999 0 0.00011062 3.3 0.00011054 3.3 0.00011064 0 0.00011056 0 0.00011066 3.3 0.00011058 3.3 0.00011068 0 0.00011059999999999999 0 0.0001107 3.3 0.00011062 3.3 0.00011072 0 0.00011064 0 0.00011074 3.3 0.00011066 3.3 0.00011076 0 0.00011067999999999999 0 0.00011077999999999999 3.3 0.0001107 3.3 0.0001108 0 0.00011072 0 0.00011082 3.3 0.00011074 3.3 0.00011084 0 0.00011075999999999999 0 0.00011085999999999999 3.3 0.00011077999999999999 3.3 0.00011088 0 0.0001108 0 0.0001109 3.3 0.00011082 3.3 0.00011092 0 0.00011083999999999999 0 0.00011093999999999999 3.3 0.00011085999999999999 3.3 0.00011096 0 0.00011088 0 0.00011098 3.3 0.0001109 3.3 0.000111 0 0.00011092 0 0.00011102 3.3 0.00011093999999999999 3.3 0.00011104 0 0.00011096 0 0.00011106 3.3 0.00011098 3.3 0.00011108 0 0.000111 0 0.0001111 3.3 0.00011101999999999999 3.3 0.00011111999999999999 0 0.00011104 0 0.00011114 3.3 0.00011106 3.3 0.00011116 0 0.00011108 0 0.00011118 3.3 0.00011109999999999999 3.3 0.00011119999999999999 0 0.00011111999999999999 0 0.00011122 3.3 0.00011114 3.3 0.00011124 0 0.00011116 0 0.00011126 3.3 0.00011117999999999999 3.3 0.00011127999999999999 0 0.00011119999999999999 0 0.0001113 3.3 0.00011122 3.3 0.00011132 0 0.00011124 0 0.00011134 3.3 0.00011126 3.3 0.00011136 0 0.00011127999999999999 0 0.00011138 3.3 0.0001113 3.3 0.0001114 0 0.00011132 0 0.00011142 3.3 0.00011134 3.3 0.00011144 0 0.00011135999999999999 0 0.00011146 3.3 0.00011138 3.3 0.00011148 0 0.0001114 0 0.0001115 3.3 0.00011142 3.3 0.00011152 0 0.00011143999999999999 0 0.00011153999999999999 3.3 0.00011146 3.3 0.00011156 0 0.00011148 0 0.00011158 3.3 0.0001115 3.3 0.0001116 0 0.00011151999999999999 0 0.00011161999999999999 3.3 0.00011153999999999999 3.3 0.00011164 0 0.00011156 0 0.00011166 3.3 0.00011158 3.3 0.00011168 0 0.00011159999999999999 0 0.00011169999999999999 3.3 0.00011161999999999999 3.3 0.00011172 0 0.00011164 0 0.00011174 3.3 0.00011166 3.3 0.00011176 0 0.00011168 0 0.00011178 3.3 0.00011169999999999999 3.3 0.0001118 0 0.00011172 0 0.00011182 3.3 0.00011174 3.3 0.00011184 0 0.00011176 0 0.00011186 3.3 0.00011177999999999999 3.3 0.00011187999999999999 0 0.0001118 0 0.0001119 3.3 0.00011182 3.3 0.00011192 0 0.00011184 0 0.00011194 3.3 0.00011185999999999999 3.3 0.00011195999999999999 0 0.00011187999999999999 0 0.00011198 3.3 0.0001119 3.3 0.000112 0 0.00011192 0 0.00011202 3.3 0.00011193999999999999 3.3 0.00011203999999999999 0 0.00011195999999999999 0 0.00011206 3.3 0.00011198 3.3 0.00011208 0 0.000112 0 0.0001121 3.3 0.00011202 3.3 0.00011212 0 0.00011203999999999999 0 0.00011214 3.3 0.00011206 3.3 0.00011216 0 0.00011208 0 0.00011218 3.3 0.0001121 3.3 0.0001122 0 0.00011211999999999999 0 0.00011221999999999999 3.3 0.00011214 3.3 0.00011224 0 0.00011216 0 0.00011226 3.3 0.00011218 3.3 0.00011228 0 0.00011219999999999999 0 0.00011229999999999999 3.3 0.00011221999999999999 3.3 0.00011232 0 0.00011224 0 0.00011234 3.3 0.00011226 3.3 0.00011236 0 0.00011227999999999999 0 0.00011237999999999999 3.3 0.00011229999999999999 3.3 0.0001124 0 0.00011232 0 0.00011242 3.3 0.00011234 3.3 0.00011244 0 0.00011236 0 0.00011246 3.3 0.00011237999999999999 3.3 0.00011248 0 0.0001124 0 0.0001125 3.3 0.00011242 3.3 0.00011252 0 0.00011244 0 0.00011254 3.3 0.00011245999999999999 3.3 0.00011255999999999999 0 0.00011248 0 0.00011258 3.3 0.0001125 3.3 0.0001126 0 0.00011252 0 0.00011262 3.3 0.00011253999999999999 3.3 0.00011263999999999999 0 0.00011255999999999999 0 0.00011266 3.3 0.00011258 3.3 0.00011268 0 0.0001126 0 0.0001127 3.3 0.00011261999999999999 3.3 0.00011271999999999999 0 0.00011263999999999999 0 0.00011274 3.3 0.00011266 3.3 0.00011276 0 0.00011268 0 0.00011278 3.3 0.0001127 3.3 0.0001128 0 0.00011271999999999999 0 0.00011282 3.3 0.00011274 3.3 0.00011284 0 0.00011276 0 0.00011286 3.3 0.00011278 3.3 0.00011288 0 0.00011279999999999999 0 0.00011289999999999999 3.3 0.00011282 3.3 0.00011292 0 0.00011284 0 0.00011294 3.3 0.00011286 3.3 0.00011296 0 0.00011287999999999999 0 0.00011297999999999999 3.3 0.00011289999999999999 3.3 0.000113 0 0.00011292 0 0.00011302 3.3 0.00011294 3.3 0.00011304 0 0.00011295999999999999 0 0.00011305999999999999 3.3 0.00011297999999999999 3.3 0.00011308 0 0.000113 0 0.0001131 3.3 0.00011302 3.3 0.00011312 0 0.00011304 0 0.00011314 3.3 0.00011305999999999999 3.3 0.00011316 0 0.00011308 0 0.00011318 3.3 0.0001131 3.3 0.0001132 0 0.00011312 0 0.00011322 3.3 0.00011313999999999999 3.3 0.00011324 0 0.00011316 0 0.00011326 3.3 0.00011318 3.3 0.00011328 0 0.0001132 0 0.0001133 3.3 0.00011321999999999999 3.3 0.00011331999999999999 0 0.00011324 0 0.00011334 3.3 0.00011326 3.3 0.00011336 0 0.00011328 0 0.00011338 3.3 0.00011329999999999999 3.3 0.00011339999999999999 0 0.00011331999999999999 0 0.00011342 3.3 0.00011334 3.3 0.00011344 0 0.00011336 0 0.00011346 3.3 0.00011338 3.3 0.00011348 0 0.00011339999999999999 0 0.0001135 3.3 0.00011342 3.3 0.00011352 0 0.00011344 0 0.00011354 3.3 0.00011346 3.3 0.00011356 0 0.00011347999999999999 0 0.00011358 3.3 0.0001135 3.3 0.0001136 0 0.00011352 0 0.00011362 3.3 0.00011354 3.3 0.00011364 0 0.00011355999999999999 0 0.00011365999999999999 3.3 0.00011358 3.3 0.00011368 0 0.0001136 0 0.0001137 3.3 0.00011362 3.3 0.00011372 0 0.00011363999999999999 0 0.00011373999999999999 3.3 0.00011365999999999999 3.3 0.00011376 0 0.00011368 0 0.00011378 3.3 0.0001137 3.3 0.0001138 0 0.00011371999999999999 0 0.00011381999999999999 3.3 0.00011373999999999999 3.3 0.00011384 0 0.00011376 0 0.00011386 3.3 0.00011378 3.3 0.00011388 0 0.0001138 0 0.0001139 3.3 0.00011381999999999999 3.3 0.00011392 0 0.00011384 0 0.00011394 3.3 0.00011386 3.3 0.00011396 0 0.00011388 0 0.00011398 3.3 0.00011389999999999999 3.3 0.00011399999999999999 0 0.00011392 0 0.00011402 3.3 0.00011394 3.3 0.00011404 0 0.00011396 0 0.00011406 3.3 0.00011397999999999999 3.3 0.00011407999999999999 0 0.00011399999999999999 0 0.0001141 3.3 0.00011402 3.3 0.00011412 0 0.00011404 0 0.00011414 3.3 0.00011405999999999999 3.3 0.00011415999999999999 0 0.00011407999999999999 0 0.00011418 3.3 0.0001141 3.3 0.0001142 0 0.00011412 0 0.00011422 3.3 0.00011414 3.3 0.00011424 0 0.00011415999999999999 0 0.00011426 3.3 0.00011418 3.3 0.00011428 0 0.0001142 0 0.0001143 3.3 0.00011422 3.3 0.00011432 0 0.00011423999999999999 0 0.00011433999999999999 3.3 0.00011426 3.3 0.00011436 0 0.00011428 0 0.00011438 3.3 0.0001143 3.3 0.0001144 0 0.00011431999999999999 0 0.00011441999999999999 3.3 0.00011433999999999999 3.3 0.00011444 0 0.00011436 0 0.00011446 3.3 0.00011438 3.3 0.00011448 0 0.00011439999999999999 0 0.00011449999999999999 3.3 0.00011441999999999999 3.3 0.00011452 0 0.00011444 0 0.00011454 3.3 0.00011446 3.3 0.00011456 0 0.00011448 0 0.00011458 3.3 0.00011449999999999999 3.3 0.0001146 0 0.00011452 0 0.00011462 3.3 0.00011454 3.3 0.00011464 0 0.00011456 0 0.00011466 3.3 0.00011457999999999999 3.3 0.00011467999999999999 0 0.0001146 0 0.0001147 3.3 0.00011462 3.3 0.00011472 0 0.00011464 0 0.00011474 3.3 0.00011465999999999999 3.3 0.00011475999999999999 0 0.00011467999999999999 0 0.00011478 3.3 0.0001147 3.3 0.0001148 0 0.00011472 0 0.00011482 3.3 0.00011473999999999999 3.3 0.00011483999999999999 0 0.00011475999999999999 0 0.00011486 3.3 0.00011478 3.3 0.00011488 0 0.0001148 0 0.0001149 3.3 0.00011482 3.3 0.00011492 0 0.00011483999999999999 0 0.00011494 3.3 0.00011486 3.3 0.00011496 0 0.00011488 0 0.00011498 3.3 0.0001149 3.3 0.000115 0 0.00011491999999999999 0 0.00011501999999999999 3.3 0.00011494 3.3 0.00011504 0 0.00011496 0 0.00011506 3.3 0.00011498 3.3 0.00011508 0 0.00011499999999999999 0 0.00011509999999999999 3.3 0.00011501999999999999 3.3 0.00011512 0 0.00011504 0 0.00011514 3.3 0.00011506 3.3 0.00011516 0 0.00011507999999999999 0 0.00011517999999999999 3.3 0.00011509999999999999 3.3 0.0001152 0 0.00011512 0 0.00011522 3.3 0.00011514 3.3 0.00011524 0 0.00011516 0 0.00011526 3.3 0.00011517999999999999 3.3 0.00011528 0 0.0001152 0 0.0001153 3.3 0.00011522 3.3 0.00011532 0 0.00011524 0 0.00011534 3.3 0.00011525999999999999 3.3 0.00011536 0 0.00011528 0 0.00011538 3.3 0.0001153 3.3 0.0001154 0 0.00011532 0 0.00011542 3.3 0.00011533999999999999 3.3 0.00011543999999999999 0 0.00011536 0 0.00011546 3.3 0.00011538 3.3 0.00011548 0 0.0001154 0 0.0001155 3.3 0.00011541999999999999 3.3 0.00011551999999999999 0 0.00011543999999999999 0 0.00011554 3.3 0.00011546 3.3 0.00011556 0 0.00011548 0 0.00011558 3.3 0.00011549999999999999 3.3 0.00011559999999999999 0 0.00011551999999999999 0 0.00011562 3.3 0.00011554 3.3 0.00011564 0 0.00011556 0 0.00011566 3.3 0.00011558 3.3 0.00011568 0 0.00011559999999999999 0 0.0001157 3.3 0.00011562 3.3 0.00011572 0 0.00011564 0 0.00011574 3.3 0.00011566 3.3 0.00011576 0 0.00011567999999999999 0 0.00011577999999999999 3.3 0.0001157 3.3 0.0001158 0 0.00011572 0 0.00011582 3.3 0.00011574 3.3 0.00011584 0 0.00011575999999999999 0 0.00011585999999999999 3.3 0.00011577999999999999 3.3 0.00011588 0 0.0001158 0 0.0001159 3.3 0.00011582 3.3 0.00011592 0 0.00011583999999999999 0 0.00011593999999999999 3.3 0.00011585999999999999 3.3 0.00011596 0 0.00011588 0 0.00011598 3.3 0.0001159 3.3 0.000116 0 0.00011592 0 0.00011602 3.3 0.00011593999999999999 3.3 0.00011604 0 0.00011596 0 0.00011606 3.3 0.00011598 3.3 0.00011608 0 0.000116 0 0.0001161 3.3 0.00011601999999999999 3.3 0.00011611999999999999 0 0.00011604 0 0.00011614 3.3 0.00011606 3.3 0.00011616 0 0.00011608 0 0.00011618 3.3 0.00011609999999999999 3.3 0.00011619999999999999 0 0.00011611999999999999 0 0.00011622 3.3 0.00011614 3.3 0.00011624 0 0.00011616 0 0.00011626 3.3 0.00011617999999999999 3.3 0.00011627999999999999 0 0.00011619999999999999 0 0.0001163 3.3 0.00011622 3.3 0.00011632 0 0.00011624 0 0.00011634 3.3 0.00011626 3.3 0.00011636 0 0.00011627999999999999 0 0.00011638 3.3 0.0001163 3.3 0.0001164 0 0.00011632 0 0.00011642 3.3 0.00011634 3.3 0.00011644 0 0.00011635999999999999 0 0.00011645999999999999 3.3 0.00011638 3.3 0.00011648 0 0.0001164 0 0.0001165 3.3 0.00011642 3.3 0.00011652 0 0.00011643999999999999 0 0.00011653999999999999 3.3 0.00011645999999999999 3.3 0.00011656 0 0.00011648 0 0.00011658 3.3 0.0001165 3.3 0.0001166 0 0.00011651999999999999 0 0.00011661999999999999 3.3 0.00011653999999999999 3.3 0.00011664 0 0.00011656 0 0.00011666 3.3 0.00011658 3.3 0.00011668 0 0.0001166 0 0.0001167 3.3 0.00011661999999999999 3.3 0.00011672 0 0.00011664 0 0.00011674 3.3 0.00011666 3.3 0.00011676 0 0.00011668 0 0.00011678 3.3 0.00011669999999999999 3.3 0.00011679999999999999 0 0.00011672 0 0.00011682 3.3 0.00011674 3.3 0.00011684 0 0.00011676 0 0.00011686 3.3 0.00011677999999999999 3.3 0.00011687999999999999 0 0.00011679999999999999 0 0.0001169 3.3 0.00011682 3.3 0.00011692 0 0.00011684 0 0.00011694 3.3 0.00011685999999999999 3.3 0.00011695999999999999 0 0.00011687999999999999 0 0.00011698 3.3 0.0001169 3.3 0.000117 0 0.00011692 0 0.00011702 3.3 0.00011694 3.3 0.00011704 0 0.00011695999999999999 0 0.00011706 3.3 0.00011698 3.3 0.00011708 0 0.000117 0 0.0001171 3.3 0.00011702 3.3 0.00011712 0 0.00011703999999999999 0 0.00011713999999999999 3.3 0.00011706 3.3 0.00011716 0 0.00011708 0 0.00011718 3.3 0.0001171 3.3 0.0001172 0 0.00011711999999999999 0 0.00011721999999999999 3.3 0.00011713999999999999 3.3 0.00011724 0 0.00011716 0 0.00011726 3.3 0.00011718 3.3 0.00011728 0 0.00011719999999999999 0 0.00011729999999999999 3.3 0.00011721999999999999 3.3 0.00011732 0 0.00011724 0 0.00011734 3.3 0.00011726 3.3 0.00011736 0 0.00011728 0 0.00011738 3.3 0.00011729999999999999 3.3 0.0001174 0 0.00011732 0 0.00011742 3.3 0.00011734 3.3 0.00011744 0 0.00011736 0 0.00011746 3.3 0.00011737999999999999 3.3 0.00011748 0 0.0001174 0 0.0001175 3.3 0.00011742 3.3 0.00011752 0 0.00011744 0 0.00011754 3.3 0.00011745999999999999 3.3 0.00011755999999999999 0 0.00011748 0 0.00011758 3.3 0.0001175 3.3 0.0001176 0 0.00011752 0 0.00011762 3.3 0.00011753999999999999 3.3 0.00011763999999999999 0 0.00011755999999999999 0 0.00011766 3.3 0.00011758 3.3 0.00011768 0 0.0001176 0 0.0001177 3.3 0.00011761999999999999 3.3 0.00011771999999999999 0 0.00011763999999999999 0 0.00011774 3.3 0.00011766 3.3 0.00011776 0 0.00011768 0 0.00011778 3.3 0.0001177 3.3 0.0001178 0 0.00011771999999999999 0 0.00011782 3.3 0.00011774 3.3 0.00011784 0 0.00011776 0 0.00011786 3.3 0.00011778 3.3 0.00011788 0 0.00011779999999999999 0 0.00011789999999999999 3.3 0.00011782 3.3 0.00011792 0 0.00011784 0 0.00011794 3.3 0.00011786 3.3 0.00011796 0 0.00011787999999999999 0 0.00011797999999999999 3.3 0.00011789999999999999 3.3 0.000118 0 0.00011792 0 0.00011802 3.3 0.00011794 3.3 0.00011804 0 0.00011795999999999999 0 0.00011805999999999999 3.3 0.00011797999999999999 3.3 0.00011808 0 0.000118 0 0.0001181 3.3 0.00011802 3.3 0.00011812 0 0.00011804 0 0.00011814 3.3 0.00011805999999999999 3.3 0.00011816 0 0.00011808 0 0.00011818 3.3 0.0001181 3.3 0.0001182 0 0.00011812 0 0.00011822 3.3 0.00011813999999999999 3.3 0.00011823999999999999 0 0.00011816 0 0.00011826 3.3 0.00011818 3.3 0.00011828 0 0.0001182 0 0.0001183 3.3 0.00011821999999999999 3.3 0.00011831999999999999 0 0.00011823999999999999 0 0.00011834 3.3 0.00011826 3.3 0.00011836 0 0.00011828 0 0.00011838 3.3 0.00011829999999999999 3.3 0.00011839999999999999 0 0.00011831999999999999 0 0.00011842 3.3 0.00011834 3.3 0.00011844 0 0.00011836 0 0.00011846 3.3 0.00011838 3.3 0.00011848 0 0.00011839999999999999 0 0.0001185 3.3 0.00011842 3.3 0.00011852 0 0.00011844 0 0.00011854 3.3 0.00011846 3.3 0.00011856 0 0.00011847999999999999 0 0.00011857999999999999 3.3 0.0001185 3.3 0.0001186 0 0.00011852 0 0.00011862 3.3 0.00011854 3.3 0.00011864 0 0.00011855999999999999 0 0.00011865999999999999 3.3 0.00011857999999999999 3.3 0.00011868 0 0.0001186 0 0.0001187 3.3 0.00011862 3.3 0.00011872 0 0.00011863999999999999 0 0.00011873999999999999 3.3 0.00011865999999999999 3.3 0.00011876 0 0.00011868 0 0.00011878 3.3 0.0001187 3.3 0.0001188 0 0.00011872 0 0.00011882 3.3 0.00011873999999999999 3.3 0.00011884 0 0.00011876 0 0.00011886 3.3 0.00011878 3.3 0.00011888 0 0.0001188 0 0.0001189 3.3 0.00011881999999999999 3.3 0.00011891999999999999 0 0.00011884 0 0.00011894 3.3 0.00011886 3.3 0.00011896 0 0.00011888 0 0.00011898 3.3 0.00011889999999999999 3.3 0.00011899999999999999 0 0.00011891999999999999 0 0.00011902 3.3 0.00011894 3.3 0.00011904 0 0.00011896 0 0.00011906 3.3 0.00011897999999999999 3.3 0.00011907999999999999 0 0.00011899999999999999 0 0.0001191 3.3 0.00011902 3.3 0.00011912 0 0.00011904 0 0.00011914 3.3 0.00011906 3.3 0.00011916 0 0.00011907999999999999 0 0.00011918 3.3 0.0001191 3.3 0.0001192 0 0.00011912 0 0.00011922 3.3 0.00011914 3.3 0.00011924 0 0.00011915999999999999 0 0.00011925999999999999 3.3 0.00011918 3.3 0.00011928 0 0.0001192 0 0.0001193 3.3 0.00011922 3.3 0.00011932 0 0.00011923999999999999 0 0.00011933999999999999 3.3 0.00011925999999999999 3.3 0.00011936 0 0.00011928 0 0.00011938 3.3 0.0001193 3.3 0.0001194 0 0.00011931999999999999 0 0.00011941999999999999 3.3 0.00011933999999999999 3.3 0.00011944 0 0.00011936 0 0.00011946 3.3 0.00011938 3.3 0.00011948 0 0.00011939999999999999 0 0.00011949999999999999 3.3 0.00011941999999999999 3.3 0.00011952 0 0.00011944 0 0.00011954 3.3 0.00011946 3.3 0.00011956 0 0.00011948 0 0.00011958 3.3 0.00011949999999999999 3.3 0.0001196 0 0.00011952 0 0.00011962 3.3 0.00011954 3.3 0.00011964 0 0.00011956 0 0.00011966 3.3 0.00011957999999999999 3.3 0.00011967999999999999 0 0.0001196 0 0.0001197 3.3 0.00011962 3.3 0.00011972 0 0.00011964 0 0.00011974 3.3 0.00011965999999999999 3.3 0.00011975999999999999 0 0.00011967999999999999 0 0.00011978 3.3 0.0001197 3.3 0.0001198 0 0.00011972 0 0.00011982 3.3 0.00011973999999999999 3.3 0.00011983999999999999 0 0.00011975999999999999 0 0.00011986 3.3 0.00011978 3.3 0.00011988 0 0.0001198 0 0.0001199 3.3 0.00011982 3.3 0.00011992 0 0.00011983999999999999 0 0.00011994 3.3 0.00011986 3.3 0.00011996 0 0.00011988 0 0.00011998 3.3 0.0001199 3.3 0.00012 0 0.00011991999999999999 0 0.00012001999999999999 3.3 0.00011994 3.3 0.00012004 0 0.00011996 0 0.00012006 3.3 0.00011998 3.3 0.00012008 0 0.00011999999999999999 0 0.00012009999999999999 3.3 0.00012001999999999999 3.3 0.00012012 0 0.00012004 0 0.00012014 3.3 0.00012006 3.3 0.00012016 0 0.00012007999999999999 0 0.00012017999999999999 3.3 0.00012009999999999999 3.3 0.0001202 0 0.00012012 0 0.00012022 3.3 0.00012014 3.3 0.00012024 0 0.00012016 0 0.00012026 3.3 0.00012017999999999999 3.3 0.00012028 0 0.0001202 0 0.0001203 3.3 0.00012022 3.3 0.00012032 0 0.00012024 0 0.00012034 3.3 0.00012025999999999999 3.3 0.00012035999999999999 0 0.00012028 0 0.00012038 3.3 0.0001203 3.3 0.0001204 0 0.00012032 0 0.00012042 3.3 0.00012033999999999999 3.3 0.00012043999999999999 0 0.00012035999999999999 0 0.00012046 3.3 0.00012038 3.3 0.00012048 0 0.0001204 0 0.0001205 3.3 0.00012041999999999999 3.3 0.00012051999999999999 0 0.00012043999999999999 0 0.00012054 3.3 0.00012046 3.3 0.00012056 0 0.00012048 0 0.00012058 3.3 0.0001205 3.3 0.0001206 0 0.00012051999999999999 0 0.00012062 3.3 0.00012054 3.3 0.00012064 0 0.00012056 0 0.00012066 3.3 0.00012058 3.3 0.00012068 0 0.00012059999999999999 0 0.00012069999999999999 3.3 0.00012062 3.3 0.00012072 0 0.00012064 0 0.00012074 3.3 0.00012066 3.3 0.00012076 0 0.00012067999999999999 0 0.00012077999999999999 3.3 0.00012069999999999999 3.3 0.0001208 0 0.00012072 0 0.00012082 3.3 0.00012074 3.3 0.00012084 0 0.00012075999999999999 0 0.00012085999999999999 3.3 0.00012077999999999999 3.3 0.00012088 0 0.0001208 0 0.0001209 3.3 0.00012082 3.3 0.00012092 0 0.00012084 0 0.00012094 3.3 0.00012085999999999999 3.3 0.00012096 0 0.00012088 0 0.00012098 3.3 0.0001209 3.3 0.000121 0 0.00012092 0 0.00012102 3.3 0.00012093999999999999 3.3 0.00012103999999999999 0 0.00012096 0 0.00012106 3.3 0.00012098 3.3 0.00012108 0 0.000121 0 0.0001211 3.3 0.00012101999999999999 3.3 0.00012111999999999999 0 0.00012103999999999999 0 0.00012114 3.3 0.00012106 3.3 0.00012116 0 0.00012108 0 0.00012118 3.3 0.00012109999999999999 3.3 0.00012119999999999999 0 0.00012111999999999999 0 0.00012122 3.3 0.00012114 3.3 0.00012124 0 0.00012116 0 0.00012126 3.3 0.00012117999999999999 3.3 0.00012127999999999999 0 0.00012119999999999999 0 0.0001213 3.3 0.00012122 3.3 0.00012132 0 0.00012124 0 0.00012134 3.3 0.00012126 3.3 0.00012136 0 0.00012127999999999999 0 0.00012137999999999999 3.3 0.0001213 3.3 0.0001214 0 0.00012132 0 0.00012142 3.3 0.00012134 3.3 0.00012144 0 0.00012135999999999999 0 0.00012145999999999999 3.3 0.00012137999999999999 3.3 0.00012148 0 0.0001214 0 0.0001215 3.3 0.00012142 3.3 0.00012152 0 0.00012143999999999999 0 0.00012153999999999999 3.3 0.00012145999999999999 3.3 0.00012156 0 0.00012148 0 0.00012158 3.3 0.0001215 3.3 0.0001216 0 0.00012151999999999999 0 0.00012161999999999999 3.3 0.00012153999999999999 3.3 0.00012164 0 0.00012156 0 0.00012166 3.3 0.00012158 3.3 0.00012168 0 0.0001216 0 0.0001217 3.3 0.00012161999999999999 3.3 0.00012172 0 0.00012164 0 0.00012174 3.3 0.00012166 3.3 0.00012176 0 0.00012168 0 0.00012178 3.3 0.00012169999999999999 3.3 0.00012179999999999999 0 0.00012172 0 0.00012182 3.3 0.00012174 3.3 0.00012184 0 0.00012176 0 0.00012186 3.3 0.00012177999999999999 3.3 0.00012187999999999999 0 0.00012179999999999999 0 0.0001219 3.3 0.00012182 3.3 0.00012192 0 0.00012184 0 0.00012194 3.3 0.00012185999999999999 3.3 0.00012195999999999999 0 0.00012187999999999999 0 0.00012198 3.3 0.0001219 3.3 0.000122 0 0.00012192 0 0.00012202 3.3 0.00012194 3.3 0.00012204 0 0.00012195999999999999 0 0.00012206 3.3 0.00012198 3.3 0.00012208 0 0.00012199999999999998 0 0.00012209999999999999 3.3 0.00012202 3.3 0.00012212 0 0.00012203999999999999 0 0.00012214 3.3 0.00012206000000000001 3.3 0.00012216 0 0.00012208 0 0.00012218 3.3 0.00012209999999999999 3.3 0.0001222 0 0.00012212 0 0.00012222 3.3 0.00012214 3.3 0.00012224 0 0.00012215999999999998 0 0.00012225999999999998 3.3 0.00012218 3.3 0.00012228 0 0.0001222 0 0.0001223 3.3 0.00012222 3.3 0.00012232 0 0.00012224 0 0.00012234 3.3 0.00012225999999999998 3.3 0.00012236 0 0.00012228 0 0.00012238 3.3 0.0001223 3.3 0.0001224 0 0.00012232 0 0.00012242 3.3 0.00012234 3.3 0.00012244 0 0.00012236 0 0.00012246 3.3 0.00012238 3.3 0.00012248 0 0.0001224 0 0.0001225 3.3 0.00012241999999999998 3.3 0.00012251999999999999 0 0.00012244 0 0.00012254 3.3 0.00012246 3.3 0.00012256 0 0.00012248 0 0.00012258 3.3 0.0001225 3.3 0.0001226 0 0.00012251999999999999 0 0.00012262 3.3 0.00012254 3.3 0.00012264 0 0.00012256 0 0.00012266 3.3 0.00012257999999999998 3.3 0.00012267999999999998 0 0.0001226 0 0.0001227 3.3 0.00012262 3.3 0.00012272 0 0.00012264 0 0.00012274 3.3 0.00012266 3.3 0.00012276 0 0.00012267999999999998 0 0.00012278 3.3 0.0001227 3.3 0.0001228 0 0.00012272 0 0.00012282 3.3 0.00012274 3.3 0.00012284 0 0.00012276 0 0.00012286 3.3 0.00012278 3.3 0.00012288 0 0.0001228 0 0.0001229 3.3 0.00012282 3.3 0.00012292 0 0.00012283999999999998 0 0.00012293999999999999 3.3 0.00012286 3.3 0.00012296 0 0.00012288 0 0.00012298 3.3 0.0001229 3.3 0.000123 0 0.00012292 0 0.00012302 3.3 0.00012293999999999999 3.3 0.00012304 0 0.00012296 0 0.00012306 3.3 0.00012298 3.3 0.00012308 0 0.000123 0 0.0001231 3.3 0.00012302 3.3 0.00012312 0 0.00012304 0 0.00012314 3.3 0.00012306 3.3 0.00012316 0 0.00012308 0 0.00012318 3.3 0.00012309999999999998 3.3 0.00012319999999999999 0 0.00012312 0 0.00012322 3.3 0.00012314 3.3 0.00012324 0 0.00012316 0 0.00012326 3.3 0.00012318 3.3 0.00012328 0 0.00012319999999999999 0 0.0001233 3.3 0.00012322 3.3 0.00012332 0 0.00012324 0 0.00012334 3.3 0.00012325999999999998 3.3 0.00012335999999999998 0 0.00012328 0 0.00012338 3.3 0.0001233 3.3 0.0001234 0 0.00012332 0 0.00012342 3.3 0.00012334 3.3 0.00012344 0 0.00012335999999999998 0 0.00012346 3.3 0.00012338 3.3 0.00012348 0 0.0001234 0 0.0001235 3.3 0.00012342 3.3 0.00012352 0 0.00012344 0 0.00012354 3.3 0.00012346 3.3 0.00012356 0 0.00012348 0 0.00012358 3.3 0.0001235 3.3 0.0001236 0 0.00012351999999999998 0 0.00012361999999999999 3.3 0.00012354 3.3 0.00012364 0 0.00012356 0 0.00012366 3.3 0.00012358 3.3 0.00012368 0 0.0001236 0 0.0001237 3.3 0.00012361999999999999 3.3 0.00012372 0 0.00012364 0 0.00012374 3.3 0.00012366 3.3 0.00012376 0 0.00012368 0 0.00012378 3.3 0.0001237 3.3 0.0001238 0 0.00012372 0 0.00012382 3.3 0.00012374 3.3 0.00012384 0 0.00012376 0 0.00012386 3.3 0.00012377999999999998 3.3 0.00012387999999999999 0 0.0001238 0 0.0001239 3.3 0.00012382 3.3 0.00012392 0 0.00012384 0 0.00012394 3.3 0.00012386 3.3 0.00012396 0 0.00012387999999999999 0 0.00012398 3.3 0.0001239 3.3 0.000124 0 0.00012392 0 0.00012402 3.3 0.00012393999999999998 3.3 0.00012403999999999998 0 0.00012396 0 0.00012406 3.3 0.00012398 3.3 0.00012408 0 0.000124 0 0.0001241 3.3 0.00012402 3.3 0.00012412 0 0.00012403999999999998 0 0.00012414 3.3 0.00012406 3.3 0.00012416 0 0.00012408 0 0.00012418 3.3 0.0001241 3.3 0.0001242 0 0.00012412 0 0.00012422 3.3 0.00012414 3.3 0.00012424 0 0.00012416 0 0.00012426 3.3 0.00012418 3.3 0.00012428 0 0.00012419999999999998 0 0.00012429999999999999 3.3 0.00012422 3.3 0.00012432 0 0.00012424 0 0.00012434 3.3 0.00012426 3.3 0.00012436 0 0.00012428 0 0.00012438 3.3 0.00012429999999999999 3.3 0.0001244 0 0.00012432 0 0.00012442 3.3 0.00012434 3.3 0.00012444 0 0.00012435999999999998 0 0.00012445999999999998 3.3 0.00012438 3.3 0.00012448 0 0.0001244 0 0.0001245 3.3 0.00012442 3.3 0.00012452 0 0.00012444 0 0.00012454 3.3 0.00012445999999999998 3.3 0.00012456 0 0.00012448 0 0.00012458 3.3 0.0001245 3.3 0.0001246 0 0.00012452 0 0.00012462 3.3 0.00012454 3.3 0.00012464 0 0.00012456 0 0.00012466 3.3 0.00012458 3.3 0.00012468 0 0.0001246 0 0.0001247 3.3 0.00012461999999999998 3.3 0.00012471999999999998 0 0.00012464 0 0.00012474 3.3 0.00012466 3.3 0.00012476 0 0.00012468 0 0.00012478 3.3 0.0001247 3.3 0.0001248 0 0.00012471999999999998 0 0.00012482 3.3 0.00012474 3.3 0.00012484 0 0.00012476 0 0.00012486 3.3 0.00012478 3.3 0.00012488 0 0.0001248 0 0.0001249 3.3 0.00012482 3.3 0.00012492 0 0.00012484 0 0.00012494 3.3 0.00012486 3.3 0.00012496 0 0.00012487999999999998 0 0.00012497999999999999 3.3 0.0001249 3.3 0.000125 0 0.00012492 0 0.00012502 3.3 0.00012494 3.3 0.00012504 0 0.00012496 0 0.00012506 3.3 0.00012497999999999999 3.3 0.00012508 0 0.000125 0 0.0001251 3.3 0.00012502 3.3 0.00012512 0 0.00012503999999999998 0 0.00012513999999999998 3.3 0.00012506 3.3 0.00012516 0 0.00012508 0 0.00012518 3.3 0.0001251 3.3 0.0001252 0 0.00012512 0 0.00012522 3.3 0.00012513999999999998 3.3 0.00012524 0 0.00012516 0 0.00012526 3.3 0.00012518 3.3 0.00012528 0 0.0001252 0 0.0001253 3.3 0.00012522 3.3 0.00012532 0 0.00012524 0 0.00012534 3.3 0.00012526 3.3 0.00012536 0 0.00012528 0 0.00012538 3.3 0.00012529999999999998 3.3 0.00012539999999999999 0 0.00012532 0 0.00012542 3.3 0.00012534 3.3 0.00012544 0 0.00012536 0 0.00012546 3.3 0.00012538 3.3 0.00012548 0 0.00012539999999999999 0 0.0001255 3.3 0.00012542 3.3 0.00012552 0 0.00012544 0 0.00012554 3.3 0.00012546 3.3 0.00012556 0 0.00012548 0 0.00012558 3.3 0.0001255 3.3 0.0001256 0 0.00012552 0 0.00012562 3.3 0.00012554 3.3 0.00012564 0 0.00012555999999999998 0 0.00012565999999999999 3.3 0.00012558 3.3 0.00012568 0 0.0001256 0 0.0001257 3.3 0.00012562 3.3 0.00012572 0 0.00012564 0 0.00012574 3.3 0.00012565999999999999 3.3 0.00012576 0 0.00012568 0 0.00012578 3.3 0.0001257 3.3 0.0001258 0 0.00012571999999999998 0 0.00012581999999999998 3.3 0.00012574 3.3 0.00012584 0 0.00012576 0 0.00012586 3.3 0.00012578 3.3 0.00012588 0 0.0001258 0 0.0001259 3.3 0.00012581999999999998 3.3 0.00012592 0 0.00012584 0 0.00012594 3.3 0.00012586 3.3 0.00012596 0 0.00012588 0 0.00012598 3.3 0.0001259 3.3 0.000126 0 0.00012592 0 0.00012602 3.3 0.00012594 3.3 0.00012604 0 0.00012596 0 0.00012606 3.3 0.00012597999999999998 3.3 0.00012607999999999999 0 0.000126 0 0.0001261 3.3 0.00012602 3.3 0.00012612 0 0.00012604 0 0.00012614 3.3 0.00012606 3.3 0.00012616 0 0.00012607999999999999 0 0.00012618 3.3 0.0001261 3.3 0.0001262 0 0.00012612 0 0.00012622 3.3 0.00012613999999999998 3.3 0.00012623999999999998 0 0.00012616 0 0.00012626 3.3 0.00012618 3.3 0.00012628 0 0.0001262 0 0.0001263 3.3 0.00012622 3.3 0.00012632 0 0.00012623999999999998 0 0.00012633999999999999 3.3 0.00012626 3.3 0.00012636 0 0.00012628 0 0.00012638 3.3 0.0001263 3.3 0.0001264 0 0.00012632 0 0.00012642 3.3 0.00012633999999999999 3.3 0.00012644 0 0.00012636 0 0.00012646 3.3 0.00012638 3.3 0.00012648 0 0.00012639999999999998 0 0.00012649999999999998 3.3 0.00012642 3.3 0.00012652 0 0.00012644 0 0.00012654 3.3 0.00012646 3.3 0.00012656 0 0.00012648 0 0.00012658 3.3 0.00012649999999999998 3.3 0.0001266 0 0.00012652 0 0.00012662 3.3 0.00012654 3.3 0.00012664 0 0.00012656 0 0.00012666 3.3 0.00012658 3.3 0.00012668 0 0.0001266 0 0.0001267 3.3 0.00012662 3.3 0.00012672 0 0.00012664 0 0.00012674 3.3 0.00012665999999999998 3.3 0.00012675999999999999 0 0.00012668 0 0.00012678 3.3 0.0001267 3.3 0.0001268 0 0.00012672 0 0.00012682 3.3 0.00012674 3.3 0.00012684 0 0.00012675999999999999 0 0.00012686 3.3 0.00012678 3.3 0.00012688 0 0.0001268 0 0.0001269 3.3 0.00012681999999999998 3.3 0.00012691999999999998 0 0.00012684 0 0.00012694 3.3 0.00012686 3.3 0.00012696 0 0.00012688 0 0.00012698 3.3 0.0001269 3.3 0.000127 0 0.00012691999999999998 0 0.00012702 3.3 0.00012694 3.3 0.00012704 0 0.00012696 0 0.00012706 3.3 0.00012698 3.3 0.00012708 0 0.000127 0 0.0001271 3.3 0.00012702 3.3 0.00012712 0 0.00012704 0 0.00012714 3.3 0.00012706 3.3 0.00012716 0 0.00012707999999999998 0 0.00012717999999999999 3.3 0.0001271 3.3 0.0001272 0 0.00012712 0 0.00012722 3.3 0.00012714 3.3 0.00012724 0 0.00012716 0 0.00012726 3.3 0.00012717999999999999 3.3 0.00012728 0 0.0001272 0 0.0001273 3.3 0.00012722 3.3 0.00012732 0 0.00012724 0 0.00012734 3.3 0.00012726 3.3 0.00012736 0 0.00012728 0 0.00012738 3.3 0.0001273 3.3 0.0001274 0 0.00012732 0 0.00012742 3.3 0.00012733999999999998 3.3 0.00012743999999999999 0 0.00012736 0 0.00012746 3.3 0.00012738 3.3 0.00012748 0 0.0001274 0 0.0001275 3.3 0.00012742 3.3 0.00012752 0 0.00012743999999999999 0 0.00012754 3.3 0.00012746 3.3 0.00012756 0 0.00012748 0 0.00012758 3.3 0.00012749999999999998 3.3 0.00012759999999999998 0 0.00012752 0 0.00012762 3.3 0.00012754 3.3 0.00012764 0 0.00012756 0 0.00012766 3.3 0.00012758 3.3 0.00012768 0 0.00012759999999999998 0 0.0001277 3.3 0.00012762 3.3 0.00012772 0 0.00012764 0 0.00012774 3.3 0.00012766 3.3 0.00012776 0 0.00012768 0 0.00012778 3.3 0.0001277 3.3 0.0001278 0 0.00012772 0 0.00012782 3.3 0.00012774 3.3 0.00012784 0 0.00012775999999999998 0 0.00012785999999999999 3.3 0.00012778 3.3 0.00012788 0 0.0001278 0 0.0001279 3.3 0.00012782 3.3 0.00012792 0 0.00012784 0 0.00012794 3.3 0.00012785999999999999 3.3 0.00012796 0 0.00012788 0 0.00012798 3.3 0.0001279 3.3 0.000128 0 0.00012792 0 0.00012802 3.3 0.00012794 3.3 0.00012804 0 0.00012796 0 0.00012806 3.3 0.00012798 3.3 0.00012808 0 0.000128 0 0.0001281 3.3 0.00012801999999999998 3.3 0.00012811999999999999 0 0.00012804 0 0.00012814 3.3 0.00012806 3.3 0.00012816 0 0.00012808 0 0.00012818 3.3 0.0001281 3.3 0.0001282 0 0.00012811999999999999 0 0.00012822 3.3 0.00012814 3.3 0.00012824 0 0.00012816 0 0.00012826 3.3 0.00012817999999999998 3.3 0.00012827999999999998 0 0.0001282 0 0.0001283 3.3 0.00012822 3.3 0.00012832 0 0.00012824 0 0.00012834 3.3 0.00012826 3.3 0.00012836 0 0.00012827999999999998 0 0.00012838 3.3 0.0001283 3.3 0.0001284 0 0.00012832 0 0.00012842 3.3 0.00012834 3.3 0.00012844 0 0.00012836 0 0.00012846 3.3 0.00012838 3.3 0.00012848 0 0.0001284 0 0.0001285 3.3 0.00012842 3.3 0.00012852 0 0.00012843999999999998 0 0.00012853999999999999 3.3 0.00012846 3.3 0.00012856 0 0.00012848 0 0.00012858 3.3 0.0001285 3.3 0.0001286 0 0.00012852 0 0.00012862 3.3 0.00012853999999999999 3.3 0.00012864 0 0.00012856 0 0.00012866 3.3 0.00012858 3.3 0.00012868 0 0.00012859999999999998 0 0.00012869999999999998 3.3 0.00012862 3.3 0.00012872 0 0.00012864 0 0.00012874 3.3 0.00012866 3.3 0.00012876 0 0.00012868 0 0.00012878 3.3 0.00012869999999999998 3.3 0.0001288 0 0.00012872 0 0.00012882 3.3 0.00012874 3.3 0.00012884 0 0.00012876 0 0.00012886 3.3 0.00012878 3.3 0.00012888 0 0.0001288 0 0.0001289 3.3 0.00012882 3.3 0.00012892 0 0.00012884 0 0.00012894 3.3 0.00012885999999999998 3.3 0.00012895999999999999 0 0.00012888 0 0.00012898 3.3 0.0001289 3.3 0.000129 0 0.00012892 0 0.00012902 3.3 0.00012894 3.3 0.00012904 0 0.00012895999999999999 0 0.00012906 3.3 0.00012898 3.3 0.00012908 0 0.000129 0 0.0001291 3.3 0.00012902 3.3 0.00012912 0 0.00012904 0 0.00012914 3.3 0.00012906 3.3 0.00012916 0 0.00012908 0 0.00012918 3.3 0.0001291 3.3 0.0001292 0 0.00012911999999999998 0 0.00012921999999999999 3.3 0.00012914 3.3 0.00012924 0 0.00012916 0 0.00012926 3.3 0.00012918 3.3 0.00012928 0 0.0001292 0 0.0001293 3.3 0.00012921999999999999 3.3 0.00012932 0 0.00012924 0 0.00012934 3.3 0.00012926 3.3 0.00012936 0 0.00012927999999999998 0 0.00012937999999999998 3.3 0.0001293 3.3 0.0001294 0 0.00012932 0 0.00012942 3.3 0.00012934 3.3 0.00012944 0 0.00012936 0 0.00012946 3.3 0.00012937999999999998 3.3 0.00012948 0 0.0001294 0 0.0001295 3.3 0.00012942 3.3 0.00012952 0 0.00012944 0 0.00012954 3.3 0.00012946 3.3 0.00012956 0 0.00012948 0 0.00012958 3.3 0.0001295 3.3 0.0001296 0 0.00012952 0 0.00012962 3.3 0.00012953999999999998 3.3 0.00012963999999999999 0 0.00012956 0 0.00012966 3.3 0.00012958 3.3 0.00012968 0 0.0001296 0 0.0001297 3.3 0.00012962 3.3 0.00012972 0 0.00012963999999999999 0 0.00012974 3.3 0.00012966 3.3 0.00012976 0 0.00012968 0 0.00012978 3.3 0.0001297 3.3 0.0001298 0 0.00012972 0 0.00012982 3.3 0.00012974 3.3 0.00012984 0 0.00012976 0 0.00012986 3.3 0.00012978 3.3 0.00012988 0 0.00012979999999999998 0 0.00012989999999999999 3.3 0.00012982 3.3 0.00012992 0 0.00012984 0 0.00012994 3.3 0.00012986 3.3 0.00012996 0 0.00012988 0 0.00012998 3.3 0.00012989999999999999 3.3 0.00013 0 0.00012992 0 0.00013002 3.3 0.00012994 3.3 0.00013004 0 0.00012995999999999998 0 0.00013005999999999998 3.3 0.00012998 3.3 0.00013008 0 0.00013 0 0.0001301 3.3 0.00013002 3.3 0.00013012 0 0.00013004 0 0.00013014 3.3 0.00013005999999999998 3.3 0.00013016 0 0.00013008 0 0.00013018 3.3 0.0001301 3.3 0.0001302 0 0.00013012 0 0.00013022 3.3 0.00013014 3.3 0.00013024 0 0.00013016 0 0.00013026 3.3 0.00013018 3.3 0.00013028 0 0.0001302 0 0.0001303 3.3 0.00013021999999999998 3.3 0.00013031999999999999 0 0.00013024 0 0.00013034 3.3 0.00013026 3.3 0.00013036 0 0.00013028 0 0.00013038 3.3 0.0001303 3.3 0.0001304 0 0.00013031999999999999 0 0.00013042 3.3 0.00013034 3.3 0.00013044 0 0.00013036 0 0.00013046 3.3 0.00013037999999999998 3.3 0.00013047999999999998 0 0.0001304 0 0.0001305 3.3 0.00013042 3.3 0.00013052 0 0.00013044 0 0.00013054 3.3 0.00013046 3.3 0.00013056 0 0.00013047999999999998 0 0.00013057999999999999 3.3 0.0001305 3.3 0.0001306 0 0.00013052 0 0.00013062 3.3 0.00013054 3.3 0.00013064 0 0.00013056 0 0.00013066 3.3 0.00013057999999999999 3.3 0.00013068 0 0.0001306 0 0.0001307 3.3 0.00013062 3.3 0.00013072 0 0.00013063999999999998 0 0.00013073999999999998 3.3 0.00013066 3.3 0.00013076 0 0.00013068 0 0.00013078 3.3 0.0001307 3.3 0.0001308 0 0.00013072 0 0.00013082 3.3 0.00013073999999999998 3.3 0.00013084 0 0.00013076 0 0.00013086 3.3 0.00013078 3.3 0.00013088 0 0.0001308 0 0.0001309 3.3 0.00013082 3.3 0.00013092 0 0.00013084 0 0.00013094 3.3 0.00013086 3.3 0.00013096 0 0.00013088 0 0.00013098 3.3 0.00013089999999999998 3.3 0.00013099999999999999 0 0.00013092 0 0.00013102 3.3 0.00013094 3.3 0.00013104 0 0.00013096 0 0.00013106 3.3 0.00013098 3.3 0.00013108 0 0.00013099999999999999 0 0.0001311 3.3 0.00013102 3.3 0.00013112 0 0.00013104 0 0.00013114 3.3 0.00013105999999999998 3.3 0.00013115999999999998 0 0.00013108 0 0.00013118 3.3 0.0001311 3.3 0.0001312 0 0.00013112 0 0.00013122 3.3 0.00013114 3.3 0.00013124 0 0.00013115999999999998 0 0.00013126 3.3 0.00013118 3.3 0.00013128 0 0.0001312 0 0.0001313 3.3 0.00013122 3.3 0.00013132 0 0.00013124 0 0.00013134 3.3 0.00013126 3.3 0.00013136 0 0.00013128 0 0.00013138 3.3 0.0001313 3.3 0.0001314 0 0.00013131999999999998 0 0.00013141999999999999 3.3 0.00013134 3.3 0.00013144 0 0.00013136 0 0.00013146 3.3 0.00013138 3.3 0.00013148 0 0.0001314 0 0.0001315 3.3 0.00013141999999999999 3.3 0.00013152 0 0.00013144 0 0.00013154 3.3 0.00013146 3.3 0.00013156 0 0.00013148 0 0.00013158 3.3 0.0001315 3.3 0.0001316 0 0.00013152 0 0.00013162 3.3 0.00013154 3.3 0.00013164 0 0.00013156 0 0.00013166 3.3 0.00013157999999999998 3.3 0.00013167999999999999 0 0.0001316 0 0.0001317 3.3 0.00013162 3.3 0.00013172 0 0.00013164 0 0.00013174 3.3 0.00013166 3.3 0.00013176 0 0.00013167999999999999 0 0.00013178 3.3 0.0001317 3.3 0.0001318 0 0.00013172 0 0.00013182 3.3 0.00013173999999999998 3.3 0.00013183999999999998 0 0.00013176 0 0.00013186 3.3 0.00013178 3.3 0.00013188 0 0.0001318 0 0.0001319 3.3 0.00013182 3.3 0.00013192 0 0.00013183999999999998 0 0.00013194 3.3 0.00013186 3.3 0.00013196 0 0.00013188 0 0.00013198 3.3 0.0001319 3.3 0.000132 0 0.00013192 0 0.00013202 3.3 0.00013194 3.3 0.00013204 0 0.00013196 0 0.00013206 3.3 0.00013198 3.3 0.00013208 0 0.00013199999999999998 0 0.00013209999999999999 3.3 0.00013202 3.3 0.00013212 0 0.00013204 0 0.00013214 3.3 0.00013206 3.3 0.00013216 0 0.00013208 0 0.00013218 3.3 0.00013209999999999999 3.3 0.0001322 0 0.00013212 0 0.00013222 3.3 0.00013214 3.3 0.00013224 0 0.00013215999999999998 0 0.00013225999999999998 3.3 0.00013218 3.3 0.00013228 0 0.0001322 0 0.0001323 3.3 0.00013222 3.3 0.00013232 0 0.00013224 0 0.00013234 3.3 0.00013225999999999998 3.3 0.00013235999999999999 0 0.00013228 0 0.00013238 3.3 0.0001323 3.3 0.0001324 0 0.00013232 0 0.00013242 3.3 0.00013234 3.3 0.00013244 0 0.00013235999999999999 0 0.00013246 3.3 0.00013238 3.3 0.00013248 0 0.0001324 0 0.0001325 3.3 0.00013241999999999998 3.3 0.00013251999999999998 0 0.00013244 0 0.00013254 3.3 0.00013246 3.3 0.00013256 0 0.00013248 0 0.00013258 3.3 0.0001325 3.3 0.0001326 0 0.00013251999999999998 0 0.00013262 3.3 0.00013254 3.3 0.00013264 0 0.00013256 0 0.00013266 3.3 0.00013258 3.3 0.00013268 0 0.0001326 0 0.0001327 3.3 0.00013262 3.3 0.00013272 0 0.00013264 0 0.00013274 3.3 0.00013266 3.3 0.00013276 0 0.00013267999999999998 0 0.00013277999999999999 3.3 0.0001327 3.3 0.0001328 0 0.00013272 0 0.00013282 3.3 0.00013274 3.3 0.00013284 0 0.00013276 0 0.00013286 3.3 0.00013277999999999999 3.3 0.00013288 0 0.0001328 0 0.0001329 3.3 0.00013282 3.3 0.00013292 0 0.00013283999999999998 0 0.00013293999999999998 3.3 0.00013286 3.3 0.00013296 0 0.00013288 0 0.00013298 3.3 0.0001329 3.3 0.000133 0 0.00013292 0 0.00013302 3.3 0.00013293999999999998 3.3 0.00013304 0 0.00013296 0 0.00013306 3.3 0.00013298 3.3 0.00013308 0 0.000133 0 0.0001331 3.3 0.00013302 3.3 0.00013312 0 0.00013304 0 0.00013314 3.3 0.00013306 3.3 0.00013316 0 0.00013308 0 0.00013318 3.3 0.00013309999999999998 3.3 0.00013319999999999999 0 0.00013312 0 0.00013322 3.3 0.00013314 3.3 0.00013324 0 0.00013316 0 0.00013326 3.3 0.00013318 3.3 0.00013328 0 0.00013319999999999999 0 0.0001333 3.3 0.00013322 3.3 0.00013332 0 0.00013324 0 0.00013334 3.3 0.00013326 3.3 0.00013336 0 0.00013328 0 0.00013338 3.3 0.0001333 3.3 0.0001334 0 0.00013332 0 0.00013342 3.3 0.00013334 3.3 0.00013344 0 0.00013335999999999998 0 0.00013345999999999999 3.3 0.00013338 3.3 0.00013348 0 0.0001334 0 0.0001335 3.3 0.00013342 3.3 0.00013352 0 0.00013344 0 0.00013354 3.3 0.00013345999999999999 3.3 0.00013356 0 0.00013348 0 0.00013358 3.3 0.0001335 3.3 0.0001336 0 0.00013351999999999998 0 0.00013361999999999998 3.3 0.00013354 3.3 0.00013364 0 0.00013356 0 0.00013366 3.3 0.00013358 3.3 0.00013368 0 0.0001336 0 0.0001337 3.3 0.00013361999999999998 3.3 0.00013372 0 0.00013364 0 0.00013374 3.3 0.00013366 3.3 0.00013376 0 0.00013368 0 0.00013378 3.3 0.0001337 3.3 0.0001338 0 0.00013372 0 0.00013382 3.3 0.00013374 3.3 0.00013384 0 0.00013376 0 0.00013386 3.3 0.00013377999999999998 3.3 0.00013387999999999999 0 0.0001338 0 0.0001339 3.3 0.00013382 3.3 0.00013392 0 0.00013384 0 0.00013394 3.3 0.00013386 3.3 0.00013396 0 0.00013387999999999999 0 0.00013398 3.3 0.0001339 3.3 0.000134 0 0.00013392 0 0.00013402 3.3 0.00013393999999999998 3.3 0.00013403999999999998 0 0.00013396 0 0.00013406 3.3 0.00013398 3.3 0.00013408 0 0.000134 0 0.0001341 3.3 0.00013402 3.3 0.00013412 0 0.00013403999999999998 0 0.00013413999999999999 3.3 0.00013406 3.3 0.00013416 0 0.00013408 0 0.00013418 3.3 0.0001341 3.3 0.0001342 0 0.00013412 0 0.00013422 3.3 0.00013413999999999999 3.3 0.00013424 0 0.00013416 0 0.00013426 3.3 0.00013418 3.3 0.00013428 0 0.00013419999999999998 0 0.00013429999999999998 3.3 0.00013422 3.3 0.00013432 0 0.00013424 0 0.00013434 3.3 0.00013426 3.3 0.00013436 0 0.00013428 0 0.00013438 3.3 0.00013429999999999998 3.3 0.0001344 0 0.00013432 0 0.00013442 3.3 0.00013434 3.3 0.00013444 0 0.00013436 0 0.00013446 3.3 0.00013438 3.3 0.00013448 0 0.0001344 0 0.0001345 3.3 0.00013442 3.3 0.00013452 0 0.00013444 0 0.00013454 3.3 0.00013445999999999998 3.3 0.00013455999999999999 0 0.00013448 0 0.00013458 3.3 0.0001345 3.3 0.0001346 0 0.00013452 0 0.00013462 3.3 0.00013454 3.3 0.00013464 0 0.00013455999999999999 0 0.00013466 3.3 0.00013458 3.3 0.00013468 0 0.0001346 0 0.0001347 3.3 0.00013461999999999998 3.3 0.00013471999999999998 0 0.00013464 0 0.00013474 3.3 0.00013466 3.3 0.00013476 0 0.00013468 0 0.00013478 3.3 0.0001347 3.3 0.0001348 0 0.00013471999999999998 0 0.00013482 3.3 0.00013474 3.3 0.00013484 0 0.00013476 0 0.00013486 3.3 0.00013478 3.3 0.00013488 0 0.0001348 0 0.0001349 3.3 0.00013482 3.3 0.00013492 0 0.00013484 0 0.00013494 3.3 0.00013486 3.3 0.00013496 0 0.00013487999999999998 0 0.00013497999999999998 3.3 0.0001349 3.3 0.000135 0 0.00013492 0 0.00013502 3.3 0.00013494 3.3 0.00013504 0 0.00013496 0 0.00013506 3.3 0.00013497999999999998 3.3 0.00013508 0 0.000135 0 0.0001351 3.3 0.00013502 3.3 0.00013512 0 0.00013504 0 0.00013514 3.3 0.00013506 3.3 0.00013516 0 0.00013508 0 0.00013518 3.3 0.0001351 3.3 0.0001352 0 0.00013512 0 0.00013522 3.3 0.00013513999999999998 3.3 0.00013523999999999999 0 0.00013516 0 0.00013526 3.3 0.00013518 3.3 0.00013528 0 0.0001352 0 0.0001353 3.3 0.00013522 3.3 0.00013532 0 0.00013523999999999999 0 0.00013534 3.3 0.00013526 3.3 0.00013536 0 0.00013528 0 0.00013538 3.3 0.00013529999999999998 3.3 0.00013539999999999998 0 0.00013532 0 0.00013542 3.3 0.00013534 3.3 0.00013544 0 0.00013536 0 0.00013546 3.3 0.00013538 3.3 0.00013548 0 0.00013539999999999998 0 0.0001355 3.3 0.00013542 3.3 0.00013552 0 0.00013544 0 0.00013554 3.3 0.00013546 3.3 0.00013556 0 0.00013548 0 0.00013558 3.3 0.0001355 3.3 0.0001356 0 0.00013552 0 0.00013562 3.3 0.00013554 3.3 0.00013564 0 0.00013555999999999998 0 0.00013565999999999999 3.3 0.00013558 3.3 0.00013568 0 0.0001356 0 0.0001357 3.3 0.00013562 3.3 0.00013572 0 0.00013564 0 0.00013574 3.3 0.00013565999999999999 3.3 0.00013576 0 0.00013568 0 0.00013578 3.3 0.0001357 3.3 0.0001358 0 0.00013572 0 0.00013582 3.3 0.00013574 3.3 0.00013584 0 0.00013576 0 0.00013586 3.3 0.00013578 3.3 0.00013588 0 0.0001358 0 0.0001359 3.3 0.00013581999999999998 3.3 0.00013591999999999999 0 0.00013584 0 0.00013594 3.3 0.00013586 3.3 0.00013596 0 0.00013588 0 0.00013598 3.3 0.0001359 3.3 0.000136 0 0.00013591999999999999 0 0.00013602 3.3 0.00013594 3.3 0.00013604 0 0.00013596 0 0.00013606 3.3 0.00013597999999999998 3.3 0.00013607999999999998 0 0.000136 0 0.0001361 3.3 0.00013602 3.3 0.00013612 0 0.00013604 0 0.00013614 3.3 0.00013606 3.3 0.00013616 0 0.00013607999999999998 0 0.00013618 3.3 0.0001361 3.3 0.0001362 0 0.00013612 0 0.00013622 3.3 0.00013614 3.3 0.00013624 0 0.00013616 0 0.00013626 3.3 0.00013618 3.3 0.00013628 0 0.0001362 0 0.0001363 3.3 0.00013622 3.3 0.00013632 0 0.00013623999999999998 0 0.00013633999999999999 3.3 0.00013626 3.3 0.00013636 0 0.00013628 0 0.00013638 3.3 0.0001363 3.3 0.0001364 0 0.00013632 0 0.00013642 3.3 0.00013633999999999999 3.3 0.00013644 0 0.00013636 0 0.00013646 3.3 0.00013638 3.3 0.00013648 0 0.00013639999999999998 0 0.00013649999999999998 3.3 0.00013642 3.3 0.00013652 0 0.00013644 0 0.00013654 3.3 0.00013646 3.3 0.00013656 0 0.00013648 0 0.00013658 3.3 0.00013649999999999998 3.3 0.00013659999999999999 0 0.00013652 0 0.00013662 3.3 0.00013654 3.3 0.00013664 0 0.00013656 0 0.00013666 3.3 0.00013658 3.3 0.00013668 0 0.00013659999999999999 0 0.0001367 3.3 0.00013662 3.3 0.00013672 0 0.00013664 0 0.00013674 3.3 0.00013665999999999998 3.3 0.00013675999999999998 0 0.00013668 0 0.00013678 3.3 0.0001367 3.3 0.0001368 0 0.00013672 0 0.00013682 3.3 0.00013674 3.3 0.00013684 0 0.00013675999999999998 0 0.00013686 3.3 0.00013678 3.3 0.00013688 0 0.0001368 0 0.0001369 3.3 0.00013682 3.3 0.00013692 0 0.00013684 0 0.00013694 3.3 0.00013686 3.3 0.00013696 0 0.00013688 0 0.00013698 3.3 0.0001369 3.3 0.000137 0 0.00013691999999999998 0 0.00013701999999999999 3.3 0.00013694 3.3 0.00013704 0 0.00013696 0 0.00013706 3.3 0.00013698 3.3 0.00013708 0 0.000137 0 0.0001371 3.3 0.00013701999999999999 3.3 0.00013712 0 0.00013704 0 0.00013714 3.3 0.00013706 3.3 0.00013716 0 0.00013707999999999998 0 0.00013717999999999998 3.3 0.0001371 3.3 0.0001372 0 0.00013712 0 0.00013722 3.3 0.00013714 3.3 0.00013724 0 0.00013716 0 0.00013726 3.3 0.00013717999999999998 3.3 0.00013728 0 0.0001372 0 0.0001373 3.3 0.00013722 3.3 0.00013732 0 0.00013724 0 0.00013734 3.3 0.00013726 3.3 0.00013736 0 0.00013728 0 0.00013738 3.3 0.0001373 3.3 0.0001374 0 0.00013732 0 0.00013742 3.3 0.00013733999999999998 3.3 0.00013743999999999999 0 0.00013736 0 0.00013746 3.3 0.00013738 3.3 0.00013748 0 0.0001374 0 0.0001375 3.3 0.00013742 3.3 0.00013752 0 0.00013743999999999999 0 0.00013754 3.3 0.00013746 3.3 0.00013756 0 0.00013748 0 0.00013758 3.3 0.0001375 3.3 0.0001376 0 0.00013752 0 0.00013762 3.3 0.00013754 3.3 0.00013764 0 0.00013756 0 0.00013766 3.3 0.00013758 3.3 0.00013768 0 0.00013759999999999998 0 0.00013769999999999999 3.3 0.00013762 3.3 0.00013772 0 0.00013764 0 0.00013774 3.3 0.00013766 3.3 0.00013776 0 0.00013768 0 0.00013778 3.3 0.00013769999999999999 3.3 0.0001378 0 0.00013772 0 0.00013782 3.3 0.00013774 3.3 0.00013784 0 0.00013775999999999998 0 0.00013785999999999998 3.3 0.00013778 3.3 0.00013788 0 0.0001378 0 0.0001379 3.3 0.00013782 3.3 0.00013792 0 0.00013784 0 0.00013794 3.3 0.00013785999999999998 3.3 0.00013796 0 0.00013788 0 0.00013798 3.3 0.0001379 3.3 0.000138 0 0.00013792 0 0.00013802 3.3 0.00013794 3.3 0.00013804 0 0.00013796 0 0.00013806 3.3 0.00013798 3.3 0.00013808 0 0.000138 0 0.0001381 3.3 0.00013801999999999998 3.3 0.00013811999999999999 0 0.00013804 0 0.00013814 3.3 0.00013806 3.3 0.00013816 0 0.00013808 0 0.00013818 3.3 0.0001381 3.3 0.0001382 0 0.00013811999999999999 0 0.00013822 3.3 0.00013814 3.3 0.00013824 0 0.00013816 0 0.00013826 3.3 0.00013817999999999998 3.3 0.00013827999999999998 0 0.0001382 0 0.0001383 3.3 0.00013822 3.3 0.00013832 0 0.00013824 0 0.00013834 3.3 0.00013826 3.3 0.00013836 0 0.00013827999999999998 0 0.00013837999999999999 3.3 0.0001383 3.3 0.0001384 0 0.00013832 0 0.00013842 3.3 0.00013834 3.3 0.00013844 0 0.00013836 0 0.00013846 3.3 0.00013837999999999999 3.3 0.00013848 0 0.0001384 0 0.0001385 3.3 0.00013842 3.3 0.00013852 0 0.00013843999999999998 0 0.00013853999999999998 3.3 0.00013846 3.3 0.00013856 0 0.00013848 0 0.00013858 3.3 0.0001385 3.3 0.0001386 0 0.00013852 0 0.00013862 3.3 0.00013853999999999998 3.3 0.00013864 0 0.00013856 0 0.00013866 3.3 0.00013858 3.3 0.00013868 0 0.0001386 0 0.0001387 3.3 0.00013862 3.3 0.00013872 0 0.00013864 0 0.00013874 3.3 0.00013866 3.3 0.00013876 0 0.00013868 0 0.00013878 3.3 0.00013869999999999998 3.3 0.00013879999999999999 0 0.00013872 0 0.00013882 3.3 0.00013874 3.3 0.00013884 0 0.00013876 0 0.00013886 3.3 0.00013878 3.3 0.00013888 0 0.00013879999999999999 0 0.0001389 3.3 0.00013882 3.3 0.00013892 0 0.00013884 0 0.00013894 3.3 0.00013885999999999998 3.3 0.00013895999999999998 0 0.00013888 0 0.00013898 3.3 0.0001389 3.3 0.000139 0 0.00013892 0 0.00013902 3.3 0.00013894 3.3 0.00013904 0 0.00013895999999999998 0 0.00013906 3.3 0.00013898 3.3 0.00013908 0 0.000139 0 0.0001391 3.3 0.00013902 3.3 0.00013912 0 0.00013904 0 0.00013914 3.3 0.00013906 3.3 0.00013916 0 0.00013908 0 0.00013918 3.3 0.0001391 3.3 0.0001392 0 0.00013911999999999998 0 0.00013921999999999999 3.3 0.00013914 3.3 0.00013924 0 0.00013916 0 0.00013926 3.3 0.00013918 3.3 0.00013928 0 0.0001392 0 0.0001393 3.3 0.00013921999999999999 3.3 0.00013932 0 0.00013924 0 0.00013934 3.3 0.00013926 3.3 0.00013936 0 0.00013928 0 0.00013938 3.3 0.0001393 3.3 0.0001394 0 0.00013932 0 0.00013942 3.3 0.00013934 3.3 0.00013944 0 0.00013936 0 0.00013946 3.3 0.00013937999999999998 3.3 0.00013947999999999999 0 0.0001394 0 0.0001395 3.3 0.00013942 3.3 0.00013952 0 0.00013944 0 0.00013954 3.3 0.00013946 3.3 0.00013956 0 0.00013947999999999999 0 0.00013958 3.3 0.0001395 3.3 0.0001396 0 0.00013952 0 0.00013962 3.3 0.00013953999999999998 3.3 0.00013963999999999998 0 0.00013956 0 0.00013966 3.3 0.00013958 3.3 0.00013968 0 0.0001396 0 0.0001397 3.3 0.00013962 3.3 0.00013972 0 0.00013963999999999998 0 0.00013974 3.3 0.00013966 3.3 0.00013976 0 0.00013968 0 0.00013978 3.3 0.0001397 3.3 0.0001398 0 0.00013972 0 0.00013982 3.3 0.00013974 3.3 0.00013984 0 0.00013976 0 0.00013986 3.3 0.00013978 3.3 0.00013988 0 0.00013979999999999998 0 0.00013989999999999999 3.3 0.00013982 3.3 0.00013992 0 0.00013984 0 0.00013994 3.3 0.00013986 3.3 0.00013996 0 0.00013988 0 0.00013998 3.3 0.00013989999999999999 3.3 0.00014 0 0.00013992 0 0.00014002 3.3 0.00013994 3.3 0.00014004 0 0.00013995999999999998 0 0.00014005999999999998 3.3 0.00013998 3.3 0.00014008 0 0.00014 0 0.0001401 3.3 0.00014002 3.3 0.00014012 0 0.00014004 0 0.00014014 3.3 0.00014005999999999998 3.3 0.00014015999999999999 0 0.00014008 0 0.00014018 3.3 0.0001401 3.3 0.0001402 0 0.00014012 0 0.00014022 3.3 0.00014014 3.3 0.00014024 0 0.00014015999999999999 0 0.00014026 3.3 0.00014018 3.3 0.00014028 0 0.0001402 0 0.0001403 3.3 0.00014021999999999998 3.3 0.00014031999999999998 0 0.00014024 0 0.00014034 3.3 0.00014026 3.3 0.00014036 0 0.00014028 0 0.00014038 3.3 0.0001403 3.3 0.0001404 0 0.00014031999999999998 0 0.00014042 3.3 0.00014034 3.3 0.00014044 0 0.00014036 0 0.00014046 3.3 0.00014038 3.3 0.00014048 0 0.0001404 0 0.0001405 3.3 0.00014042 3.3 0.00014052 0 0.00014044 0 0.00014054 3.3 0.00014046 3.3 0.00014056 0 0.00014047999999999998 0 0.00014057999999999999 3.3 0.0001405 3.3 0.0001406 0 0.00014052 0 0.00014062 3.3 0.00014054 3.3 0.00014064 0 0.00014056 0 0.00014066 3.3 0.00014057999999999999 3.3 0.00014068 0 0.0001406 0 0.0001407 3.3 0.00014062 3.3 0.00014072 0 0.00014063999999999998 0 0.00014073999999999998 3.3 0.00014066 3.3 0.00014076 0 0.00014068 0 0.00014078 3.3 0.0001407 3.3 0.0001408 0 0.00014072 0 0.00014082 3.3 0.00014073999999999998 3.3 0.00014084 0 0.00014076 0 0.00014086 3.3 0.00014078 3.3 0.00014088 0 0.0001408 0 0.0001409 3.3 0.00014082 3.3 0.00014092 0 0.00014084 0 0.00014094 3.3 0.00014086 3.3 0.00014096 0 0.00014088 0 0.00014098 3.3 0.00014089999999999998 3.3 0.00014099999999999998 0 0.00014092 0 0.00014102 3.3 0.00014094 3.3 0.00014104 0 0.00014096 0 0.00014106 3.3 0.00014098 3.3 0.00014108 0 0.00014099999999999998 0 0.0001411 3.3 0.00014102 3.3 0.00014112 0 0.00014104 0 0.00014114 3.3 0.00014106 3.3 0.00014116 0 0.00014108 0 0.00014118 3.3 0.0001411 3.3 0.0001412 0 0.00014112 0 0.00014122 3.3 0.00014114 3.3 0.00014124 0 0.00014115999999999998 0 0.00014125999999999999 3.3 0.00014118 3.3 0.00014128 0 0.0001412 0 0.0001413 3.3 0.00014122 3.3 0.00014132 0 0.00014124 0 0.00014134 3.3 0.00014125999999999999 3.3 0.00014136 0 0.00014128 0 0.00014138 3.3 0.0001413 3.3 0.0001414 0 0.00014131999999999998 0 0.00014141999999999998 3.3 0.00014134 3.3 0.00014144 0 0.00014136 0 0.00014146 3.3 0.00014138 3.3 0.00014148 0 0.0001414 0 0.0001415 3.3 0.00014141999999999998 3.3 0.00014152 0 0.00014144 0 0.00014154 3.3 0.00014146 3.3 0.00014156 0 0.00014148 0 0.00014158 3.3 0.0001415 3.3 0.0001416 0 0.00014152 0 0.00014162 3.3 0.00014154 3.3 0.00014164 0 0.00014156 0 0.00014166 3.3 0.00014157999999999998 3.3 0.00014167999999999999 0 0.0001416 0 0.0001417 3.3 0.00014162 3.3 0.00014172 0 0.00014164 0 0.00014174 3.3 0.00014166 3.3 0.00014176 0 0.00014167999999999999 0 0.00014178 3.3 0.0001417 3.3 0.0001418 0 0.00014172 0 0.00014182 3.3 0.00014173999999999998 3.3 0.00014183999999999998 0 0.00014176 0 0.00014186 3.3 0.00014178 3.3 0.00014188 0 0.0001418 0 0.0001419 3.3 0.00014182 3.3 0.00014192 0 0.00014183999999999998 0 0.00014193999999999999 3.3 0.00014186 3.3 0.00014196 0 0.00014188 0 0.00014198 3.3 0.0001419 3.3 0.000142 0 0.00014192 0 0.00014202 3.3 0.00014193999999999999 3.3 0.00014204 0 0.00014196 0 0.00014206 3.3 0.00014198 3.3 0.00014208 0 0.00014199999999999998 0 0.00014209999999999998 3.3 0.00014202 3.3 0.00014212 0 0.00014204 0 0.00014214 3.3 0.00014206 3.3 0.00014216 0 0.00014208 0 0.00014218 3.3 0.00014209999999999998 3.3 0.0001422 0 0.00014212 0 0.00014222 3.3 0.00014214 3.3 0.00014224 0 0.00014216 0 0.00014226 3.3 0.00014218 3.3 0.00014228 0 0.0001422 0 0.0001423 3.3 0.00014222 3.3 0.00014232 0 0.00014224 0 0.00014234 3.3 0.00014225999999999998 3.3 0.00014235999999999999 0 0.00014228 0 0.00014238 3.3 0.0001423 3.3 0.0001424 0 0.00014232 0 0.00014242 3.3 0.00014234 3.3 0.00014244 0 0.00014235999999999999 0 0.00014246 3.3 0.00014238 3.3 0.00014248 0 0.0001424 0 0.0001425 3.3 0.00014241999999999998 3.3 0.00014251999999999998 0 0.00014244 0 0.00014254 3.3 0.00014246 3.3 0.00014256 0 0.00014248 0 0.00014258 3.3 0.0001425 3.3 0.0001426 0 0.00014251999999999998 0 0.00014261999999999999 3.3 0.00014254 3.3 0.00014264 0 0.00014256 0 0.00014266 3.3 0.00014258 3.3 0.00014268 0 0.0001426 0 0.0001427 3.3 0.00014261999999999999 3.3 0.00014272 0 0.00014264 0 0.00014274 3.3 0.00014266 3.3 0.00014276 0 0.00014267999999999998 0 0.00014277999999999998 3.3 0.0001427 3.3 0.0001428 0 0.00014272 0 0.00014282 3.3 0.00014274 3.3 0.00014284 0 0.00014276 0 0.00014286 3.3 0.00014277999999999998 3.3 0.00014288 0 0.0001428 0 0.0001429 3.3 0.00014282 3.3 0.00014292 0 0.00014284 0 0.00014294 3.3 0.00014286 3.3 0.00014296 0 0.00014288 0 0.00014298 3.3 0.0001429 3.3 0.000143 0 0.00014292 0 0.00014302 3.3 0.00014293999999999998 3.3 0.00014303999999999999 0 0.00014296 0 0.00014306 3.3 0.00014298 3.3 0.00014308 0 0.000143 0 0.0001431 3.3 0.00014302 3.3 0.00014312 0 0.00014303999999999999 0 0.00014314 3.3 0.00014306 3.3 0.00014316 0 0.00014308 0 0.00014318 3.3 0.00014309999999999998 3.3 0.00014319999999999998 0 0.00014312 0 0.00014322 3.3 0.00014314 3.3 0.00014324 0 0.00014316 0 0.00014326 3.3 0.00014318 3.3 0.00014328 0 0.00014319999999999998 0 0.0001433 3.3 0.00014322 3.3 0.00014332 0 0.00014324 0 0.00014334 3.3 0.00014326 3.3 0.00014336 0 0.00014328 0 0.00014338 3.3 0.0001433 3.3 0.0001434 0 0.00014332 0 0.00014342 3.3 0.00014334 3.3 0.00014344 0 0.00014335999999999998 0 0.00014345999999999999 3.3 0.00014338 3.3 0.00014348 0 0.0001434 0 0.0001435 3.3 0.00014342 3.3 0.00014352 0 0.00014344 0 0.00014354 3.3 0.00014345999999999999 3.3 0.00014356 0 0.00014348 0 0.00014358 3.3 0.0001435 3.3 0.0001436 0 0.00014351999999999998 0 0.00014361999999999998 3.3 0.00014354 3.3 0.00014364 0 0.00014356 0 0.00014366 3.3 0.00014358 3.3 0.00014368 0 0.0001436 0 0.0001437 3.3 0.00014361999999999998 3.3 0.00014371999999999999 0 0.00014364 0 0.00014374 3.3 0.00014366 3.3 0.00014376 0 0.00014368 0 0.00014378 3.3 0.0001437 3.3 0.0001438 0 0.00014371999999999999 0 0.00014382 3.3 0.00014374 3.3 0.00014384 0 0.00014376 0 0.00014386 3.3 0.00014377999999999998 3.3 0.00014387999999999998 0 0.0001438 0 0.0001439 3.3 0.00014382 3.3 0.00014392 0 0.00014384 0 0.00014394 3.3 0.00014386 3.3 0.00014396 0 0.00014387999999999998 0 0.00014398 3.3 0.0001439 3.3 0.000144 0 0.00014392 0 0.00014402 3.3 0.00014394 3.3 0.00014404 0 0.00014396 0 0.00014406 3.3 0.00014398 3.3 0.00014408 0 0.000144 0 0.0001441 3.3 0.00014402 3.3 0.00014412 0 0.00014403999999999998 0 0.00014413999999999999 3.3 0.00014406 3.3 0.00014416 0 0.00014408 0 0.00014418 3.3 0.0001441 3.3 0.0001442 0 0.00014412 0 0.00014422 3.3 0.00014413999999999999 3.3 0.00014424 0 0.00014416 0 0.00014426 3.3 0.00014418 3.3 0.00014428 0 0.00014419999999999998 0 0.00014429999999999998 3.3 0.00014422 3.3 0.00014432 0 0.00014424 0 0.00014434 3.3 0.00014426 3.3 0.00014436 0 0.00014428 0 0.00014438 3.3 0.00014429999999999998 3.3 0.00014439999999999999 0 0.00014432 0 0.00014442 3.3 0.00014434 3.3 0.00014444 0 0.00014436 0 0.00014446 3.3 0.00014438 3.3 0.00014448 0 0.00014439999999999999 0 0.0001445 3.3 0.00014442 3.3 0.00014452 0 0.00014444 0 0.00014454 3.3 0.00014445999999999998 3.3 0.00014455999999999998 0 0.00014448 0 0.00014458 3.3 0.0001445 3.3 0.0001446 0 0.00014452 0 0.00014462 3.3 0.00014454 3.3 0.00014464 0 0.00014455999999999998 0 0.00014466 3.3 0.00014458 3.3 0.00014468 0 0.0001446 0 0.0001447 3.3 0.00014462 3.3 0.00014472 0 0.00014464 0 0.00014474 3.3 0.00014466 3.3 0.00014476 0 0.00014468 0 0.00014478 3.3 0.0001447 3.3 0.0001448 0 0.00014471999999999998 0 0.00014481999999999999 3.3 0.00014474 3.3 0.00014484 0 0.00014476 0 0.00014486 3.3 0.00014478 3.3 0.00014488 0 0.0001448 0 0.0001449 3.3 0.00014481999999999999 3.3 0.00014492 0 0.00014484 0 0.00014494 3.3 0.00014486 3.3 0.00014496 0 0.00014487999999999998 0 0.00014497999999999998 3.3 0.0001449 3.3 0.000145 0 0.00014492 0 0.00014502 3.3 0.00014494 3.3 0.00014504 0 0.00014496 0 0.00014506 3.3 0.00014497999999999998 3.3 0.00014508 0 0.000145 0 0.0001451 3.3 0.00014502 3.3 0.00014512 0 0.00014504 0 0.00014514 3.3 0.00014506 3.3 0.00014516 0 0.00014508 0 0.00014518 3.3 0.0001451 3.3 0.0001452 0 0.00014512 0 0.00014522 3.3 0.00014513999999999998 3.3 0.00014523999999999998 0 0.00014516 0 0.00014526 3.3 0.00014518 3.3 0.00014528 0 0.0001452 0 0.0001453 3.3 0.00014522 3.3 0.00014532 0 0.00014523999999999998 0 0.00014534 3.3 0.00014526 3.3 0.00014536 0 0.00014528 0 0.00014538 3.3 0.0001453 3.3 0.0001454 0 0.00014532 0 0.00014542 3.3 0.00014534 3.3 0.00014544 0 0.00014536 0 0.00014546 3.3 0.00014538 3.3 0.00014548 0 0.00014539999999999998 0 0.00014549999999999999 3.3 0.00014542 3.3 0.00014552 0 0.00014544 0 0.00014554 3.3 0.00014546 3.3 0.00014556 0 0.00014548 0 0.00014558 3.3 0.00014549999999999999 3.3 0.0001456 0 0.00014552 0 0.00014562 3.3 0.00014554 3.3 0.00014564 0 0.00014555999999999998 0 0.00014565999999999998 3.3 0.00014558 3.3 0.00014568 0 0.0001456 0 0.0001457 3.3 0.00014562 3.3 0.00014572 0 0.00014564 0 0.00014574 3.3 0.00014565999999999998 3.3 0.00014576 0 0.00014568 0 0.00014578 3.3 0.0001457 3.3 0.0001458 0 0.00014572 0 0.00014582 3.3 0.00014574 3.3 0.00014584 0 0.00014576 0 0.00014586 3.3 0.00014578 3.3 0.00014588 0 0.0001458 0 0.0001459 3.3 0.00014581999999999998 3.3 0.00014591999999999999 0 0.00014584 0 0.00014594 3.3 0.00014586 3.3 0.00014596 0 0.00014588 0 0.00014598 3.3 0.0001459 3.3 0.000146 0 0.00014591999999999999 0 0.00014602 3.3 0.00014594 3.3 0.00014604 0 0.00014596 0 0.00014606 3.3 0.00014597999999999998 3.3 0.00014607999999999998 0 0.000146 0 0.0001461 3.3 0.00014602 3.3 0.00014612 0 0.00014604 0 0.00014614 3.3 0.00014606 3.3 0.00014616 0 0.00014607999999999998 0 0.00014617999999999999 3.3 0.0001461 3.3 0.0001462 0 0.00014612 0 0.00014622 3.3 0.00014614 3.3 0.00014624 0 0.00014616 0 0.00014626 3.3 0.00014617999999999999 3.3 0.00014628 0 0.0001462 0 0.0001463 3.3 0.00014622 3.3 0.00014632 0 0.00014623999999999998 0 0.00014633999999999998 3.3 0.00014626 3.3 0.00014636 0 0.00014628 0 0.00014638 3.3 0.0001463 3.3 0.0001464 0 0.00014632 0 0.00014642 3.3 0.00014633999999999998 3.3 0.00014644 0 0.00014636 0 0.00014646 3.3 0.00014638 3.3 0.00014648 0 0.0001464 0 0.0001465 3.3 0.00014642 3.3 0.00014652 0 0.00014644 0 0.00014654 3.3 0.00014646 3.3 0.00014656 0 0.00014648 0 0.00014658 3.3 0.00014649999999999998 3.3 0.00014659999999999999 0 0.00014652 0 0.00014662 3.3 0.00014654 3.3 0.00014664 0 0.00014656 0 0.00014666 3.3 0.00014658 3.3 0.00014668 0 0.00014659999999999999 0 0.0001467 3.3 0.00014662 3.3 0.00014672 0 0.00014664 0 0.00014674 3.3 0.00014665999999999998 3.3 0.00014675999999999998 0 0.00014668 0 0.00014678 3.3 0.0001467 3.3 0.0001468 0 0.00014672 0 0.00014682 3.3 0.00014674 3.3 0.00014684 0 0.00014675999999999998 0 0.00014685999999999999 3.3 0.00014678 3.3 0.00014688 0 0.0001468 0 0.0001469 3.3 0.00014682 3.3 0.00014692 0 0.00014684 0 0.00014694 3.3 0.00014685999999999999 3.3 0.00014696 0 0.00014688 0 0.00014698 3.3 0.0001469 3.3 0.000147 0 0.00014691999999999998 0 0.00014701999999999998 3.3 0.00014694 3.3 0.00014704 0 0.00014696 0 0.00014706 3.3 0.00014698 3.3 0.00014708 0 0.000147 0 0.0001471 3.3 0.00014701999999999998 3.3 0.00014712 0 0.00014704 0 0.00014714 3.3 0.00014706 3.3 0.00014716 0 0.00014708 0 0.00014718 3.3 0.0001471 3.3 0.0001472 0 0.00014712 0 0.00014722 3.3 0.00014714 3.3 0.00014724 0 0.00014716 0 0.00014726 3.3 0.00014717999999999998 3.3 0.00014727999999999999 0 0.0001472 0 0.0001473 3.3 0.00014722 3.3 0.00014732 0 0.00014724 0 0.00014734 3.3 0.00014726 3.3 0.00014736 0 0.00014727999999999999 0 0.00014738 3.3 0.0001473 3.3 0.0001474 0 0.00014732 0 0.00014742 3.3 0.00014733999999999998 3.3 0.00014743999999999998 0 0.00014736 0 0.00014746 3.3 0.00014738 3.3 0.00014748 0 0.0001474 0 0.0001475 3.3 0.00014742 3.3 0.00014752 0 0.00014743999999999998 0 0.00014754 3.3 0.00014746 3.3 0.00014756 0 0.00014748 0 0.00014758 3.3 0.0001475 3.3 0.0001476 0 0.00014752 0 0.00014762 3.3 0.00014754 3.3 0.00014764 0 0.00014756 0 0.00014766 3.3 0.00014758 3.3 0.00014768 0 0.00014759999999999998 0 0.00014769999999999999 3.3 0.00014762 3.3 0.00014772 0 0.00014764 0 0.00014774 3.3 0.00014766 3.3 0.00014776 0 0.00014768 0 0.00014778 3.3 0.00014769999999999999 3.3 0.0001478 0 0.00014772 0 0.00014782 3.3 0.00014774 3.3 0.00014784 0 0.00014775999999999998 0 0.00014785999999999998 3.3 0.00014778 3.3 0.00014788 0 0.0001478 0 0.0001479 3.3 0.00014782 3.3 0.00014792 0 0.00014784 0 0.00014794 3.3 0.00014785999999999998 3.3 0.00014795999999999999 0 0.00014788 0 0.00014798 3.3 0.0001479 3.3 0.000148 0 0.00014792 0 0.00014802 3.3 0.00014794 3.3 0.00014804 0 0.00014795999999999999 0 0.00014806 3.3 0.00014798 3.3 0.00014808 0 0.000148 0 0.0001481 3.3 0.00014801999999999998 3.3 0.00014811999999999998 0 0.00014804 0 0.00014814 3.3 0.00014806 3.3 0.00014816 0 0.00014808 0 0.00014818 3.3 0.0001481 3.3 0.0001482 0 0.00014811999999999998 0 0.00014822 3.3 0.00014814 3.3 0.00014824 0 0.00014816 0 0.00014826 3.3 0.00014818 3.3 0.00014828 0 0.0001482 0 0.0001483 3.3 0.00014822 3.3 0.00014832 0 0.00014824 0 0.00014834 3.3 0.00014826 3.3 0.00014836 0 0.00014827999999999998 0 0.00014837999999999999 3.3 0.0001483 3.3 0.0001484 0 0.00014832 0 0.00014842 3.3 0.00014834 3.3 0.00014844 0 0.00014836 0 0.00014846 3.3 0.00014837999999999999 3.3 0.00014848 0 0.0001484 0 0.0001485 3.3 0.00014842 3.3 0.00014852 0 0.00014843999999999998 0 0.00014853999999999998 3.3 0.00014846 3.3 0.00014856 0 0.00014848 0 0.00014858 3.3 0.0001485 3.3 0.0001486 0 0.00014852 0 0.00014862 3.3 0.00014853999999999998 3.3 0.00014863999999999999 0 0.00014856 0 0.00014866 3.3 0.00014858 3.3 0.00014868 0 0.0001486 0 0.0001487 3.3 0.00014862 3.3 0.00014872 0 0.00014863999999999999 0 0.00014874 3.3 0.00014866 3.3 0.00014876 0 0.00014868 0 0.00014878 3.3 0.00014869999999999998 3.3 0.00014879999999999998 0 0.00014872 0 0.00014882 3.3 0.00014874 3.3 0.00014884 0 0.00014876 0 0.00014886 3.3 0.00014878 3.3 0.00014888 0 0.00014879999999999998 0 0.0001489 3.3 0.00014882 3.3 0.00014892 0 0.00014884 0 0.00014894 3.3 0.00014886 3.3 0.00014896 0 0.00014888 0 0.00014898 3.3 0.0001489 3.3 0.000149 0 0.00014892 0 0.00014902 3.3 0.00014894 3.3 0.00014904 0 0.00014895999999999998 0 0.00014905999999999999 3.3 0.00014898 3.3 0.00014908 0 0.000149 0 0.0001491 3.3 0.00014902 3.3 0.00014912 0 0.00014904 0 0.00014914 3.3 0.00014905999999999999 3.3 0.00014916 0 0.00014908 0 0.00014918 3.3 0.0001491 3.3 0.0001492 0 0.00014911999999999998 0 0.00014921999999999998 3.3 0.00014914 3.3 0.00014924 0 0.00014916 0 0.00014926 3.3 0.00014918 3.3 0.00014928 0 0.0001492 0 0.0001493 3.3 0.00014921999999999998 3.3 0.00014932 0 0.00014924 0 0.00014934 3.3 0.00014926 3.3 0.00014936 0 0.00014928 0 0.00014938 3.3 0.0001493 3.3 0.0001494 0 0.00014932 0 0.00014942 3.3 0.00014934 3.3 0.00014944 0 0.00014936 0 0.00014946 3.3 0.00014937999999999998 3.3 0.00014947999999999999 0 0.0001494 0 0.0001495 3.3 0.00014942 3.3 0.00014952 0 0.00014944 0 0.00014954 3.3 0.00014946 3.3 0.00014956 0 0.00014947999999999999 0 0.00014958 3.3 0.0001495 3.3 0.0001496 0 0.00014952 0 0.00014962 3.3 0.00014953999999999998 3.3 0.00014963999999999998 0 0.00014956 0 0.00014966 3.3 0.00014958 3.3 0.00014968 0 0.0001496 0 0.0001497 3.3 0.00014962 3.3 0.00014972 0 0.00014963999999999998 0 0.00014973999999999999 3.3 0.00014966 3.3 0.00014976 0 0.00014968 0 0.00014978 3.3 0.0001497 3.3 0.0001498 0 0.00014972 0 0.00014982 3.3 0.00014973999999999999 3.3 0.00014984 0 0.00014976 0 0.00014986 3.3 0.00014978 3.3 0.00014988 0 0.00014979999999999998 0 0.00014989999999999998 3.3 0.00014982 3.3 0.00014992 0 0.00014984 0 0.00014994 3.3 0.00014986 3.3 0.00014996 0 0.00014988 0 0.00014998 3.3 0.00014989999999999998 3.3 0.00015 0 0.00014992 0 0.00015002 3.3 0.00014994 3.3 0.00015004 0 0.00014996 0 0.00015006 3.3 0.00014998 3.3 0.00015008 0 0.00015 0 0.0001501 3.3 0.00015002 3.3 0.00015012 0 0.00015004 0 0.00015014 3.3 0.00015005999999999998 3.3 0.00015015999999999999 0 0.00015008 0 0.00015018 3.3 0.0001501 3.3 0.0001502 0 0.00015012 0 0.00015022 3.3 0.00015014 3.3 0.00015024 0 0.00015015999999999999 0 0.00015026 3.3 0.00015018 3.3 0.00015028 0 0.0001502 0 0.0001503 3.3 0.00015021999999999998 3.3 0.00015031999999999998 0 0.00015024 0 0.00015034 3.3 0.00015026 3.3 0.00015036 0 0.00015028 0 0.00015038 3.3 0.0001503 3.3 0.0001504 0 0.00015031999999999998 0 0.00015041999999999999 3.3 0.00015034 3.3 0.00015044 0 0.00015036 0 0.00015046 3.3 0.00015038 3.3 0.00015048 0 0.0001504 0 0.0001505 3.3 0.00015041999999999999 3.3 0.00015052 0 0.00015044 0 0.00015054 3.3 0.00015046 3.3 0.00015056 0 0.00015047999999999998 0 0.00015057999999999998 3.3 0.0001505 3.3 0.0001506 0 0.00015052 0 0.00015062 3.3 0.00015054 3.3 0.00015064 0 0.00015056 0 0.00015066 3.3 0.00015057999999999998 3.3 0.00015068 0 0.0001506 0 0.0001507 3.3 0.00015062 3.3 0.00015072 0 0.00015064 0 0.00015074 3.3 0.00015066 3.3 0.00015076 0 0.00015068 0 0.00015078 3.3 0.0001507 3.3 0.0001508 0 0.00015072 0 0.00015082 3.3 0.00015073999999999998 3.3 0.00015083999999999999 0 0.00015076 0 0.00015086 3.3 0.00015078 3.3 0.00015088 0 0.0001508 0 0.0001509 3.3 0.00015082 3.3 0.00015092 0 0.00015083999999999999 0 0.00015094 3.3 0.00015086 3.3 0.00015096 0 0.00015088 0 0.00015098 3.3 0.00015089999999999998 3.3 0.00015099999999999998 0 0.00015092 0 0.00015102 3.3 0.00015094 3.3 0.00015104 0 0.00015096 0 0.00015106 3.3 0.00015098 3.3 0.00015108 0 0.00015099999999999998 0 0.0001511 3.3 0.00015102 3.3 0.00015112 0 0.00015104 0 0.00015114 3.3 0.00015106 3.3 0.00015116 0 0.00015108 0 0.00015118 3.3 0.0001511 3.3 0.0001512 0 0.00015112 0 0.00015122 3.3 0.00015114 3.3 0.00015124 0 0.00015115999999999998 0 0.00015125999999999998 3.3 0.00015118 3.3 0.00015128 0 0.0001512 0 0.0001513 3.3 0.00015122 3.3 0.00015132 0 0.00015124 0 0.00015134 3.3 0.00015125999999999998 3.3 0.00015136 0 0.00015128 0 0.00015138 3.3 0.0001513 3.3 0.0001514 0 0.00015131999999999998 0 0.00015141999999999998 3.3 0.00015134 3.3 0.00015144 0 0.00015136 0 0.00015146 3.3 0.00015138 3.3 0.00015148 0 0.0001514 0 0.0001515 3.3 0.00015141999999999998 3.3 0.00015151999999999999 0 0.00015144 0 0.00015154 3.3 0.00015146 3.3 0.00015156 0 0.00015148 0 0.00015158 3.3 0.0001515 3.3 0.0001516 0 0.00015151999999999999 0 0.00015162 3.3 0.00015154 3.3 0.00015164 0 0.00015156 0 0.00015166 3.3 0.00015157999999999998 3.3 0.00015167999999999998 0 0.0001516 0 0.0001517 3.3 0.00015162 3.3 0.00015172 0 0.00015164 0 0.00015174 3.3 0.00015166 3.3 0.00015176 0 0.00015167999999999998 0 0.00015178 3.3 0.0001517 3.3 0.0001518 0 0.00015172 0 0.00015182 3.3 0.00015174 3.3 0.00015184 0 0.00015176 0 0.00015186 3.3 0.00015178 3.3 0.00015188 0 0.0001518 0 0.0001519 3.3 0.00015182 3.3 0.00015192 0 0.00015183999999999998 0 0.00015193999999999999 3.3 0.00015186 3.3 0.00015196 0 0.00015188 0 0.00015198 3.3 0.0001519 3.3 0.000152 0 0.00015192 0 0.00015202 3.3 0.00015193999999999999 3.3 0.00015204 0 0.00015196 0 0.00015206 3.3 0.00015198 3.3 0.00015208 0 0.00015199999999999998 0 0.00015209999999999998 3.3 0.00015202 3.3 0.00015212 0 0.00015204 0 0.00015214 3.3 0.00015206 3.3 0.00015216 0 0.00015208 0 0.00015218 3.3 0.00015209999999999998 3.3 0.00015219999999999999 0 0.00015212 0 0.00015222 3.3 0.00015214 3.3 0.00015224 0 0.00015216 0 0.00015226 3.3 0.00015218 3.3 0.00015228 0 0.00015219999999999999 0 0.0001523 3.3 0.00015222 3.3 0.00015232 0 0.00015224 0 0.00015234 3.3 0.00015225999999999998 3.3 0.00015235999999999998 0 0.00015228 0 0.00015238 3.3 0.0001523 3.3 0.0001524 0 0.00015232 0 0.00015242 3.3 0.00015234 3.3 0.00015244 0 0.00015235999999999998 0 0.00015246 3.3 0.00015238 3.3 0.00015248 0 0.0001524 0 0.0001525 3.3 0.00015242 3.3 0.00015252 0 0.00015244 0 0.00015254 3.3 0.00015246 3.3 0.00015256 0 0.00015248 0 0.00015258 3.3 0.0001525 3.3 0.0001526 0 0.00015251999999999998 0 0.00015261999999999999 3.3 0.00015254 3.3 0.00015264 0 0.00015256 0 0.00015266 3.3 0.00015258 3.3 0.00015268 0 0.0001526 0 0.0001527 3.3 0.00015261999999999999 3.3 0.00015272 0 0.00015264 0 0.00015274 3.3 0.00015266 3.3 0.00015276 0 0.00015267999999999998 0 0.00015277999999999998 3.3 0.0001527 3.3 0.0001528 0 0.00015272 0 0.00015282 3.3 0.00015274 3.3 0.00015284 0 0.00015276 0 0.00015286 3.3 0.00015277999999999998 3.3 0.00015287999999999999 0 0.0001528 0 0.0001529 3.3 0.00015282 3.3 0.00015292 0 0.00015284 0 0.00015294 3.3 0.00015286 3.3 0.00015296 0 0.00015287999999999999 0 0.00015298 3.3 0.0001529 3.3 0.000153 0 0.00015292 0 0.00015302 3.3 0.00015293999999999998 3.3 0.00015303999999999998 0 0.00015296 0 0.00015306 3.3 0.00015298 3.3 0.00015308 0 0.000153 0 0.0001531 3.3 0.00015302 3.3 0.00015312 0 0.00015303999999999998 0 0.00015314 3.3 0.00015306 3.3 0.00015316 0 0.00015308 0 0.00015318 3.3 0.0001531 3.3 0.0001532 0 0.00015312 0 0.00015322 3.3 0.00015314 3.3 0.00015324 0 0.00015316 0 0.00015326 3.3 0.00015318 3.3 0.00015328 0 0.00015319999999999998 0 0.00015329999999999999 3.3 0.00015322 3.3 0.00015332 0 0.00015324 0 0.00015334 3.3 0.00015326 3.3 0.00015336 0 0.00015328 0 0.00015338 3.3 0.00015329999999999999 3.3 0.0001534 0 0.00015332 0 0.00015342 3.3 0.00015334 3.3 0.00015344 0 0.00015335999999999998 0 0.00015345999999999998 3.3 0.00015338 3.3 0.00015348 0 0.0001534 0 0.0001535 3.3 0.00015342 3.3 0.00015352 0 0.00015344 0 0.00015354 3.3 0.00015345999999999998 3.3 0.00015356 0 0.00015348 0 0.00015358 3.3 0.0001535 3.3 0.0001536 0 0.00015352 0 0.00015362 3.3 0.00015354 3.3 0.00015364 0 0.00015356 0 0.00015366 3.3 0.00015358 3.3 0.00015368 0 0.0001536 0 0.0001537 3.3 0.00015361999999999998 3.3 0.00015371999999999999 0 0.00015364 0 0.00015374 3.3 0.00015366 3.3 0.00015376 0 0.00015368 0 0.00015378 3.3 0.0001537 3.3 0.0001538 0 0.00015371999999999999 0 0.00015382 3.3 0.00015374 3.3 0.00015384 0 0.00015376 0 0.00015386 3.3 0.00015377999999999998 3.3 0.00015387999999999998 0 0.0001538 0 0.0001539 3.3 0.00015382 3.3 0.00015392 0 0.00015384 0 0.00015394 3.3 0.00015386 3.3 0.00015396 0 0.00015387999999999998 0 0.00015397999999999999 3.3 0.0001539 3.3 0.000154 0 0.00015392 0 0.00015402 3.3 0.00015394 3.3 0.00015404 0 0.00015396 0 0.00015406 3.3 0.00015397999999999999 3.3 0.00015408 0 0.000154 0 0.0001541 3.3 0.00015402 3.3 0.00015412 0 0.00015403999999999998 0 0.00015413999999999998 3.3 0.00015406 3.3 0.00015416 0 0.00015408 0 0.00015418 3.3 0.0001541 3.3 0.0001542 0 0.00015412 0 0.00015422 3.3 0.00015413999999999998 3.3 0.00015424 0 0.00015416 0 0.00015426 3.3 0.00015418 3.3 0.00015428 0 0.0001542 0 0.0001543 3.3 0.00015422 3.3 0.00015432 0 0.00015424 0 0.00015434 3.3 0.00015426 3.3 0.00015436 0 0.00015428 0 0.00015438 3.3 0.00015429999999999998 3.3 0.00015439999999999999 0 0.00015432 0 0.00015442 3.3 0.00015434 3.3 0.00015444 0 0.00015436 0 0.00015446 3.3 0.00015438 3.3 0.00015448 0 0.00015439999999999999 0 0.0001545 3.3 0.00015442 3.3 0.00015452 0 0.00015444 0 0.00015454 3.3 0.00015445999999999998 3.3 0.00015455999999999998 0 0.00015448 0 0.00015458 3.3 0.0001545 3.3 0.0001546 0 0.00015452 0 0.00015462 3.3 0.00015454 3.3 0.00015464 0 0.00015455999999999998 0 0.00015465999999999999 3.3 0.00015458 3.3 0.00015468 0 0.0001546 0 0.0001547 3.3 0.00015462 3.3 0.00015472 0 0.00015464 0 0.00015474 3.3 0.00015465999999999999 3.3 0.00015476 0 0.00015468 0 0.00015478 3.3 0.0001547 3.3 0.0001548 0 0.00015471999999999998 0 0.00015481999999999998 3.3 0.00015474 3.3 0.00015484 0 0.00015476 0 0.00015486 3.3 0.00015478 3.3 0.00015488 0 0.0001548 0 0.0001549 3.3 0.00015481999999999998 3.3 0.00015492 0 0.00015484 0 0.00015494 3.3 0.00015486 3.3 0.00015496 0 0.00015488 0 0.00015498 3.3 0.0001549 3.3 0.000155 0 0.00015492 0 0.00015502 3.3 0.00015494 3.3 0.00015504 0 0.00015496 0 0.00015506 3.3 0.00015497999999999998 3.3 0.00015507999999999999 0 0.000155 0 0.0001551 3.3 0.00015502 3.3 0.00015512 0 0.00015504 0 0.00015514 3.3 0.00015506 3.3 0.00015516 0 0.00015507999999999999 0 0.00015518 3.3 0.0001551 3.3 0.0001552 0 0.00015512 0 0.00015522 3.3 0.00015513999999999998 3.3 0.00015523999999999998 0 0.00015516 0 0.00015526 3.3 0.00015518 3.3 0.00015528 0 0.0001552 0 0.0001553 3.3 0.00015522 3.3 0.00015532 0 0.00015523999999999998 0 0.00015534 3.3 0.00015526 3.3 0.00015536 0 0.00015528 0 0.00015538 3.3 0.0001553 3.3 0.0001554 0 0.00015532 0 0.00015542 3.3 0.00015534 3.3 0.00015544 0 0.00015536 0 0.00015546 3.3 0.00015538 3.3 0.00015548 0 0.00015539999999999998 0 0.00015549999999999999 3.3 0.00015542 3.3 0.00015552 0 0.00015544 0 0.00015554 3.3 0.00015546 3.3 0.00015556 0 0.00015548 0 0.00015558 3.3 0.00015549999999999999 3.3 0.0001556 0 0.00015552 0 0.00015562 3.3 0.00015554 3.3 0.00015564 0 0.00015555999999999998 0 0.00015565999999999998 3.3 0.00015558 3.3 0.00015568 0 0.0001556 0 0.0001557 3.3 0.00015562 3.3 0.00015572 0 0.00015564 0 0.00015574 3.3 0.00015565999999999998 3.3 0.00015575999999999999 0 0.00015568 0 0.00015578 3.3 0.0001557 3.3 0.0001558 0 0.00015572 0 0.00015582 3.3 0.00015574 3.3 0.00015584 0 0.00015575999999999999 0 0.00015586 3.3 0.00015578 3.3 0.00015588 0 0.0001558 0 0.0001559 3.3 0.00015581999999999998 3.3 0.00015591999999999998 0 0.00015584 0 0.00015594 3.3 0.00015586 3.3 0.00015596 0 0.00015588 0 0.00015598 3.3 0.0001559 3.3 0.000156 0 0.00015591999999999998 0 0.00015602 3.3 0.00015594 3.3 0.00015604 0 0.00015596 0 0.00015606 3.3 0.00015598 3.3 0.00015608 0 0.000156 0 0.0001561 3.3 0.00015602 3.3 0.00015612 0 0.00015604 0 0.00015614 3.3 0.00015606 3.3 0.00015616 0 0.00015607999999999998 0 0.00015617999999999999 3.3 0.0001561 3.3 0.0001562 0 0.00015612 0 0.00015622 3.3 0.00015614 3.3 0.00015624 0 0.00015616 0 0.00015626 3.3 0.00015617999999999999 3.3 0.00015628 0 0.0001562 0 0.0001563 3.3 0.00015622 3.3 0.00015632 0 0.00015623999999999998 0 0.00015633999999999998 3.3 0.00015626 3.3 0.00015636 0 0.00015628 0 0.00015638 3.3 0.0001563 3.3 0.0001564 0 0.00015632 0 0.00015642 3.3 0.00015633999999999998 3.3 0.00015643999999999999 0 0.00015636 0 0.00015646 3.3 0.00015638 3.3 0.00015648 0 0.0001564 0 0.0001565 3.3 0.00015642 3.3 0.00015652 0 0.00015643999999999999 0 0.00015654 3.3 0.00015646 3.3 0.00015656 0 0.00015648 0 0.00015658 3.3 0.00015649999999999998 3.3 0.00015659999999999998 0 0.00015652 0 0.00015662 3.3 0.00015654 3.3 0.00015664 0 0.00015656 0 0.00015666 3.3 0.00015658 3.3 0.00015668 0 0.00015659999999999998 0 0.0001567 3.3 0.00015662 3.3 0.00015672 0 0.00015664 0 0.00015674 3.3 0.00015666 3.3 0.00015676 0 0.00015668 0 0.00015678 3.3 0.0001567 3.3 0.0001568 0 0.00015672 0 0.00015682 3.3 0.00015674 3.3 0.00015684 0 0.00015675999999999998 0 0.00015685999999999999 3.3 0.00015678 3.3 0.00015688 0 0.0001568 0 0.0001569 3.3 0.00015682 3.3 0.00015692 0 0.00015684 0 0.00015694 3.3 0.00015685999999999999 3.3 0.00015696 0 0.00015688 0 0.00015698 3.3 0.0001569 3.3 0.000157 0 0.00015691999999999998 0 0.00015701999999999998 3.3 0.00015694 3.3 0.00015704 0 0.00015696 0 0.00015706 3.3 0.00015698 3.3 0.00015708 0 0.000157 0 0.0001571 3.3 0.00015701999999999998 3.3 0.00015712 0 0.00015704 0 0.00015714 3.3 0.00015706 3.3 0.00015716 0 0.00015708 0 0.00015718 3.3 0.0001571 3.3 0.0001572 0 0.00015712 0 0.00015722 3.3 0.00015714 3.3 0.00015724 0 0.00015716 0 0.00015726 3.3 0.00015717999999999998 3.3 0.00015727999999999998 0 0.0001572 0 0.0001573 3.3 0.00015722 3.3 0.00015732 0 0.00015724 0 0.00015734 3.3 0.00015726 3.3 0.00015736 0 0.00015727999999999998 0 0.00015738 3.3 0.0001573 3.3 0.0001574 0 0.00015732 0 0.00015742 3.3 0.00015733999999999998 3.3 0.00015743999999999998 0 0.00015736 0 0.00015746 3.3 0.00015738 3.3 0.00015748 0 0.0001574 0 0.0001575 3.3 0.00015742 3.3 0.00015752 0 0.00015743999999999998 0 0.00015753999999999999 3.3 0.00015746 3.3 0.00015756 0 0.00015748 0 0.00015758 3.3 0.0001575 3.3 0.0001576 0 0.00015752 0 0.00015762 3.3 0.00015753999999999999 3.3 0.00015764 0 0.00015756 0 0.00015766 3.3 0.00015758 3.3 0.00015768 0 0.00015759999999999998 0 0.00015769999999999998 3.3 0.00015762 3.3 0.00015772 0 0.00015764 0 0.00015774 3.3 0.00015766 3.3 0.00015776 0 0.00015768 0 0.00015778 3.3 0.00015769999999999998 3.3 0.0001578 0 0.00015772 0 0.00015782 3.3 0.00015774 3.3 0.00015784 0 0.00015776 0 0.00015786 3.3 0.00015778 3.3 0.00015788 0 0.0001578 0 0.0001579 3.3 0.00015782 3.3 0.00015792 0 0.00015784 0 0.00015794 3.3 0.00015785999999999998 3.3 0.00015795999999999999 0 0.00015788 0 0.00015798 3.3 0.0001579 3.3 0.000158 0 0.00015792 0 0.00015802 3.3 0.00015794 3.3 0.00015804 0 0.00015795999999999999 0 0.00015806 3.3 0.00015798 3.3 0.00015808 0 0.000158 0 0.0001581 3.3 0.00015801999999999998 3.3 0.00015811999999999998 0 0.00015804 0 0.00015814 3.3 0.00015806 3.3 0.00015816 0 0.00015808 0 0.00015818 3.3 0.0001581 3.3 0.0001582 0 0.00015811999999999998 0 0.00015821999999999999 3.3 0.00015814 3.3 0.00015824 0 0.00015816 0 0.00015826 3.3 0.00015818 3.3 0.00015828 0 0.0001582 0 0.0001583 3.3 0.00015821999999999999 3.3 0.00015832 0 0.00015824 0 0.00015834 3.3 0.00015826 3.3 0.00015836 0 0.00015827999999999998 0 0.00015837999999999998 3.3 0.0001583 3.3 0.0001584 0 0.00015832 0 0.00015842 3.3 0.00015834 3.3 0.00015844 0 0.00015836 0 0.00015846 3.3 0.00015837999999999998 3.3 0.00015848 0 0.0001584 0 0.0001585 3.3 0.00015842 3.3 0.00015852 0 0.00015844 0 0.00015854 3.3 0.00015846 3.3 0.00015856 0 0.00015848 0 0.00015858 3.3 0.0001585 3.3 0.0001586 0 0.00015852 0 0.00015862 3.3 0.00015853999999999998 3.3 0.00015863999999999999 0 0.00015856 0 0.00015866 3.3 0.00015858 3.3 0.00015868 0 0.0001586 0 0.0001587 3.3 0.00015862 3.3 0.00015872 0 0.00015863999999999999 0 0.00015874 3.3 0.00015866 3.3 0.00015876 0 0.00015868 0 0.00015878 3.3 0.00015869999999999998 3.3 0.00015879999999999998 0 0.00015872 0 0.00015882 3.3 0.00015874 3.3 0.00015884 0 0.00015876 0 0.00015886 3.3 0.00015878 3.3 0.00015888 0 0.00015879999999999998 0 0.00015889999999999999 3.3 0.00015882 3.3 0.00015892 0 0.00015884 0 0.00015894 3.3 0.00015886 3.3 0.00015896 0 0.00015888 0 0.00015898 3.3 0.00015889999999999999 3.3 0.000159 0 0.00015892 0 0.00015902 3.3 0.00015894 3.3 0.00015904 0 0.00015895999999999998 0 0.00015905999999999998 3.3 0.00015898 3.3 0.00015908 0 0.000159 0 0.0001591 3.3 0.00015902 3.3 0.00015912 0 0.00015904 0 0.00015914 3.3 0.00015905999999999998 3.3 0.00015916 0 0.00015908 0 0.00015918 3.3 0.0001591 3.3 0.0001592 0 0.00015911999999999998 0 0.00015921999999999998 3.3 0.00015914 3.3 0.00015924 0 0.00015916 0 0.00015926 3.3 0.00015918 3.3 0.00015928 0 0.0001592 0 0.0001593 3.3 0.00015921999999999998 3.3 0.00015931999999999999 0 0.00015924 0 0.00015934 3.3 0.00015926 3.3 0.00015936 0 0.00015928 0 0.00015938 3.3 0.0001593 3.3 0.0001594 0 0.00015931999999999999 0 0.00015942 3.3 0.00015934 3.3 0.00015944 0 0.00015936 0 0.00015946 3.3 0.00015937999999999998 3.3 0.00015947999999999998 0 0.0001594 0 0.0001595 3.3 0.00015942 3.3 0.00015952 0 0.00015944 0 0.00015954 3.3 0.00015946 3.3 0.00015956 0 0.00015947999999999998 0 0.00015958 3.3 0.0001595 3.3 0.0001596 0 0.00015952 0 0.00015962 3.3 0.00015954 3.3 0.00015964 0 0.00015956 0 0.00015966 3.3 0.00015958 3.3 0.00015968 0 0.0001596 0 0.0001597 3.3 0.00015962 3.3 0.00015972 0 0.00015963999999999998 0 0.00015973999999999999 3.3 0.00015966 3.3 0.00015976 0 0.00015968 0 0.00015978 3.3 0.0001597 3.3 0.0001598 0 0.00015972 0 0.00015982 3.3 0.00015973999999999999 3.3 0.00015984 0 0.00015976 0 0.00015986 3.3 0.00015978 3.3 0.00015988 0 0.00015979999999999998 0 0.00015989999999999998 3.3 0.00015982 3.3 0.00015992 0 0.00015984 0 0.00015994 3.3 0.00015986 3.3 0.00015996 0 0.00015988 0 0.00015998 3.3 0.00015989999999999998 3.3 0.00015999999999999999 0 0.00015992 0 0.00016002 3.3 0.00015994 3.3 0.00016004 0 0.00015996 0 0.00016006 3.3 0.00015998 3.3 0.00016008 0 0.00015999999999999999 0 0.0001601 3.3 0.00016002 3.3 0.00016012 0 0.00016004 0 0.00016014 3.3 0.00016005999999999998 3.3 0.00016015999999999998 0 0.00016008 0 0.00016018 3.3 0.0001601 3.3 0.0001602 0 0.00016012 0 0.00016022 3.3 0.00016014 3.3 0.00016024 0 0.00016015999999999998 0 0.00016026 3.3 0.00016018 3.3 0.00016028 0 0.0001602 0 0.0001603 3.3 0.00016022 3.3 0.00016032 0 0.00016024 0 0.00016034 3.3 0.00016026 3.3 0.00016036 0 0.00016028 0 0.00016038 3.3 0.0001603 3.3 0.0001604 0 0.00016031999999999998 0 0.00016041999999999999 3.3 0.00016034 3.3 0.00016044 0 0.00016036 0 0.00016046 3.3 0.00016038 3.3 0.00016048 0 0.0001604 0 0.0001605 3.3 0.00016041999999999999 3.3 0.00016052 0 0.00016044 0 0.00016054 3.3 0.00016046 3.3 0.00016056 0 0.00016047999999999998 0 0.00016057999999999998 3.3 0.0001605 3.3 0.0001606 0 0.00016052 0 0.00016062 3.3 0.00016054 3.3 0.00016064 0 0.00016056 0 0.00016066 3.3 0.00016057999999999998 3.3 0.00016067999999999999 0 0.0001606 0 0.0001607 3.3 0.00016062 3.3 0.00016072 0 0.00016064 0 0.00016074 3.3 0.00016066 3.3 0.00016076 0 0.00016067999999999999 0 0.00016078 3.3 0.0001607 3.3 0.0001608 0 0.00016072 0 0.00016082 3.3 0.00016073999999999998 3.3 0.00016083999999999998 0 0.00016076 0 0.00016086 3.3 0.00016078 3.3 0.00016088 0 0.0001608 0 0.0001609 3.3 0.00016082 3.3 0.00016092 0 0.00016083999999999998 0 0.00016094 3.3 0.00016086 3.3 0.00016096 0 0.00016088 0 0.00016098 3.3 0.0001609 3.3 0.000161 0 0.00016092 0 0.00016102 3.3 0.00016094 3.3 0.00016104 0 0.00016096 0 0.00016106 3.3 0.00016098 3.3 0.00016108 0 0.00016099999999999998 0 0.00016109999999999999 3.3 0.00016102 3.3 0.00016112 0 0.00016104 0 0.00016114 3.3 0.00016106 3.3 0.00016116 0 0.00016108 0 0.00016118 3.3 0.00016109999999999999 3.3 0.0001612 0 0.00016112 0 0.00016122 3.3 0.00016114 3.3 0.00016124 0 0.00016115999999999998 0 0.00016125999999999998 3.3 0.00016118 3.3 0.00016128 0 0.0001612 0 0.0001613 3.3 0.00016122 3.3 0.00016132 0 0.00016124 0 0.00016134 3.3 0.00016125999999999998 3.3 0.00016136 0 0.00016128 0 0.00016138 3.3 0.0001613 3.3 0.0001614 0 0.00016132 0 0.00016142 3.3 0.00016134 3.3 0.00016144 0 0.00016136 0 0.00016146 3.3 0.00016138 3.3 0.00016148 0 0.0001614 0 0.0001615 3.3 0.00016141999999999998 3.3 0.00016151999999999998 0 0.00016144 0 0.00016154 3.3 0.00016146 3.3 0.00016156 0 0.00016148 0 0.00016158 3.3 0.0001615 3.3 0.0001616 0 0.00016151999999999998 0 0.00016162 3.3 0.00016154 3.3 0.00016164 0 0.00016156 0 0.00016166 3.3 0.00016157999999999998 3.3 0.00016167999999999998 0 0.0001616 0 0.0001617 3.3 0.00016162 3.3 0.00016172 0 0.00016164 0 0.00016174 3.3 0.00016166 3.3 0.00016176 0 0.00016167999999999998 0 0.00016177999999999999 3.3 0.0001617 3.3 0.0001618 0 0.00016172 0 0.00016182 3.3 0.00016174 3.3 0.00016184 0 0.00016176 0 0.00016186 3.3 0.00016177999999999999 3.3 0.00016188 0 0.0001618 0 0.0001619 3.3 0.00016182 3.3 0.00016192 0 0.00016183999999999998 0 0.00016193999999999998 3.3 0.00016186 3.3 0.00016196 0 0.00016188 0 0.00016198 3.3 0.0001619 3.3 0.000162 0 0.00016192 0 0.00016202 3.3 0.00016193999999999998 3.3 0.00016204 0 0.00016196 0 0.00016206 3.3 0.00016198 3.3 0.00016208 0 0.000162 0 0.0001621 3.3 0.00016202 3.3 0.00016212 0 0.00016204 0 0.00016214 3.3 0.00016206 3.3 0.00016216 0 0.00016208 0 0.00016218 3.3 0.00016209999999999998 3.3 0.00016219999999999999 0 0.00016212 0 0.00016222 3.3 0.00016214 3.3 0.00016224 0 0.00016216 0 0.00016226 3.3 0.00016218 3.3 0.00016228 0 0.00016219999999999999 0 0.0001623 3.3 0.00016222 3.3 0.00016232 0 0.00016224 0 0.00016234 3.3 0.00016225999999999998 3.3 0.00016235999999999998 0 0.00016228 0 0.00016238 3.3 0.0001623 3.3 0.0001624 0 0.00016232 0 0.00016242 3.3 0.00016234 3.3 0.00016244 0 0.00016235999999999998 0 0.00016245999999999999 3.3 0.00016238 3.3 0.00016248 0 0.0001624 0 0.0001625 3.3 0.00016242 3.3 0.00016252 0 0.00016244 0 0.00016254 3.3 0.00016245999999999999 3.3 0.00016256 0 0.00016248 0 0.00016258 3.3 0.0001625 3.3 0.0001626 0 0.00016251999999999998 0 0.00016261999999999998 3.3 0.00016254 3.3 0.00016264 0 0.00016256 0 0.00016266 3.3 0.00016258 3.3 0.00016268 0 0.0001626 0 0.0001627 3.3 0.00016261999999999998 3.3 0.00016272 0 0.00016264 0 0.00016274 3.3 0.00016266 3.3 0.00016276 0 0.00016268 0 0.00016278 3.3 0.0001627 3.3 0.0001628 0 0.00016272 0 0.00016282 3.3 0.00016274 3.3 0.00016284 0 0.00016276 0 0.00016286 3.3 0.00016277999999999998 3.3 0.00016287999999999999 0 0.0001628 0 0.0001629 3.3 0.00016282 3.3 0.00016292 0 0.00016284 0 0.00016294 3.3 0.00016286 3.3 0.00016296 0 0.00016287999999999999 0 0.00016298 3.3 0.0001629 3.3 0.000163 0 0.00016292 0 0.00016302 3.3 0.00016293999999999998 3.3 0.00016303999999999998 0 0.00016296 0 0.00016306 3.3 0.00016298 3.3 0.00016308 0 0.000163 0 0.0001631 3.3 0.00016302 3.3 0.00016312 0 0.00016303999999999998 0 0.00016313999999999999 3.3 0.00016306 3.3 0.00016316 0 0.00016308 0 0.00016318 3.3 0.0001631 3.3 0.0001632 0 0.00016312 0 0.00016322 3.3 0.00016313999999999999 3.3 0.00016324 0 0.00016316 0 0.00016326 3.3 0.00016318 3.3 0.00016328 0 0.00016319999999999998 0 0.00016329999999999998 3.3 0.00016322 3.3 0.00016332 0 0.00016324 0 0.00016334 3.3 0.00016326 3.3 0.00016336 0 0.00016328 0 0.00016338 3.3 0.00016329999999999998 3.3 0.0001634 0 0.00016332 0 0.00016342 3.3 0.00016334 3.3 0.00016344 0 0.00016335999999999998 0 0.00016345999999999998 3.3 0.00016338 3.3 0.00016348 0 0.0001634 0 0.0001635 3.3 0.00016342 3.3 0.00016352 0 0.00016344 0 0.00016354 3.3 0.00016345999999999998 3.3 0.00016355999999999999 0 0.00016348 0 0.00016358 3.3 0.0001635 3.3 0.0001636 0 0.00016352 0 0.00016362 3.3 0.00016354 3.3 0.00016364 0 0.00016355999999999999 0 0.00016366 3.3 0.00016358 3.3 0.00016368 0 0.0001636 0 0.0001637 3.3 0.00016361999999999998 3.3 0.00016371999999999998 0 0.00016364 0 0.00016374 3.3 0.00016366 3.3 0.00016376 0 0.00016368 0 0.00016378 3.3 0.0001637 3.3 0.0001638 0 0.00016371999999999998 0 0.00016382 3.3 0.00016374 3.3 0.00016384 0 0.00016376 0 0.00016386 3.3 0.00016378 3.3 0.00016388 0 0.0001638 0 0.0001639 3.3 0.00016382 3.3 0.00016392 0 0.00016384 0 0.00016394 3.3 0.00016386 3.3 0.00016396 0 0.00016387999999999998 0 0.00016397999999999999 3.3 0.0001639 3.3 0.000164 0 0.00016392 0 0.00016402 3.3 0.00016394 3.3 0.00016404 0 0.00016396 0 0.00016406 3.3 0.00016397999999999999 3.3 0.00016408 0 0.000164 0 0.0001641 3.3 0.00016402 3.3 0.00016412 0 0.00016403999999999998 0 0.00016413999999999998 3.3 0.00016406 3.3 0.00016416 0 0.00016408 0 0.00016418 3.3 0.0001641 3.3 0.0001642 0 0.00016412 0 0.00016422 3.3 0.00016413999999999998 3.3 0.00016423999999999999 0 0.00016416 0 0.00016426 3.3 0.00016418 3.3 0.00016428 0 0.0001642 0 0.0001643 3.3 0.00016422 3.3 0.00016432 0 0.00016423999999999999 0 0.00016434 3.3 0.00016426 3.3 0.00016436 0 0.00016428 0 0.00016438 3.3 0.00016429999999999998 3.3 0.00016439999999999998 0 0.00016432 0 0.00016442 3.3 0.00016434 3.3 0.00016444 0 0.00016436 0 0.00016446 3.3 0.00016438 3.3 0.00016448 0 0.00016439999999999998 0 0.0001645 3.3 0.00016442 3.3 0.00016452 0 0.00016444 0 0.00016454 3.3 0.00016446 3.3 0.00016456 0 0.00016448 0 0.00016458 3.3 0.0001645 3.3 0.0001646 0 0.00016452 0 0.00016462 3.3 0.00016454 3.3 0.00016464 0 0.00016455999999999998 0 0.00016465999999999999 3.3 0.00016458 3.3 0.00016468 0 0.0001646 0 0.0001647 3.3 0.00016462 3.3 0.00016472 0 0.00016464 0 0.00016474 3.3 0.00016465999999999999 3.3 0.00016476 0 0.00016468 0 0.00016478 3.3 0.0001647 3.3 0.0001648 0 0.00016471999999999998 0 0.00016481999999999998 3.3 0.00016474 3.3 0.00016484 0 0.00016476 0 0.00016486 3.3 0.00016478 3.3 0.00016488 0 0.0001648 0 0.0001649 3.3 0.00016481999999999998 3.3 0.00016491999999999999 0 0.00016484 0 0.00016494 3.3 0.00016486 3.3 0.00016496 0 0.00016488 0 0.00016498 3.3 0.0001649 3.3 0.000165 0 0.00016491999999999999 0 0.00016502 3.3 0.00016494 3.3 0.00016504 0 0.00016496 0 0.00016506 3.3 0.00016497999999999998 3.3 0.00016507999999999998 0 0.000165 0 0.0001651 3.3 0.00016502 3.3 0.00016512 0 0.00016504 0 0.00016514 3.3 0.00016506 3.3 0.00016516 0 0.00016507999999999998 0 0.00016518 3.3 0.0001651 3.3 0.0001652 0 0.00016512 0 0.00016522 3.3 0.00016513999999999998 3.3 0.00016523999999999998 0 0.00016516 0 0.00016526 3.3 0.00016518 3.3 0.00016528 0 0.0001652 0 0.0001653 3.3 0.00016522 3.3 0.00016532 0 0.00016523999999999998 0 0.00016533999999999999 3.3 0.00016526 3.3 0.00016536 0 0.00016528 0 0.00016538 3.3 0.0001653 3.3 0.0001654 0 0.00016532 0 0.00016542 3.3 0.00016533999999999999 3.3 0.00016544 0 0.00016536 0 0.00016546 3.3 0.00016538 3.3 0.00016548 0 0.00016539999999999998 0 0.00016549999999999998 3.3 0.00016542 3.3 0.00016552 0 0.00016544 0 0.00016554 3.3 0.00016546 3.3 0.00016556 0 0.00016548 0 0.00016558 3.3 0.00016549999999999998 3.3 0.0001656 0 0.00016552 0 0.00016562 3.3 0.00016554 3.3 0.00016564 0 0.00016556 0 0.00016566 3.3 0.00016558 3.3 0.00016568 0 0.0001656 0 0.0001657 3.3 0.00016562 3.3 0.00016572 0 0.00016564 0 0.00016574 3.3 0.00016565999999999998 3.3 0.00016575999999999999 0 0.00016568 0 0.00016578 3.3 0.0001657 3.3 0.0001658 0 0.00016572 0 0.00016582 3.3 0.00016574 3.3 0.00016584 0 0.00016575999999999999 0 0.00016586 3.3 0.00016578 3.3 0.00016588 0 0.0001658 0 0.0001659 3.3 0.00016581999999999998 3.3 0.00016591999999999998 0 0.00016584 0 0.00016594 3.3 0.00016586 3.3 0.00016596 0 0.00016588 0 0.00016598 3.3 0.0001659 3.3 0.000166 0 0.00016591999999999998 0 0.00016601999999999999 3.3 0.00016594 3.3 0.00016604 0 0.00016596 0 0.00016606 3.3 0.00016598 3.3 0.00016608 0 0.000166 0 0.0001661 3.3 0.00016601999999999999 3.3 0.00016612 0 0.00016604 0 0.00016614 3.3 0.00016606 3.3 0.00016616 0 0.00016607999999999998 0 0.00016617999999999998 3.3 0.0001661 3.3 0.0001662 0 0.00016612 0 0.00016622 3.3 0.00016614 3.3 0.00016624 0 0.00016616 0 0.00016626 3.3 0.00016617999999999998 3.3 0.00016628 0 0.0001662 0 0.0001663 3.3 0.00016622 3.3 0.00016632 0 0.00016624 0 0.00016634 3.3 0.00016626 3.3 0.00016636 0 0.00016628 0 0.00016638 3.3 0.0001663 3.3 0.0001664 0 0.00016632 0 0.00016642 3.3 0.00016633999999999998 3.3 0.00016643999999999999 0 0.00016636 0 0.00016646 3.3 0.00016638 3.3 0.00016648 0 0.0001664 0 0.0001665 3.3 0.00016642 3.3 0.00016652 0 0.00016643999999999999 0 0.00016654 3.3 0.00016646 3.3 0.00016656 0 0.00016648 0 0.00016658 3.3 0.00016649999999999998 3.3 0.00016659999999999998 0 0.00016652 0 0.00016662 3.3 0.00016654 3.3 0.00016664 0 0.00016656 0 0.00016666 3.3 0.00016658 3.3 0.00016668 0 0.00016659999999999998 0 0.00016669999999999999 3.3 0.00016662 3.3 0.00016672 0 0.00016664 0 0.00016674 3.3 0.00016666 3.3 0.00016676 0 0.00016668 0 0.00016678 3.3 0.00016669999999999999 3.3 0.0001668 0 0.00016672 0 0.00016682 3.3 0.00016674 3.3 0.00016684 0 0.00016675999999999998 0 0.00016685999999999998 3.3 0.00016678 3.3 0.00016688 0 0.0001668 0 0.0001669 3.3 0.00016682 3.3 0.00016692 0 0.00016684 0 0.00016694 3.3 0.00016685999999999998 3.3 0.00016696 0 0.00016688 0 0.00016698 3.3 0.0001669 3.3 0.000167 0 0.00016691999999999998 0 0.00016701999999999998 3.3 0.00016694 3.3 0.00016704 0 0.00016696 0 0.00016706 3.3 0.00016698 3.3 0.00016708 0 0.000167 0 0.0001671 3.3 0.00016701999999999998 3.3 0.00016711999999999999 0 0.00016704 0 0.00016714 3.3 0.00016706 3.3 0.00016716 0 0.00016708 0 0.00016718 3.3 0.0001671 3.3 0.0001672 0 0.00016711999999999999 0 0.00016722 3.3 0.00016714 3.3 0.00016724 0 0.00016716 0 0.00016726 3.3 0.00016717999999999998 3.3 0.00016727999999999998 0 0.0001672 0 0.0001673 3.3 0.00016722 3.3 0.00016732 0 0.00016724 0 0.00016734 3.3 0.00016726 3.3 0.00016736 0 0.00016727999999999998 0 0.00016738 3.3 0.0001673 3.3 0.0001674 0 0.00016732 0 0.00016742 3.3 0.00016734 3.3 0.00016744 0 0.00016736 0 0.00016746 3.3 0.00016738 3.3 0.00016748 0 0.0001674 0 0.0001675 3.3 0.00016742 3.3 0.00016752 0 0.00016743999999999998 0 0.00016753999999999998 3.3 0.00016746 3.3 0.00016756 0 0.00016748 0 0.00016758 3.3 0.0001675 3.3 0.0001676 0 0.00016752 0 0.00016762 3.3 0.00016753999999999998 3.3 0.00016764 0 0.00016756 0 0.00016766 3.3 0.00016758 3.3 0.00016768 0 0.00016759999999999998 0 0.00016769999999999998 3.3 0.00016762 3.3 0.00016772 0 0.00016764 0 0.00016774 3.3 0.00016766 3.3 0.00016776 0 0.00016768 0 0.00016778 3.3 0.00016769999999999998 3.3 0.00016779999999999999 0 0.00016772 0 0.00016782 3.3 0.00016774 3.3 0.00016784 0 0.00016776 0 0.00016786 3.3 0.00016778 3.3 0.00016788 0 0.00016779999999999999 0 0.0001679 3.3 0.00016782 3.3 0.00016792 0 0.00016784 0 0.00016794 3.3 0.00016785999999999998 3.3 0.00016795999999999998 0 0.00016788 0 0.00016798 3.3 0.0001679 3.3 0.000168 0 0.00016792 0 0.00016802 3.3 0.00016794 3.3 0.00016804 0 0.00016795999999999998 0 0.00016806 3.3 0.00016798 3.3 0.00016808 0 0.000168 0 0.0001681 3.3 0.00016802 3.3 0.00016812 0 0.00016804 0 0.00016814 3.3 0.00016806 3.3 0.00016816 0 0.00016808 0 0.00016818 3.3 0.0001681 3.3 0.0001682 0 0.00016811999999999998 0 0.00016821999999999999 3.3 0.00016814 3.3 0.00016824 0 0.00016816 0 0.00016826 3.3 0.00016818 3.3 0.00016828 0 0.0001682 0 0.0001683 3.3 0.00016821999999999999 3.3 0.00016832 0 0.00016824 0 0.00016834 3.3 0.00016826 3.3 0.00016836 0 0.00016827999999999998 0 0.00016837999999999998 3.3 0.0001683 3.3 0.0001684 0 0.00016832 0 0.00016842 3.3 0.00016834 3.3 0.00016844 0 0.00016836 0 0.00016846 3.3 0.00016837999999999998 3.3 0.00016847999999999999 0 0.0001684 0 0.0001685 3.3 0.00016842 3.3 0.00016852 0 0.00016844 0 0.00016854 3.3 0.00016846 3.3 0.00016856 0 0.00016847999999999999 0 0.00016858 3.3 0.0001685 3.3 0.0001686 0 0.00016852 0 0.00016862 3.3 0.00016853999999999998 3.3 0.00016863999999999998 0 0.00016856 0 0.00016866 3.3 0.00016858 3.3 0.00016868 0 0.0001686 0 0.0001687 3.3 0.00016862 3.3 0.00016872 0 0.00016863999999999998 0 0.00016874 3.3 0.00016866 3.3 0.00016876 0 0.00016868 0 0.00016878 3.3 0.0001687 3.3 0.0001688 0 0.00016872 0 0.00016882 3.3 0.00016874 3.3 0.00016884 0 0.00016876 0 0.00016886 3.3 0.00016878 3.3 0.00016888 0 0.00016879999999999998 0 0.00016889999999999999 3.3 0.00016882 3.3 0.00016892 0 0.00016884 0 0.00016894 3.3 0.00016886 3.3 0.00016896 0 0.00016888 0 0.00016898 3.3 0.00016889999999999999 3.3 0.000169 0 0.00016892 0 0.00016902 3.3 0.00016894 3.3 0.00016904 0 0.00016895999999999998 0 0.00016905999999999998 3.3 0.00016898 3.3 0.00016908 0 0.000169 0 0.0001691 3.3 0.00016902 3.3 0.00016912 0 0.00016904 0 0.00016914 3.3 0.00016905999999999998 3.3 0.00016915999999999999 0 0.00016908 0 0.00016918 3.3 0.0001691 3.3 0.0001692 0 0.00016912 0 0.00016922 3.3 0.00016914 3.3 0.00016924 0 0.00016915999999999999 0 0.00016926 3.3 0.00016918 3.3 0.00016928 0 0.0001692 0 0.0001693 3.3 0.00016921999999999998 3.3 0.00016931999999999998 0 0.00016924 0 0.00016934 3.3 0.00016926 3.3 0.00016936 0 0.00016928 0 0.00016938 3.3 0.0001693 3.3 0.0001694 0 0.00016931999999999998 0 0.00016942 3.3 0.00016934 3.3 0.00016944 0 0.00016936 0 0.00016946 3.3 0.00016937999999999998 3.3 0.00016947999999999998 0 0.0001694 0 0.0001695 3.3 0.00016942 3.3 0.00016952 0 0.00016944 0 0.00016954 3.3 0.00016946 3.3 0.00016956 0 0.00016947999999999998 0 0.00016957999999999999 3.3 0.0001695 3.3 0.0001696 0 0.00016952 0 0.00016962 3.3 0.00016954 3.3 0.00016964 0 0.00016956 0 0.00016966 3.3 0.00016957999999999999 3.3 0.00016968 0 0.0001696 0 0.0001697 3.3 0.00016962 3.3 0.00016972 0 0.00016963999999999998 0 0.00016973999999999998 3.3 0.00016966 3.3 0.00016976 0 0.00016968 0 0.00016978 3.3 0.0001697 3.3 0.0001698 0 0.00016972 0 0.00016982 3.3 0.00016973999999999998 3.3 0.00016984 0 0.00016976 0 0.00016986 3.3 0.00016978 3.3 0.00016988 0 0.0001698 0 0.0001699 3.3 0.00016982 3.3 0.00016992 0 0.00016984 0 0.00016994 3.3 0.00016986 3.3 0.00016996 0 0.00016988 0 0.00016998 3.3 0.00016989999999999998 3.3 0.00016999999999999999 0 0.00016992 0 0.00017002 3.3 0.00016994 3.3 0.00017004 0 0.00016996 0 0.00017006 3.3 0.00016998 3.3 0.00017008 0 0.00016999999999999999 0 0.0001701 3.3 0.00017002 3.3 0.00017012 0 0.00017004 0 0.00017014 3.3 0.00017005999999999998 3.3 0.00017015999999999998 0 0.00017008 0 0.00017018 3.3 0.0001701 3.3 0.0001702 0 0.00017012 0 0.00017022 3.3 0.00017014 3.3 0.00017024 0 0.00017015999999999998 0 0.00017025999999999999 3.3 0.00017018 3.3 0.00017028 0 0.0001702 0 0.0001703 3.3 0.00017022 3.3 0.00017032 0 0.00017024 0 0.00017034 3.3 0.00017025999999999999 3.3 0.00017036 0 0.00017028 0 0.00017038 3.3 0.0001703 3.3 0.0001704 0 0.00017031999999999998 0 0.00017041999999999998 3.3 0.00017034 3.3 0.00017044 0 0.00017036 0 0.00017046 3.3 0.00017038 3.3 0.00017048 0 0.0001704 0 0.0001705 3.3 0.00017041999999999998 3.3 0.00017052 0 0.00017044 0 0.00017054 3.3 0.00017046 3.3 0.00017056 0 0.00017048 0 0.00017058 3.3 0.0001705 3.3 0.0001706 0 0.00017052 0 0.00017062 3.3 0.00017054 3.3 0.00017064 0 0.00017056 0 0.00017066 3.3 0.00017057999999999998 3.3 0.00017067999999999999 0 0.0001706 0 0.0001707 3.3 0.00017062 3.3 0.00017072 0 0.00017064 0 0.00017074 3.3 0.00017066 3.3 0.00017076 0 0.00017067999999999999 0 0.00017078 3.3 0.0001707 3.3 0.0001708 0 0.00017072 0 0.00017082 3.3 0.00017073999999999998 3.3 0.00017083999999999998 0 0.00017076 0 0.00017086 3.3 0.00017078 3.3 0.00017088 0 0.0001708 0 0.0001709 3.3 0.00017082 3.3 0.00017092 0 0.00017083999999999998 0 0.00017093999999999999 3.3 0.00017086 3.3 0.00017096 0 0.00017088 0 0.00017098 3.3 0.0001709 3.3 0.000171 0 0.00017092 0 0.00017102 3.3 0.00017093999999999999 3.3 0.00017104 0 0.00017096 0 0.00017106 3.3 0.00017098 3.3 0.00017108 0 0.00017099999999999998 0 0.00017109999999999998 3.3 0.00017102 3.3 0.00017112 0 0.00017104 0 0.00017114 3.3 0.00017106 3.3 0.00017116 0 0.00017108 0 0.00017118 3.3 0.00017109999999999998 3.3 0.0001712 0 0.00017112 0 0.00017122 3.3 0.00017114 3.3 0.00017124 0 0.00017115999999999998 0 0.00017125999999999998 3.3 0.00017118 3.3 0.00017128 0 0.0001712 0 0.0001713 3.3 0.00017122 3.3 0.00017132 0 0.00017124 0 0.00017134 3.3 0.00017125999999999998 3.3 0.00017135999999999999 0 0.00017128 0 0.00017138 3.3 0.0001713 3.3 0.0001714 0 0.00017132 0 0.00017142 3.3 0.00017134 3.3 0.00017144 0 0.00017135999999999999 0 0.00017146 3.3 0.00017138 3.3 0.00017148 0 0.0001714 0 0.0001715 3.3 0.00017141999999999998 3.3 0.00017151999999999998 0 0.00017144 0 0.00017154 3.3 0.00017146 3.3 0.00017156 0 0.00017148 0 0.00017158 3.3 0.0001715 3.3 0.0001716 0 0.00017151999999999998 0 0.00017162 3.3 0.00017154 3.3 0.00017164 0 0.00017156 0 0.00017166 3.3 0.00017158 3.3 0.00017168 0 0.0001716 0 0.0001717 3.3 0.00017162 3.3 0.00017172 0 0.00017164 0 0.00017174 3.3 0.00017166 3.3 0.00017176 0 0.00017167999999999998 0 0.00017177999999999999 3.3 0.0001717 3.3 0.0001718 0 0.00017172 0 0.00017182 3.3 0.00017174 3.3 0.00017184 0 0.00017176 0 0.00017186 3.3 0.00017177999999999999 3.3 0.00017188 0 0.0001718 0 0.0001719 3.3 0.00017182 3.3 0.00017192 0 0.00017183999999999998 0 0.00017193999999999998 3.3 0.00017186 3.3 0.00017196 0 0.00017188 0 0.00017198 3.3 0.0001719 3.3 0.000172 0 0.00017192 0 0.00017202 3.3 0.00017193999999999998 3.3 0.00017203999999999999 0 0.00017196 0 0.00017206 3.3 0.00017198 3.3 0.00017208 0 0.000172 0 0.0001721 3.3 0.00017202 3.3 0.00017212 0 0.00017203999999999999 0 0.00017214 3.3 0.00017206 3.3 0.00017216 0 0.00017208 0 0.00017218 3.3 0.00017209999999999998 3.3 0.00017219999999999998 0 0.00017212 0 0.00017222 3.3 0.00017214 3.3 0.00017224 0 0.00017216 0 0.00017226 3.3 0.00017218 3.3 0.00017228 0 0.00017219999999999998 0 0.0001723 3.3 0.00017222 3.3 0.00017232 0 0.00017224 0 0.00017234 3.3 0.00017226 3.3 0.00017236 0 0.00017228 0 0.00017238 3.3 0.0001723 3.3 0.0001724 0 0.00017232 0 0.00017242 3.3 0.00017234 3.3 0.00017244 0 0.00017235999999999998 0 0.00017245999999999999 3.3 0.00017238 3.3 0.00017248 0 0.0001724 0 0.0001725 3.3 0.00017242 3.3 0.00017252 0 0.00017244 0 0.00017254 3.3 0.00017245999999999999 3.3 0.00017256 0 0.00017248 0 0.00017258 3.3 0.0001725 3.3 0.0001726 0 0.00017251999999999998 0 0.00017261999999999998 3.3 0.00017254 3.3 0.00017264 0 0.00017256 0 0.00017266 3.3 0.00017258 3.3 0.00017268 0 0.0001726 0 0.0001727 3.3 0.00017261999999999998 3.3 0.00017271999999999999 0 0.00017264 0 0.00017274 3.3 0.00017266 3.3 0.00017276 0 0.00017268 0 0.00017278 3.3 0.0001727 3.3 0.0001728 0 0.00017271999999999999 0 0.00017282 3.3 0.00017274 3.3 0.00017284 0 0.00017276 0 0.00017286 3.3 0.00017277999999999998 3.3 0.00017287999999999998 0 0.0001728 0 0.0001729 3.3 0.00017282 3.3 0.00017292 0 0.00017284 0 0.00017294 3.3 0.00017286 3.3 0.00017296 0 0.00017287999999999998 0 0.00017298 3.3 0.0001729 3.3 0.000173 0 0.00017292 0 0.00017302 3.3 0.00017293999999999998 3.3 0.00017303999999999998 0 0.00017296 0 0.00017306 3.3 0.00017298 3.3 0.00017308 0 0.000173 0 0.0001731 3.3 0.00017302 3.3 0.00017312 0 0.00017303999999999998 0 0.00017313999999999999 3.3 0.00017306 3.3 0.00017316 0 0.00017308 0 0.00017318 3.3 0.0001731 3.3 0.0001732 0 0.00017312 0 0.00017322 3.3 0.00017313999999999999 3.3 0.00017324 0 0.00017316 0 0.00017326 3.3 0.00017318 3.3 0.00017328 0 0.00017319999999999998 0 0.00017329999999999998 3.3 0.00017322 3.3 0.00017332 0 0.00017324 0 0.00017334 3.3 0.00017326 3.3 0.00017336 0 0.00017328 0 0.00017338 3.3 0.00017329999999999998 3.3 0.00017339999999999999 0 0.00017332 0 0.00017342 3.3 0.00017334 3.3 0.00017344 0 0.00017336 0 0.00017346 3.3 0.00017338 3.3 0.00017348 0 0.00017339999999999999 0 0.0001735 3.3 0.00017342 3.3 0.00017352 0 0.00017344 0 0.00017354 3.3 0.00017345999999999998 3.3 0.00017355999999999998 0 0.00017348 0 0.00017358 3.3 0.0001735 3.3 0.0001736 0 0.00017352 0 0.00017362 3.3 0.00017354 3.3 0.00017364 0 0.00017355999999999998 0 0.00017366 3.3 0.00017358 3.3 0.00017368 0 0.0001736 0 0.0001737 3.3 0.00017361999999999998 3.3 0.00017371999999999998 0 0.00017364 0 0.00017374 3.3 0.00017366 3.3 0.00017376 0 0.00017368 0 0.00017378 3.3 0.0001737 3.3 0.0001738 0 0.00017371999999999998 0 0.00017381999999999999 3.3 0.00017374 3.3 0.00017384 0 0.00017376 0 0.00017386 3.3 0.00017378 3.3 0.00017388 0 0.0001738 0 0.0001739 3.3 0.00017381999999999999 3.3 0.00017392 0 0.00017384 0 0.00017394 3.3 0.00017386 3.3 0.00017396 0 0.00017387999999999998 0 0.00017397999999999998 3.3 0.0001739 3.3 0.000174 0 0.00017392 0 0.00017402 3.3 0.00017394 3.3 0.00017404 0 0.00017396 0 0.00017406 3.3 0.00017397999999999998 3.3 0.00017408 0 0.000174 0 0.0001741 3.3 0.00017402 3.3 0.00017412 0 0.00017404 0 0.00017414 3.3 0.00017406 3.3 0.00017416 0 0.00017408 0 0.00017418 3.3 0.0001741 3.3 0.0001742 0 0.00017412 0 0.00017422 3.3 0.00017413999999999998 3.3 0.00017423999999999999 0 0.00017416 0 0.00017426 3.3 0.00017418 3.3 0.00017428 0 0.0001742 0 0.0001743 3.3 0.00017422 3.3 0.00017432 0 0.00017423999999999999 0 0.00017434 3.3 0.00017426 3.3 0.00017436 0 0.00017428 0 0.00017438 3.3 0.00017429999999999998 3.3 0.00017439999999999998 0 0.00017432 0 0.00017442 3.3 0.00017434 3.3 0.00017444 0 0.00017436 0 0.00017446 3.3 0.00017438 3.3 0.00017448 0 0.00017439999999999998 0 0.00017449999999999999 3.3 0.00017442 3.3 0.00017452 0 0.00017444 0 0.00017454 3.3 0.00017446 3.3 0.00017456 0 0.00017448 0 0.00017458 3.3 0.00017449999999999999 3.3 0.0001746 0 0.00017452 0 0.00017462 3.3 0.00017454 3.3 0.00017464 0 0.00017455999999999998 0 0.00017465999999999998 3.3 0.00017458 3.3 0.00017468 0 0.0001746 0 0.0001747 3.3 0.00017462 3.3 0.00017472 0 0.00017464 0 0.00017474 3.3 0.00017465999999999998 3.3 0.00017476 0 0.00017468 0 0.00017478 3.3 0.0001747 3.3 0.0001748 0 0.00017471999999999998 0 0.00017481999999999998 3.3 0.00017474 3.3 0.00017484 0 0.00017476 0 0.00017486 3.3 0.00017478 3.3 0.00017488 0 0.0001748 0 0.0001749 3.3 0.00017481999999999998 3.3 0.00017491999999999999 0 0.00017484 0 0.00017494 3.3 0.00017486 3.3 0.00017496 0 0.00017488 0 0.00017498 3.3 0.0001749 3.3 0.000175 0 0.00017491999999999999 0 0.00017502 3.3 0.00017494 3.3 0.00017504 0 0.00017496 0 0.00017506 3.3 0.00017497999999999998 3.3 0.00017507999999999998 0 0.000175 0 0.0001751 3.3 0.00017502 3.3 0.00017512 0 0.00017504 0 0.00017514 3.3 0.00017506 3.3 0.00017516 0 0.00017507999999999998 0 0.00017517999999999999 3.3 0.0001751 3.3 0.0001752 0 0.00017512 0 0.00017522 3.3 0.00017514 3.3 0.00017524 0 0.00017516 0 0.00017526 3.3 0.00017517999999999999 3.3 0.00017528 0 0.0001752 0 0.0001753 3.3 0.00017522 3.3 0.00017532 0 0.00017523999999999998 0 0.00017533999999999998 3.3 0.00017526 3.3 0.00017536 0 0.00017528 0 0.00017538 3.3 0.0001753 3.3 0.0001754 0 0.00017532 0 0.00017542 3.3 0.00017533999999999998 3.3 0.00017544 0 0.00017536 0 0.00017546 3.3 0.00017538 3.3 0.00017548 0 0.00017539999999999998 0 0.00017549999999999998 3.3 0.00017542 3.3 0.00017552 0 0.00017544 0 0.00017554 3.3 0.00017546 3.3 0.00017556 0 0.00017548 0 0.00017558 3.3 0.00017549999999999998 3.3 0.00017559999999999999 0 0.00017552 0 0.00017562 3.3 0.00017554 3.3 0.00017564 0 0.00017556 0 0.00017566 3.3 0.00017558 3.3 0.00017568 0 0.00017559999999999999 0 0.0001757 3.3 0.00017562 3.3 0.00017572 0 0.00017564 0 0.00017574 3.3 0.00017565999999999998 3.3 0.00017575999999999998 0 0.00017568 0 0.00017578 3.3 0.0001757 3.3 0.0001758 0 0.00017572 0 0.00017582 3.3 0.00017574 3.3 0.00017584 0 0.00017575999999999998 0 0.00017586 3.3 0.00017578 3.3 0.00017588 0 0.0001758 0 0.0001759 3.3 0.00017582 3.3 0.00017592 0 0.00017584 0 0.00017594 3.3 0.00017586 3.3 0.00017596 0 0.00017588 0 0.00017598 3.3 0.0001759 3.3 0.000176 0 0.00017591999999999998 0 0.00017601999999999999 3.3 0.00017594 3.3 0.00017604 0 0.00017596 0 0.00017606 3.3 0.00017598 3.3 0.00017608 0 0.000176 0 0.0001761 3.3 0.00017601999999999999 3.3 0.00017612 0 0.00017604 0 0.00017614 3.3 0.00017606 3.3 0.00017616 0 0.00017607999999999998 0 0.00017617999999999998 3.3 0.0001761 3.3 0.0001762 0 0.00017612 0 0.00017622 3.3 0.00017614 3.3 0.00017624 0 0.00017616 0 0.00017626 3.3 0.00017617999999999998 3.3 0.00017627999999999999 0 0.0001762 0 0.0001763 3.3 0.00017622 3.3 0.00017632 0 0.00017624 0 0.00017634 3.3 0.00017626 3.3 0.00017636 0 0.00017627999999999999 0 0.00017638 3.3 0.0001763 3.3 0.0001764 0 0.00017632 0 0.00017642 3.3 0.00017633999999999998 3.3 0.00017643999999999998 0 0.00017636 0 0.00017646 3.3 0.00017638 3.3 0.00017648 0 0.0001764 0 0.0001765 3.3 0.00017642 3.3 0.00017652 0 0.00017643999999999998 0 0.00017654 3.3 0.00017646 3.3 0.00017656 0 0.00017648 0 0.00017658 3.3 0.00017649999999999998 3.3 0.00017659999999999998 0 0.00017652 0 0.00017662 3.3 0.00017654 3.3 0.00017664 0 0.00017656 0 0.00017666 3.3 0.00017658 3.3 0.00017668 0 0.00017659999999999998 0 0.00017669999999999999 3.3 0.00017662 3.3 0.00017672 0 0.00017664 0 0.00017674 3.3 0.00017666 3.3 0.00017676 0 0.00017668 0 0.00017678 3.3 0.00017669999999999999 3.3 0.0001768 0 0.00017672 0 0.00017682 3.3 0.00017674 3.3 0.00017684 0 0.00017675999999999998 0 0.00017685999999999998 3.3 0.00017678 3.3 0.00017688 0 0.0001768 0 0.0001769 3.3 0.00017682 3.3 0.00017692 0 0.00017684 0 0.00017694 3.3 0.00017685999999999998 3.3 0.00017695999999999999 0 0.00017688 0 0.00017698 3.3 0.0001769 3.3 0.000177 0 0.00017692 0 0.00017702 3.3 0.00017694 3.3 0.00017704 0 0.00017695999999999999 0 0.00017706 3.3 0.00017698 3.3 0.00017708 0 0.000177 0 0.0001771 3.3 0.00017701999999999998 3.3 0.00017711999999999998 0 0.00017704 0 0.00017714 3.3 0.00017706 3.3 0.00017716 0 0.00017708 0 0.00017718 3.3 0.0001771 3.3 0.0001772 0 0.00017711999999999998 0 0.00017722 3.3 0.00017714 3.3 0.00017724 0 0.00017716 0 0.00017726 3.3 0.00017717999999999998 3.3 0.00017727999999999998 0 0.0001772 0 0.0001773 3.3 0.00017722 3.3 0.00017732 0 0.00017724 0 0.00017734 3.3 0.00017726 3.3 0.00017736 0 0.00017727999999999998 0 0.00017737999999999999 3.3 0.0001773 3.3 0.0001774 0 0.00017732 0 0.00017742 3.3 0.00017734 3.3 0.00017744 0 0.00017736 0 0.00017746 3.3 0.00017737999999999999 3.3 0.00017748 0 0.0001774 0 0.0001775 3.3 0.00017742 3.3 0.00017752 0 0.00017743999999999998 0 0.00017753999999999998 3.3 0.00017746 3.3 0.00017756 0 0.00017748 0 0.00017758 3.3 0.0001775 3.3 0.0001776 0 0.00017752 0 0.00017762 3.3 0.00017753999999999998 3.3 0.00017764 0 0.00017756 0 0.00017766 3.3 0.00017758 3.3 0.00017768 0 0.0001776 0 0.0001777 3.3 0.00017762 3.3 0.00017772 0 0.00017764 0 0.00017774 3.3 0.00017766 3.3 0.00017776 0 0.00017768 0 0.00017778 3.3 0.00017769999999999998 3.3 0.00017779999999999998 0 0.00017772 0 0.00017782 3.3 0.00017774 3.3 0.00017784 0 0.00017776 0 0.00017786 3.3 0.00017778 3.3 0.00017788 0 0.00017779999999999998 0 0.0001779 3.3 0.00017782 3.3 0.00017792 0 0.00017784 0 0.00017794 3.3 0.00017785999999999998 3.3 0.00017795999999999998 0 0.00017788 0 0.00017798 3.3 0.0001779 3.3 0.000178 0 0.00017792 0 0.00017802 3.3 0.00017794 3.3 0.00017804 0 0.00017795999999999998 0 0.00017805999999999999 3.3 0.00017798 3.3 0.00017808 0 0.000178 0 0.0001781 3.3 0.00017802 3.3 0.00017812 0 0.00017804 0 0.00017814 3.3 0.00017805999999999999 3.3 0.00017816 0 0.00017808 0 0.00017818 3.3 0.0001781 3.3 0.0001782 0 0.00017811999999999998 0 0.00017821999999999998 3.3 0.00017814 3.3 0.00017824 0 0.00017816 0 0.00017826 3.3 0.00017818 3.3 0.00017828 0 0.0001782 0 0.0001783 3.3 0.00017821999999999998 3.3 0.00017832 0 0.00017824 0 0.00017834 3.3 0.00017826 3.3 0.00017836 0 0.00017828 0 0.00017838 3.3 0.0001783 3.3 0.0001784 0 0.00017832 0 0.00017842 3.3 0.00017834 3.3 0.00017844 0 0.00017836 0 0.00017846 3.3 0.00017837999999999998 3.3 0.00017847999999999999 0 0.0001784 0 0.0001785 3.3 0.00017842 3.3 0.00017852 0 0.00017844 0 0.00017854 3.3 0.00017846 3.3 0.00017856 0 0.00017847999999999999 0 0.00017858 3.3 0.0001785 3.3 0.0001786 0 0.00017852 0 0.00017862 3.3 0.00017853999999999998 3.3 0.00017863999999999998 0 0.00017856 0 0.00017866 3.3 0.00017858 3.3 0.00017868 0 0.0001786 0 0.0001787 3.3 0.00017862 3.3 0.00017872 0 0.00017863999999999998 0 0.00017873999999999999 3.3 0.00017866 3.3 0.00017876 0 0.00017868 0 0.00017878 3.3 0.0001787 3.3 0.0001788 0 0.00017872 0 0.00017882 3.3 0.00017873999999999999 3.3 0.00017884 0 0.00017876 0 0.00017886 3.3 0.00017878 3.3 0.00017888 0 0.00017879999999999998 0 0.00017889999999999998 3.3 0.00017882 3.3 0.00017892 0 0.00017884 0 0.00017894 3.3 0.00017886 3.3 0.00017896 0 0.00017888 0 0.00017898 3.3 0.00017889999999999998 3.3 0.000179 0 0.00017892 0 0.00017902 3.3 0.00017894 3.3 0.00017904 0 0.00017895999999999998 0 0.00017905999999999998 3.3 0.00017898 3.3 0.00017908 0 0.000179 0 0.0001791 3.3 0.00017902 3.3 0.00017912 0 0.00017904 0 0.00017914 3.3 0.00017905999999999998 3.3 0.00017915999999999999 0 0.00017908 0 0.00017918 3.3 0.0001791 3.3 0.0001792 0 0.00017912 0 0.00017922 3.3 0.00017914 3.3 0.00017924 0 0.00017915999999999999 0 0.00017926 3.3 0.00017918 3.3 0.00017928 0 0.0001792 0 0.0001793 3.3 0.00017921999999999998 3.3 0.00017931999999999998 0 0.00017924 0 0.00017934 3.3 0.00017926 3.3 0.00017936 0 0.00017928 0 0.00017938 3.3 0.0001793 3.3 0.0001794 0 0.00017931999999999998 0 0.00017941999999999999 3.3 0.00017934 3.3 0.00017944 0 0.00017936 0 0.00017946 3.3 0.00017938 3.3 0.00017948 0 0.0001794 0 0.0001795 3.3 0.00017941999999999999 3.3 0.00017952 0 0.00017944 0 0.00017954 3.3 0.00017946 3.3 0.00017956 0 0.00017947999999999998 0 0.00017957999999999998 3.3 0.0001795 3.3 0.0001796 0 0.00017952 0 0.00017962 3.3 0.00017954 3.3 0.00017964 0 0.00017956 0 0.00017966 3.3 0.00017957999999999998 3.3 0.00017968 0 0.0001796 0 0.0001797 3.3 0.00017962 3.3 0.00017972 0 0.00017963999999999998 0 0.00017973999999999998 3.3 0.00017966 3.3 0.00017976 0 0.00017968 0 0.00017978 3.3 0.0001797 3.3 0.0001798 0 0.00017972 0 0.00017982 3.3 0.00017973999999999998 3.3 0.00017983999999999999 0 0.00017976 0 0.00017986 3.3 0.00017978 3.3 0.00017988 0 0.0001798 0 0.0001799 3.3 0.00017982 3.3 0.00017992 0 0.00017983999999999999 0 0.00017994 3.3 0.00017986 3.3 0.00017996 0 0.00017988 0 0.00017998 3.3 0.00017989999999999998 3.3 0.00017999999999999998 0 0.00017992 0 0.00018002 3.3 0.00017994 3.3 0.00018004 0 0.00017996 0 0.00018006 3.3 0.00017998 3.3 0.00018008 0 0.00017999999999999998 0 0.0001801 3.3 0.00018002 3.3 0.00018012 0 0.00018004 0 0.00018014 3.3 0.00018006 3.3 0.00018016 0 0.00018008 0 0.00018018 3.3 0.0001801 3.3 0.0001802 0 0.00018012 0 0.00018022 3.3 0.00018014 3.3 0.00018024 0 0.00018015999999999998 0 0.00018025999999999999 3.3 0.00018018 3.3 0.00018028 0 0.0001802 0 0.0001803 3.3 0.00018022 3.3 0.00018032 0 0.00018024 0 0.00018034 3.3 0.00018025999999999999 3.3 0.00018036 0 0.00018028 0 0.00018038 3.3 0.0001803 3.3 0.0001804 0 0.00018031999999999998 0 0.00018041999999999998 3.3 0.00018034 3.3 0.00018044 0 0.00018036 0 0.00018046 3.3 0.00018038 3.3 0.00018048 0 0.0001804 0 0.0001805 3.3 0.00018041999999999998 3.3 0.00018051999999999999 0 0.00018044 0 0.00018054 3.3 0.00018046 3.3 0.00018056 0 0.00018048 0 0.00018058 3.3 0.0001805 3.3 0.0001806 0 0.00018051999999999999 0 0.00018062 3.3 0.00018054 3.3 0.00018064 0 0.00018056 0 0.00018066 3.3 0.00018057999999999998 3.3 0.00018067999999999998 0 0.0001806 0 0.0001807 3.3 0.00018062 3.3 0.00018072 0 0.00018064 0 0.00018074 3.3 0.00018066 3.3 0.00018076 0 0.00018067999999999998 0 0.00018078 3.3 0.0001807 3.3 0.0001808 0 0.00018072 0 0.00018082 3.3 0.00018073999999999998 3.3 0.00018083999999999998 0 0.00018076 0 0.00018086 3.3 0.00018078 3.3 0.00018088 0 0.0001808 0 0.0001809 3.3 0.00018082 3.3 0.00018092 0 0.00018083999999999998 0 0.00018093999999999999 3.3 0.00018086 3.3 0.00018096 0 0.00018088 0 0.00018098 3.3 0.0001809 3.3 0.000181 0 0.00018092 0 0.00018102 3.3 0.00018093999999999999 3.3 0.00018104 0 0.00018096 0 0.00018106 3.3 0.00018098 3.3 0.00018108 0 0.00018099999999999998 0 0.00018109999999999998 3.3 0.00018102 3.3 0.00018112 0 0.00018104 0 0.00018114 3.3 0.00018106 3.3 0.00018116 0 0.00018108 0 0.00018118 3.3 0.00018109999999999998 3.3 0.00018119999999999999 0 0.00018112 0 0.00018122 3.3 0.00018114 3.3 0.00018124 0 0.00018116 0 0.00018126 3.3 0.00018118 3.3 0.00018128 0 0.00018119999999999999 0 0.0001813 3.3 0.00018122 3.3 0.00018132 0 0.00018124 0 0.00018134 3.3 0.00018125999999999998 3.3 0.00018135999999999998 0 0.00018128 0 0.00018138 3.3 0.0001813 3.3 0.0001814 0 0.00018132 0 0.00018142 3.3 0.00018134 3.3 0.00018144 0 0.00018135999999999998 0 0.00018146 3.3 0.00018138 3.3 0.00018148 0 0.0001814 0 0.0001815 3.3 0.00018141999999999998 3.3 0.00018151999999999998 0 0.00018144 0 0.00018154 3.3 0.00018146 3.3 0.00018156 0 0.00018148 0 0.00018158 3.3 0.0001815 3.3 0.0001816 0 0.00018151999999999998 0 0.00018161999999999999 3.3 0.00018154 3.3 0.00018164 0 0.00018156 0 0.00018166 3.3 0.00018158 3.3 0.00018168 0 0.0001816 0 0.0001817 3.3 0.00018161999999999999 3.3 0.00018172 0 0.00018164 0 0.00018174 3.3 0.00018166 3.3 0.00018176 0 0.00018167999999999998 0 0.00018177999999999998 3.3 0.0001817 3.3 0.0001818 0 0.00018172 0 0.00018182 3.3 0.00018174 3.3 0.00018184 0 0.00018176 0 0.00018186 3.3 0.00018177999999999998 3.3 0.00018188 0 0.0001818 0 0.0001819 3.3 0.00018182 3.3 0.00018192 0 0.00018184 0 0.00018194 3.3 0.00018186 3.3 0.00018196 0 0.00018188 0 0.00018198 3.3 0.0001819 3.3 0.000182 0 0.00018192 0 0.00018202 3.3 0.00018193999999999998 3.3 0.00018203999999999999 0 0.00018196 0 0.00018206 3.3 0.00018198 3.3 0.00018208 0 0.000182 0 0.0001821 3.3 0.00018202 3.3 0.00018212 0 0.00018203999999999999 0 0.00018214 3.3 0.00018206 3.3 0.00018216 0 0.00018208 0 0.00018218 3.3 0.00018209999999999998 3.3 0.00018219999999999998 0 0.00018212 0 0.00018222 3.3 0.00018214 3.3 0.00018224 0 0.00018216 0 0.00018226 3.3 0.00018218 3.3 0.00018228 0 0.00018219999999999998 0 0.00018229999999999999 3.3 0.00018222 3.3 0.00018232 0 0.00018224 0 0.00018234 3.3 0.00018226 3.3 0.00018236 0 0.00018228 0 0.00018238 3.3 0.00018229999999999999 3.3 0.0001824 0 0.00018232 0 0.00018242 3.3 0.00018234 3.3 0.00018244 0 0.00018235999999999998 0 0.00018245999999999998 3.3 0.00018238 3.3 0.00018248 0 0.0001824 0 0.0001825 3.3 0.00018242 3.3 0.00018252 0 0.00018244 0 0.00018254 3.3 0.00018245999999999998 3.3 0.00018256 0 0.00018248 0 0.00018258 3.3 0.0001825 3.3 0.0001826 0 0.00018251999999999998 0 0.00018261999999999998 3.3 0.00018254 3.3 0.00018264 0 0.00018256 0 0.00018266 3.3 0.00018258 3.3 0.00018268 0 0.0001826 0 0.0001827 3.3 0.00018261999999999998 3.3 0.00018271999999999999 0 0.00018264 0 0.00018274 3.3 0.00018266 3.3 0.00018276 0 0.00018268 0 0.00018278 3.3 0.0001827 3.3 0.0001828 0 0.00018271999999999999 0 0.00018282 3.3 0.00018274 3.3 0.00018284 0 0.00018276 0 0.00018286 3.3 0.00018277999999999998 3.3 0.00018287999999999998 0 0.0001828 0 0.0001829 3.3 0.00018282 3.3 0.00018292 0 0.00018284 0 0.00018294 3.3 0.00018286 3.3 0.00018296 0 0.00018287999999999998 0 0.00018297999999999999 3.3 0.0001829 3.3 0.000183 0 0.00018292 0 0.00018302 3.3 0.00018294 3.3 0.00018304 0 0.00018296 0 0.00018306 3.3 0.00018297999999999999 3.3 0.00018308 0 0.000183 0 0.0001831 3.3 0.00018302 3.3 0.00018312 0 0.00018303999999999998 0 0.00018313999999999998 3.3 0.00018306 3.3 0.00018316 0 0.00018308 0 0.00018318 3.3 0.0001831 3.3 0.0001832 0 0.00018312 0 0.00018322 3.3 0.00018313999999999998 3.3 0.00018324 0 0.00018316 0 0.00018326 3.3 0.00018318 3.3 0.00018328 0 0.00018319999999999998 0 0.00018329999999999998 3.3 0.00018322 3.3 0.00018332 0 0.00018324 0 0.00018334 3.3 0.00018326 3.3 0.00018336 0 0.00018328 0 0.00018338 3.3 0.00018329999999999998 3.3 0.00018339999999999999 0 0.00018332 0 0.00018342 3.3 0.00018334 3.3 0.00018344 0 0.00018336 0 0.00018346 3.3 0.00018338 3.3 0.00018348 0 0.00018339999999999999 0 0.0001835 3.3 0.00018342 3.3 0.00018352 0 0.00018344 0 0.00018354 3.3 0.00018345999999999998 3.3 0.00018355999999999998 0 0.00018348 0 0.00018358 3.3 0.0001835 3.3 0.0001836 0 0.00018352 0 0.00018362 3.3 0.00018354 3.3 0.00018364 0 0.00018355999999999998 0 0.00018366 3.3 0.00018358 3.3 0.00018368 0 0.0001836 0 0.0001837 3.3 0.00018362 3.3 0.00018372 0 0.00018364 0 0.00018374 3.3 0.00018366 3.3 0.00018376 0 0.00018368 0 0.00018378 3.3 0.0001837 3.3 0.0001838 0 0.00018371999999999998 0 0.00018381999999999998 3.3 0.00018374 3.3 0.00018384 0 0.00018376 0 0.00018386 3.3 0.00018378 3.3 0.00018388 0 0.0001838 0 0.0001839 3.3 0.00018381999999999998 3.3 0.00018392 0 0.00018384 0 0.00018394 3.3 0.00018386 3.3 0.00018396 0 0.00018387999999999998 0 0.00018397999999999998 3.3 0.0001839 3.3 0.000184 0 0.00018392 0 0.00018402 3.3 0.00018394 3.3 0.00018404 0 0.00018396 0 0.00018406 3.3 0.00018397999999999998 3.3 0.00018407999999999999 0 0.000184 0 0.0001841 3.3 0.00018402 3.3 0.00018412 0 0.00018404 0 0.00018414 3.3 0.00018406 3.3 0.00018416 0 0.00018407999999999999 0 0.00018418 3.3 0.0001841 3.3 0.0001842 0 0.00018412 0 0.00018422 3.3 0.00018413999999999998 3.3 0.00018423999999999998 0 0.00018416 0 0.00018426 3.3 0.00018418 3.3 0.00018428 0 0.0001842 0 0.0001843 3.3 0.00018422 3.3 0.00018432 0 0.00018423999999999998 0 0.00018434 3.3 0.00018426 3.3 0.00018436 0 0.00018428 0 0.00018438 3.3 0.00018429999999999998 3.3 0.00018439999999999998 0 0.00018432 0 0.00018442 3.3 0.00018434 3.3 0.00018444 0 0.00018436 0 0.00018446 3.3 0.00018438 3.3 0.00018448 0 0.00018439999999999998 0 0.00018449999999999999 3.3 0.00018442 3.3 0.00018452 0 0.00018444 0 0.00018454 3.3 0.00018446 3.3 0.00018456 0 0.00018448 0 0.00018458 3.3 0.00018449999999999999 3.3 0.0001846 0 0.00018452 0 0.00018462 3.3 0.00018454 3.3 0.00018464 0 0.00018455999999999998 0 0.00018465999999999998 3.3 0.00018458 3.3 0.00018468 0 0.0001846 0 0.0001847 3.3 0.00018462 3.3 0.00018472 0 0.00018464 0 0.00018474 3.3 0.00018465999999999998 3.3 0.00018475999999999999 0 0.00018468 0 0.00018478 3.3 0.0001847 3.3 0.0001848 0 0.00018472 0 0.00018482 3.3 0.00018474 3.3 0.00018484 0 0.00018475999999999999 0 0.00018486 3.3 0.00018478 3.3 0.00018488 0 0.0001848 0 0.0001849 3.3 0.00018481999999999998 3.3 0.00018491999999999998 0 0.00018484 0 0.00018494 3.3 0.00018486 3.3 0.00018496 0 0.00018488 0 0.00018498 3.3 0.0001849 3.3 0.000185 0 0.00018491999999999998 0 0.00018502 3.3 0.00018494 3.3 0.00018504 0 0.00018496 0 0.00018506 3.3 0.00018497999999999998 3.3 0.00018507999999999998 0 0.000185 0 0.0001851 3.3 0.00018502 3.3 0.00018512 0 0.00018504 0 0.00018514 3.3 0.00018506 3.3 0.00018516 0 0.00018507999999999998 0 0.00018517999999999999 3.3 0.0001851 3.3 0.0001852 0 0.00018512 0 0.00018522 3.3 0.00018514 3.3 0.00018524 0 0.00018516 0 0.00018526 3.3 0.00018517999999999999 3.3 0.00018528 0 0.0001852 0 0.0001853 3.3 0.00018522 3.3 0.00018532 0 0.00018523999999999998 0 0.00018533999999999998 3.3 0.00018526 3.3 0.00018536 0 0.00018528 0 0.00018538 3.3 0.0001853 3.3 0.0001854 0 0.00018532 0 0.00018542 3.3 0.00018533999999999998 3.3 0.00018543999999999999 0 0.00018536 0 0.00018546 3.3 0.00018538 3.3 0.00018548 0 0.0001854 0 0.0001855 3.3 0.00018542 3.3 0.00018552 0 0.00018543999999999999 0 0.00018554 3.3 0.00018546 3.3 0.00018556 0 0.00018548 0 0.00018558 3.3 0.00018549999999999998 3.3 0.00018559999999999998 0 0.00018552 0 0.00018562 3.3 0.00018554 3.3 0.00018564 0 0.00018556 0 0.00018566 3.3 0.00018558 3.3 0.00018568 0 0.00018559999999999998 0 0.0001857 3.3 0.00018562 3.3 0.00018572 0 0.00018564 0 0.00018574 3.3 0.00018565999999999998 3.3 0.00018575999999999998 0 0.00018568 0 0.00018578 3.3 0.0001857 3.3 0.0001858 0 0.00018572 0 0.00018582 3.3 0.00018574 3.3 0.00018584 0 0.00018575999999999998 0 0.00018585999999999999 3.3 0.00018578 3.3 0.00018588 0 0.0001858 0 0.0001859 3.3 0.00018582 3.3 0.00018592 0 0.00018584 0 0.00018594 3.3 0.00018585999999999999 3.3 0.00018596 0 0.00018588 0 0.00018598 3.3 0.0001859 3.3 0.000186 0 0.00018591999999999998 0 0.00018601999999999998 3.3 0.00018594 3.3 0.00018604 0 0.00018596 0 0.00018606 3.3 0.00018598 3.3 0.00018608 0 0.000186 0 0.0001861 3.3 0.00018601999999999998 3.3 0.00018612 0 0.00018604 0 0.00018614 3.3 0.00018606 3.3 0.00018616 0 0.00018608 0 0.00018618 3.3 0.0001861 3.3 0.0001862 0 0.00018612 0 0.00018622 3.3 0.00018614 3.3 0.00018624 0 0.00018616 0 0.00018626 3.3 0.00018617999999999998 3.3 0.00018627999999999999 0 0.0001862 0 0.0001863 3.3 0.00018622 3.3 0.00018632 0 0.00018624 0 0.00018634 3.3 0.00018626 3.3 0.00018636 0 0.00018627999999999999 0 0.00018638 3.3 0.0001863 3.3 0.0001864 0 0.00018632 0 0.00018642 3.3 0.00018633999999999998 3.3 0.00018643999999999998 0 0.00018636 0 0.00018646 3.3 0.00018638 3.3 0.00018648 0 0.0001864 0 0.0001865 3.3 0.00018642 3.3 0.00018652 0 0.00018643999999999998 0 0.00018653999999999999 3.3 0.00018646 3.3 0.00018656 0 0.00018648 0 0.00018658 3.3 0.0001865 3.3 0.0001866 0 0.00018652 0 0.00018662 3.3 0.00018653999999999999 3.3 0.00018664 0 0.00018656 0 0.00018666 3.3 0.00018658 3.3 0.00018668 0 0.00018659999999999998 0 0.00018669999999999998 3.3 0.00018662 3.3 0.00018672 0 0.00018664 0 0.00018674 3.3 0.00018666 3.3 0.00018676 0 0.00018668 0 0.00018678 3.3 0.00018669999999999998 3.3 0.0001868 0 0.00018672 0 0.00018682 3.3 0.00018674 3.3 0.00018684 0 0.00018675999999999998 0 0.00018685999999999998 3.3 0.00018678 3.3 0.00018688 0 0.0001868 0 0.0001869 3.3 0.00018682 3.3 0.00018692 0 0.00018684 0 0.00018694 3.3 0.00018685999999999998 3.3 0.00018695999999999999 0 0.00018688 0 0.00018698 3.3 0.0001869 3.3 0.000187 0 0.00018692 0 0.00018702 3.3 0.00018694 3.3 0.00018704 0 0.00018695999999999999 0 0.00018706 3.3 0.00018698 3.3 0.00018708 0 0.000187 0 0.0001871 3.3 0.00018701999999999998 3.3 0.00018711999999999998 0 0.00018704 0 0.00018714 3.3 0.00018706 3.3 0.00018716 0 0.00018708 0 0.00018718 3.3 0.0001871 3.3 0.0001872 0 0.00018711999999999998 0 0.00018721999999999999 3.3 0.00018714 3.3 0.00018724 0 0.00018716 0 0.00018726 3.3 0.00018718 3.3 0.00018728 0 0.0001872 0 0.0001873 3.3 0.00018721999999999999 3.3 0.00018732 0 0.00018724 0 0.00018734 3.3 0.00018726 3.3 0.00018736 0 0.00018727999999999998 0 0.00018737999999999998 3.3 0.0001873 3.3 0.0001874 0 0.00018732 0 0.00018742 3.3 0.00018734 3.3 0.00018744 0 0.00018736 0 0.00018746 3.3 0.00018737999999999998 3.3 0.00018748 0 0.0001874 0 0.0001875 3.3 0.00018742 3.3 0.00018752 0 0.00018743999999999998 0 0.00018753999999999998 3.3 0.00018746 3.3 0.00018756 0 0.00018748 0 0.00018758 3.3 0.0001875 3.3 0.0001876 0 0.00018752 0 0.00018762 3.3 0.00018753999999999998 3.3 0.00018763999999999999 0 0.00018756 0 0.00018766 3.3 0.00018758 3.3 0.00018768 0 0.0001876 0 0.0001877 3.3 0.00018762 3.3 0.00018772 0 0.00018763999999999999 0 0.00018774 3.3 0.00018766 3.3 0.00018776 0 0.00018768 0 0.00018778 3.3 0.00018769999999999998 3.3 0.00018779999999999998 0 0.00018772 0 0.00018782 3.3 0.00018774 3.3 0.00018784 0 0.00018776 0 0.00018786 3.3 0.00018778 3.3 0.00018788 0 0.00018779999999999998 0 0.0001879 3.3 0.00018782 3.3 0.00018792 0 0.00018784 0 0.00018794 3.3 0.00018786 3.3 0.00018796 0 0.00018788 0 0.00018798 3.3 0.0001879 3.3 0.000188 0 0.00018792 0 0.00018802 3.3 0.00018794 3.3 0.00018804 0 0.00018795999999999998 0 0.00018805999999999998 3.3 0.00018798 3.3 0.00018808 0 0.000188 0 0.0001881 3.3 0.00018802 3.3 0.00018812 0 0.00018804 0 0.00018814 3.3 0.00018805999999999998 3.3 0.00018816 0 0.00018808 0 0.00018818 3.3 0.0001881 3.3 0.0001882 0 0.00018811999999999998 0 0.00018821999999999998 3.3 0.00018814 3.3 0.00018824 0 0.00018816 0 0.00018826 3.3 0.00018818 3.3 0.00018828 0 0.0001882 0 0.0001883 3.3 0.00018821999999999998 3.3 0.00018831999999999999 0 0.00018824 0 0.00018834 3.3 0.00018826 3.3 0.00018836 0 0.00018828 0 0.00018838 3.3 0.0001883 3.3 0.0001884 0 0.00018831999999999999 0 0.00018842 3.3 0.00018834 3.3 0.00018844 0 0.00018836 0 0.00018846 3.3 0.00018837999999999998 3.3 0.00018847999999999998 0 0.0001884 0 0.0001885 3.3 0.00018842 3.3 0.00018852 0 0.00018844 0 0.00018854 3.3 0.00018846 3.3 0.00018856 0 0.00018847999999999998 0 0.00018858 3.3 0.0001885 3.3 0.0001886 0 0.00018852 0 0.00018862 3.3 0.00018853999999999998 3.3 0.00018863999999999998 0 0.00018856 0 0.00018866 3.3 0.00018858 3.3 0.00018868 0 0.0001886 0 0.0001887 3.3 0.00018862 3.3 0.00018872 0 0.00018863999999999998 0 0.00018873999999999999 3.3 0.00018866 3.3 0.00018876 0 0.00018868 0 0.00018878 3.3 0.0001887 3.3 0.0001888 0 0.00018872 0 0.00018882 3.3 0.00018873999999999999 3.3 0.00018884 0 0.00018876 0 0.00018886 3.3 0.00018878 3.3 0.00018888 0 0.00018879999999999998 0 0.00018889999999999998 3.3 0.00018882 3.3 0.00018892 0 0.00018884 0 0.00018894 3.3 0.00018886 3.3 0.00018896 0 0.00018888 0 0.00018898 3.3 0.00018889999999999998 3.3 0.00018899999999999999 0 0.00018892 0 0.00018902 3.3 0.00018894 3.3 0.00018904 0 0.00018896 0 0.00018906 3.3 0.00018898 3.3 0.00018908 0 0.00018899999999999999 0 0.0001891 3.3 0.00018902 3.3 0.00018912 0 0.00018904 0 0.00018914 3.3 0.00018905999999999998 3.3 0.00018915999999999998 0 0.00018908 0 0.00018918 3.3 0.0001891 3.3 0.0001892 0 0.00018912 0 0.00018922 3.3 0.00018914 3.3 0.00018924 0 0.00018915999999999998 0 0.00018926 3.3 0.00018918 3.3 0.00018928 0 0.0001892 0 0.0001893 3.3 0.00018921999999999998 3.3 0.00018931999999999998 0 0.00018924 0 0.00018934 3.3 0.00018926 3.3 0.00018936 0 0.00018928 0 0.00018938 3.3 0.0001893 3.3 0.0001894 0 0.00018931999999999998 0 0.00018941999999999999 3.3 0.00018934 3.3 0.00018944 0 0.00018936 0 0.00018946 3.3 0.00018938 3.3 0.00018948 0 0.0001894 0 0.0001895 3.3 0.00018941999999999999 3.3 0.00018952 0 0.00018944 0 0.00018954 3.3 0.00018946 3.3 0.00018956 0 0.00018947999999999998 0 0.00018957999999999998 3.3 0.0001895 3.3 0.0001896 0 0.00018952 0 0.00018962 3.3 0.00018954 3.3 0.00018964 0 0.00018956 0 0.00018966 3.3 0.00018957999999999998 3.3 0.00018967999999999999 0 0.0001896 0 0.0001897 3.3 0.00018962 3.3 0.00018972 0 0.00018964 0 0.00018974 3.3 0.00018966 3.3 0.00018976 0 0.00018967999999999999 0 0.00018978 3.3 0.0001897 3.3 0.0001898 0 0.00018972 0 0.00018982 3.3 0.00018973999999999998 3.3 0.00018983999999999998 0 0.00018976 0 0.00018986 3.3 0.00018978 3.3 0.00018988 0 0.0001898 0 0.0001899 3.3 0.00018982 3.3 0.00018992 0 0.00018983999999999998 0 0.00018994 3.3 0.00018986 3.3 0.00018996 0 0.00018988 0 0.00018998 3.3 0.00018989999999999998 3.3 0.00018999999999999998 0 0.00018992 0 0.00019002 3.3 0.00018994 3.3 0.00019004 0 0.00018996 0 0.00019006 3.3 0.00018998 3.3 0.00019008 0 0.00018999999999999998 0 0.00019009999999999999 3.3 0.00019002 3.3 0.00019012 0 0.00019004 0 0.00019014 3.3 0.00019006 3.3 0.00019016 0 0.00019008 0 0.00019018 3.3 0.00019009999999999999 3.3 0.0001902 0 0.00019012 0 0.00019022 3.3 0.00019014 3.3 0.00019024 0 0.00019015999999999998 0 0.00019025999999999998 3.3 0.00019018 3.3 0.00019028 0 0.0001902 0 0.0001903 3.3 0.00019022 3.3 0.00019032 0 0.00019024 0 0.00019034 3.3 0.00019025999999999998 3.3 0.00019036 0 0.00019028 0 0.00019038 3.3 0.0001903 3.3 0.0001904 0 0.00019031999999999998 0 0.00019041999999999998 3.3 0.00019034 3.3 0.00019044 0 0.00019036 0 0.00019046 3.3 0.00019038 3.3 0.00019048 0 0.0001904 0 0.0001905 3.3 0.00019041999999999998 3.3 0.00019051999999999999 0 0.00019044 0 0.00019054 3.3 0.00019046 3.3 0.00019056 0 0.00019048 0 0.00019058 3.3 0.0001905 3.3 0.0001906 0 0.00019051999999999999 0 0.00019062 3.3 0.00019054 3.3 0.00019064 0 0.00019056 0 0.00019066 3.3 0.00019057999999999998 3.3 0.00019067999999999998 0 0.0001906 0 0.0001907 3.3 0.00019062 3.3 0.00019072 0 0.00019064 0 0.00019074 3.3 0.00019066 3.3 0.00019076 0 0.00019067999999999998 0 0.00019077999999999999 3.3 0.0001907 3.3 0.0001908 0 0.00019072 0 0.00019082 3.3 0.00019074 3.3 0.00019084 0 0.00019076 0 0.00019086 3.3 0.00019077999999999999 3.3 0.00019088 0 0.0001908 0 0.0001909 3.3 0.00019082 3.3 0.00019092 0 0.00019083999999999998 0 0.00019093999999999998 3.3 0.00019086 3.3 0.00019096 0 0.00019088 0 0.00019098 3.3 0.0001909 3.3 0.000191 0 0.00019092 0 0.00019102 3.3 0.00019093999999999998 3.3 0.00019104 0 0.00019096 0 0.00019106 3.3 0.00019098 3.3 0.00019108 0 0.00019099999999999998 0 0.00019109999999999998 3.3 0.00019102 3.3 0.00019112 0 0.00019104 0 0.00019114 3.3 0.00019106 3.3 0.00019116 0 0.00019108 0 0.00019118 3.3 0.00019109999999999998 3.3 0.00019119999999999999 0 0.00019112 0 0.00019122 3.3 0.00019114 3.3 0.00019124 0 0.00019116 0 0.00019126 3.3 0.00019118 3.3 0.00019128 0 0.00019119999999999999 0 0.0001913 3.3 0.00019122 3.3 0.00019132 0 0.00019124 0 0.00019134 3.3 0.00019125999999999998 3.3 0.00019135999999999998 0 0.00019128 0 0.00019138 3.3 0.0001913 3.3 0.0001914 0 0.00019132 0 0.00019142 3.3 0.00019134 3.3 0.00019144 0 0.00019135999999999998 0 0.00019145999999999999 3.3 0.00019138 3.3 0.00019148 0 0.0001914 0 0.0001915 3.3 0.00019142 3.3 0.00019152 0 0.00019144 0 0.00019154 3.3 0.00019145999999999999 3.3 0.00019156 0 0.00019148 0 0.00019158 3.3 0.0001915 3.3 0.0001916 0 0.00019151999999999998 0 0.00019161999999999998 3.3 0.00019154 3.3 0.00019164 0 0.00019156 0 0.00019166 3.3 0.00019158 3.3 0.00019168 0 0.0001916 0 0.0001917 3.3 0.00019161999999999998 3.3 0.00019172 0 0.00019164 0 0.00019174 3.3 0.00019166 3.3 0.00019176 0 0.00019167999999999998 0 0.00019177999999999998 3.3 0.0001917 3.3 0.0001918 0 0.00019172 0 0.00019182 3.3 0.00019174 3.3 0.00019184 0 0.00019176 0 0.00019186 3.3 0.00019177999999999998 3.3 0.00019187999999999999 0 0.0001918 0 0.0001919 3.3 0.00019182 3.3 0.00019192 0 0.00019184 0 0.00019194 3.3 0.00019186 3.3 0.00019196 0 0.00019187999999999999 0 0.00019198 3.3 0.0001919 3.3 0.000192 0 0.00019192 0 0.00019202 3.3 0.00019193999999999998 3.3 0.00019203999999999998 0 0.00019196 0 0.00019206 3.3 0.00019198 3.3 0.00019208 0 0.000192 0 0.0001921 3.3 0.00019202 3.3 0.00019212 0 0.00019203999999999998 0 0.00019214 3.3 0.00019206 3.3 0.00019216 0 0.00019208 0 0.00019218 3.3 0.00019209999999999998 3.3 0.00019219999999999998 0 0.00019212 0 0.00019222 3.3 0.00019214 3.3 0.00019224 0 0.00019216 0 0.00019226 3.3 0.00019218 3.3 0.00019228 0 0.00019219999999999998 0 0.00019229999999999999 3.3 0.00019222 3.3 0.00019232 0 0.00019224 0 0.00019234 3.3 0.00019226 3.3 0.00019236 0 0.00019228 0 0.00019238 3.3 0.00019229999999999999 3.3 0.0001924 0 0.00019232 0 0.00019242 3.3 0.00019234 3.3 0.00019244 0 0.00019235999999999998 0 0.00019245999999999998 3.3 0.00019238 3.3 0.00019248 0 0.0001924 0 0.0001925 3.3 0.00019242 3.3 0.00019252 0 0.00019244 0 0.00019254 3.3 0.00019245999999999998 3.3 0.00019255999999999999 0 0.00019248 0 0.00019258 3.3 0.0001925 3.3 0.0001926 0 0.00019252 0 0.00019262 3.3 0.00019254 3.3 0.00019264 0 0.00019255999999999999 0 0.00019266 3.3 0.00019258 3.3 0.00019268 0 0.0001926 0 0.0001927 3.3 0.00019261999999999998 3.3 0.00019271999999999998 0 0.00019264 0 0.00019274 3.3 0.00019266 3.3 0.00019276 0 0.00019268 0 0.00019278 3.3 0.0001927 3.3 0.0001928 0 0.00019271999999999998 0 0.00019282 3.3 0.00019274 3.3 0.00019284 0 0.00019276 0 0.00019286 3.3 0.00019277999999999998 3.3 0.00019287999999999998 0 0.0001928 0 0.0001929 3.3 0.00019282 3.3 0.00019292 0 0.00019284 0 0.00019294 3.3 0.00019286 3.3 0.00019296 0 0.00019287999999999998 0 0.00019297999999999999 3.3 0.0001929 3.3 0.000193 0 0.00019292 0 0.00019302 3.3 0.00019294 3.3 0.00019304 0 0.00019296 0 0.00019306 3.3 0.00019297999999999999 3.3 0.00019308 0 0.000193 0 0.0001931 3.3 0.00019302 3.3 0.00019312 0 0.00019303999999999998 0 0.00019313999999999998 3.3 0.00019306 3.3 0.00019316 0 0.00019308 0 0.00019318 3.3 0.0001931 3.3 0.0001932 0 0.00019312 0 0.00019322 3.3 0.00019313999999999998 3.3 0.00019323999999999999 0 0.00019316 0 0.00019326 3.3 0.00019318 3.3 0.00019328 0 0.0001932 0 0.0001933 3.3 0.00019322 3.3 0.00019332 0 0.00019323999999999999 0 0.00019334 3.3 0.00019326 3.3 0.00019336 0 0.00019328 0 0.00019338 3.3 0.00019329999999999998 3.3 0.00019339999999999998 0 0.00019332 0 0.00019342 3.3 0.00019334 3.3 0.00019344 0 0.00019336 0 0.00019346 3.3 0.00019338 3.3 0.00019348 0 0.00019339999999999998 0 0.0001935 3.3 0.00019342 3.3 0.00019352 0 0.00019344 0 0.00019354 3.3 0.00019345999999999998 3.3 0.00019355999999999998 0 0.00019348 0 0.00019358 3.3 0.0001935 3.3 0.0001936 0 0.00019352 0 0.00019362 3.3 0.00019354 3.3 0.00019364 0 0.00019355999999999998 0 0.00019365999999999999 3.3 0.00019358 3.3 0.00019368 0 0.0001936 0 0.0001937 3.3 0.00019362 3.3 0.00019372 0 0.00019364 0 0.00019374 3.3 0.00019365999999999999 3.3 0.00019376 0 0.00019368 0 0.00019378 3.3 0.0001937 3.3 0.0001938 0 0.00019371999999999998 0 0.00019381999999999998 3.3 0.00019374 3.3 0.00019384 0 0.00019376 0 0.00019386 3.3 0.00019378 3.3 0.00019388 0 0.0001938 0 0.0001939 3.3 0.00019381999999999998 3.3 0.00019392 0 0.00019384 0 0.00019394 3.3 0.00019386 3.3 0.00019396 0 0.00019388 0 0.00019398 3.3 0.0001939 3.3 0.000194 0 0.00019392 0 0.00019402 3.3 0.00019394 3.3 0.00019404 0 0.00019396 0 0.00019406 3.3 0.00019397999999999998 3.3 0.00019407999999999998 0 0.000194 0 0.0001941 3.3 0.00019402 3.3 0.00019412 0 0.00019404 0 0.00019414 3.3 0.00019406 3.3 0.00019416 0 0.00019407999999999998 0 0.00019418 3.3 0.0001941 3.3 0.0001942 0 0.00019412 0 0.00019422 3.3 0.00019413999999999998 3.3 0.00019423999999999998 0 0.00019416 0 0.00019426 3.3 0.00019418 3.3 0.00019428 0 0.0001942 0 0.0001943 3.3 0.00019422 3.3 0.00019432 0 0.00019423999999999998 0 0.00019433999999999999 3.3 0.00019426 3.3 0.00019436 0 0.00019428 0 0.00019438 3.3 0.0001943 3.3 0.0001944 0 0.00019432 0 0.00019442 3.3 0.00019433999999999999 3.3 0.00019444 0 0.00019436 0 0.00019446 3.3 0.00019438 3.3 0.00019448 0 0.00019439999999999998 0 0.00019449999999999998 3.3 0.00019442 3.3 0.00019452 0 0.00019444 0 0.00019454 3.3 0.00019446 3.3 0.00019456 0 0.00019448 0 0.00019458 3.3 0.00019449999999999998 3.3 0.0001946 0 0.00019452 0 0.00019462 3.3 0.00019454 3.3 0.00019464 0 0.00019455999999999998 0 0.00019465999999999998 3.3 0.00019458 3.3 0.00019468 0 0.0001946 0 0.0001947 3.3 0.00019462 3.3 0.00019472 0 0.00019464 0 0.00019474 3.3 0.00019465999999999998 3.3 0.00019475999999999999 0 0.00019468 0 0.00019478 3.3 0.0001947 3.3 0.0001948 0 0.00019472 0 0.00019482 3.3 0.00019474 3.3 0.00019484 0 0.00019475999999999999 0 0.00019486 3.3 0.00019478 3.3 0.00019488 0 0.0001948 0 0.0001949 3.3 0.00019481999999999998 3.3 0.00019491999999999998 0 0.00019484 0 0.00019494 3.3 0.00019486 3.3 0.00019496 0 0.00019488 0 0.00019498 3.3 0.0001949 3.3 0.000195 0 0.00019491999999999998 0 0.00019501999999999999 3.3 0.00019494 3.3 0.00019504 0 0.00019496 0 0.00019506 3.3 0.00019498 3.3 0.00019508 0 0.000195 0 0.0001951 3.3 0.00019501999999999999 3.3 0.00019512 0 0.00019504 0 0.00019514 3.3 0.00019506 3.3 0.00019516 0 0.00019507999999999998 0 0.00019517999999999998 3.3 0.0001951 3.3 0.0001952 0 0.00019512 0 0.00019522 3.3 0.00019514 3.3 0.00019524 0 0.00019516 0 0.00019526 3.3 0.00019517999999999998 3.3 0.00019528 0 0.0001952 0 0.0001953 3.3 0.00019522 3.3 0.00019532 0 0.00019523999999999998 0 0.00019533999999999998 3.3 0.00019526 3.3 0.00019536 0 0.00019528 0 0.00019538 3.3 0.0001953 3.3 0.0001954 0 0.00019532 0 0.00019542 3.3 0.00019533999999999998 3.3 0.00019543999999999999 0 0.00019536 0 0.00019546 3.3 0.00019538 3.3 0.00019548 0 0.0001954 0 0.0001955 3.3 0.00019542 3.3 0.00019552 0 0.00019543999999999999 0 0.00019554 3.3 0.00019546 3.3 0.00019556 0 0.00019548 0 0.00019558 3.3 0.00019549999999999998 3.3 0.00019559999999999998 0 0.00019552 0 0.00019562 3.3 0.00019554 3.3 0.00019564 0 0.00019556 0 0.00019566 3.3 0.00019558 3.3 0.00019568 0 0.00019559999999999998 0 0.00019569999999999999 3.3 0.00019562 3.3 0.00019572 0 0.00019564 0 0.00019574 3.3 0.00019566 3.3 0.00019576 0 0.00019568 0 0.00019578 3.3 0.00019569999999999999 3.3 0.0001958 0 0.00019572 0 0.00019582 3.3 0.00019574 3.3 0.00019584 0 0.00019575999999999998 0 0.00019585999999999998 3.3 0.00019578 3.3 0.00019588 0 0.0001958 0 0.0001959 3.3 0.00019582 3.3 0.00019592 0 0.00019584 0 0.00019594 3.3 0.00019585999999999998 3.3 0.00019596 0 0.00019588 0 0.00019598 3.3 0.0001959 3.3 0.000196 0 0.00019591999999999998 0 0.00019601999999999998 3.3 0.00019594 3.3 0.00019604 0 0.00019596 0 0.00019606 3.3 0.00019598 3.3 0.00019608 0 0.000196 0 0.0001961 3.3 0.00019601999999999998 3.3 0.00019611999999999999 0 0.00019604 0 0.00019614 3.3 0.00019606 3.3 0.00019616 0 0.00019608 0 0.00019618 3.3 0.0001961 3.3 0.0001962 0 0.00019611999999999999 0 0.00019622 3.3 0.00019614 3.3 0.00019624 0 0.00019616 0 0.00019626 3.3 0.00019617999999999998 3.3 0.00019627999999999998 0 0.0001962 0 0.0001963 3.3 0.00019622 3.3 0.00019632 0 0.00019624 0 0.00019634 3.3 0.00019626 3.3 0.00019636 0 0.00019627999999999998 0 0.00019638 3.3 0.0001963 3.3 0.0001964 0 0.00019632 0 0.00019642 3.3 0.00019633999999999998 3.3 0.00019643999999999998 0 0.00019636 0 0.00019646 3.3 0.00019638 3.3 0.00019648 0 0.0001964 0 0.0001965 3.3 0.00019642 3.3 0.00019652 0 0.00019643999999999998 0 0.00019653999999999999 3.3 0.00019646 3.3 0.00019656 0 0.00019648 0 0.00019658 3.3 0.0001965 3.3 0.0001966 0 0.00019652 0 0.00019662 3.3 0.00019653999999999999 3.3 0.00019664 0 0.00019656 0 0.00019666 3.3 0.00019658 3.3 0.00019668 0 0.00019659999999999998 0 0.00019669999999999998 3.3 0.00019662 3.3 0.00019672 0 0.00019664 0 0.00019674 3.3 0.00019666 3.3 0.00019676 0 0.00019668 0 0.00019678 3.3 0.00019669999999999998 3.3 0.00019679999999999999 0 0.00019672 0 0.00019682 3.3 0.00019674 3.3 0.00019684 0 0.00019676 0 0.00019686 3.3 0.00019678 3.3 0.00019688 0 0.00019679999999999999 0 0.0001969 3.3 0.00019682 3.3 0.00019692 0 0.00019684 0 0.00019694 3.3 0.00019685999999999998 3.3 0.00019695999999999998 0 0.00019688 0 0.00019698 3.3 0.0001969 3.3 0.000197 0 0.00019692 0 0.00019702 3.3 0.00019694 3.3 0.00019704 0 0.00019695999999999998 0 0.00019706 3.3 0.00019698 3.3 0.00019708 0 0.000197 0 0.0001971 3.3 0.00019701999999999998 3.3 0.00019711999999999998 0 0.00019704 0 0.00019714 3.3 0.00019706 3.3 0.00019716 0 0.00019708 0 0.00019718 3.3 0.0001971 3.3 0.0001972 0 0.00019711999999999998 0 0.00019721999999999999 3.3 0.00019714 3.3 0.00019724 0 0.00019716 0 0.00019726 3.3 0.00019718 3.3 0.00019728 0 0.0001972 0 0.0001973 3.3 0.00019721999999999999 3.3 0.00019732 0 0.00019724 0 0.00019734 3.3 0.00019726 3.3 0.00019736 0 0.00019727999999999998 0 0.00019737999999999998 3.3 0.0001973 3.3 0.0001974 0 0.00019732 0 0.00019742 3.3 0.00019734 3.3 0.00019744 0 0.00019736 0 0.00019746 3.3 0.00019737999999999998 3.3 0.00019747999999999999 0 0.0001974 0 0.0001975 3.3 0.00019742 3.3 0.00019752 0 0.00019744 0 0.00019754 3.3 0.00019746 3.3 0.00019756 0 0.00019747999999999999 0 0.00019758 3.3 0.0001975 3.3 0.0001976 0 0.00019752 0 0.00019762 3.3 0.00019753999999999998 3.3 0.00019763999999999998 0 0.00019756 0 0.00019766 3.3 0.00019758 3.3 0.00019768 0 0.0001976 0 0.0001977 3.3 0.00019762 3.3 0.00019772 0 0.00019763999999999998 0 0.00019774 3.3 0.00019766 3.3 0.00019776 0 0.00019768 0 0.00019778 3.3 0.00019769999999999998 3.3 0.00019779999999999998 0 0.00019772 0 0.00019782 3.3 0.00019774 3.3 0.00019784 0 0.00019776 0 0.00019786 3.3 0.00019778 3.3 0.00019788 0 0.00019779999999999998 0 0.00019789999999999999 3.3 0.00019782 3.3 0.00019792 0 0.00019784 0 0.00019794 3.3 0.00019786 3.3 0.00019796 0 0.00019788 0 0.00019798 3.3 0.00019789999999999999 3.3 0.000198 0 0.00019792 0 0.00019802 3.3 0.00019794 3.3 0.00019804 0 0.00019795999999999998 0 0.00019805999999999998 3.3 0.00019798 3.3 0.00019808 0 0.000198 0 0.0001981 3.3 0.00019802 3.3 0.00019812 0 0.00019804 0 0.00019814 3.3 0.00019805999999999998 3.3 0.00019816 0 0.00019808 0 0.00019818 3.3 0.0001981 3.3 0.0001982 0 0.00019811999999999998 0 0.00019821999999999998 3.3 0.00019814 3.3 0.00019824 0 0.00019816 0 0.00019826 3.3 0.00019818 3.3 0.00019828 0 0.0001982 0 0.0001983 3.3 0.00019821999999999998 3.3 0.00019831999999999999 0 0.00019824 0 0.00019834 3.3 0.00019826 3.3 0.00019836 0 0.00019828 0 0.00019838 3.3 0.0001983 3.3 0.0001984 0 0.00019831999999999999 0 0.00019842 3.3 0.00019834 3.3 0.00019844 0 0.00019836 0 0.00019846 3.3 0.00019837999999999998 3.3 0.00019847999999999998 0 0.0001984 0 0.0001985 3.3 0.00019842 3.3 0.00019852 0 0.00019844 0 0.00019854 3.3 0.00019846 3.3 0.00019856 0 0.00019847999999999998 0 0.00019857999999999999 3.3 0.0001985 3.3 0.0001986 0 0.00019852 0 0.00019862 3.3 0.00019854 3.3 0.00019864 0 0.00019856 0 0.00019866 3.3 0.00019857999999999999 3.3 0.00019868 0 0.0001986 0 0.0001987 3.3 0.00019862 3.3 0.00019872 0 0.00019863999999999998 0 0.00019873999999999998 3.3 0.00019866 3.3 0.00019876 0 0.00019868 0 0.00019878 3.3 0.0001987 3.3 0.0001988 0 0.00019872 0 0.00019882 3.3 0.00019873999999999998 3.3 0.00019884 0 0.00019876 0 0.00019886 3.3 0.00019878 3.3 0.00019888 0 0.00019879999999999998 0 0.00019889999999999998 3.3 0.00019882 3.3 0.00019892 0 0.00019884 0 0.00019894 3.3 0.00019886 3.3 0.00019896 0 0.00019888 0 0.00019898 3.3 0.00019889999999999998 3.3 0.00019899999999999999 0 0.00019892 0 0.00019902 3.3 0.00019894 3.3 0.00019904 0 0.00019896 0 0.00019906 3.3 0.00019898 3.3 0.00019908 0 0.00019899999999999999 0 0.0001991 3.3 0.00019902 3.3 0.00019912 0 0.00019904 0 0.00019914 3.3 0.00019905999999999998 3.3 0.00019915999999999998 0 0.00019908 0 0.00019918 3.3 0.0001991 3.3 0.0001992 0 0.00019912 0 0.00019922 3.3 0.00019914 3.3 0.00019924 0 0.00019915999999999998 0 0.00019925999999999999 3.3 0.00019918 3.3 0.00019928 0 0.0001992 0 0.0001993 3.3 0.00019922 3.3 0.00019932 0 0.00019924 0 0.00019934 3.3 0.00019925999999999999 3.3 0.00019936 0 0.00019928 0 0.00019938 3.3 0.0001993 3.3 0.0001994 0 0.00019931999999999998 0 0.00019941999999999998 3.3 0.00019934 3.3 0.00019944 0 0.00019936 0 0.00019946 3.3 0.00019938 3.3 0.00019948 0 0.0001994 0 0.0001995 3.3 0.00019941999999999998 3.3 0.00019952 0 0.00019944 0 0.00019954 3.3 0.00019946 3.3 0.00019956 0 0.00019947999999999998 0 0.00019957999999999998 3.3 0.0001995 3.3 0.0001996 0 0.00019952 0 0.00019962 3.3 0.00019954 3.3 0.00019964 0 0.00019956 0 0.00019966 3.3 0.00019957999999999998 3.3 0.00019967999999999999 0 0.0001996 0 0.0001997 3.3 0.00019962 3.3 0.00019972 0 0.00019964 0 0.00019974 3.3 0.00019966 3.3 0.00019976 0 0.00019967999999999999 0 0.00019978 3.3 0.0001997 3.3 0.0001998 0 0.00019972 0 0.00019982 3.3 0.00019973999999999998 3.3 0.00019983999999999998 0 0.00019976 0 0.00019986 3.3 0.00019978 3.3 0.00019988 0 0.0001998 0 0.0001999 3.3 0.00019982 3.3 0.00019992 0 0.00019983999999999998 0 0.00019993999999999999 3.3 0.00019986 3.3 0.00019996 0 0.00019988 0 0.00019998 3.3 0.00019989999999999998 3.3 0.00019999999999999998 0 0.00019992 0 0.00020002 3.3 0.00019993999999999999 3.3 0.00020004 0 0.00019996 0 0.00020006 3.3 0.00019998 3.3 0.00020008 0 0.00019999999999999998 0 0.00020009999999999998 3.3 0.00020002 3.3 0.00020012 0 0.00020004 0 0.00020014 3.3 0.00020006 3.3 0.00020016 0 0.00020008 0 0.00020018 3.3 0.00020009999999999998 3.3 0.0002002 0 0.00020012 0 0.00020022 3.3 0.00020014 3.3 0.00020024 0 0.00020015999999999998 0 0.00020025999999999998 3.3 0.00020018 3.3 0.00020028 0 0.0002002 0 0.0002003 3.3 0.00020022 3.3 0.00020032 0 0.00020024 0 0.00020034 3.3 0.00020025999999999998 3.3 0.00020035999999999999 0 0.00020028 0 0.00020038 3.3 0.0002003 3.3 0.0002004 0 0.00020032 0 0.00020042 3.3 0.00020034 3.3 0.00020044 0 0.00020035999999999999 0 0.00020046 3.3 0.00020038 3.3 0.00020048 0 0.0002004 0 0.0002005 3.3 0.00020041999999999998 3.3 0.00020051999999999998 0 0.00020044 0 0.00020054 3.3 0.00020046 3.3 0.00020056 0 0.00020048 0 0.00020058 3.3 0.0002005 3.3 0.0002006 0 0.00020051999999999998 0 0.00020062 3.3 0.00020054 3.3 0.00020064 0 0.00020056 0 0.00020066 3.3 0.00020057999999999998 3.3 0.00020067999999999998 0 0.0002006 0 0.0002007 3.3 0.00020062 3.3 0.00020072 0 0.00020064 0 0.00020074 3.3 0.00020066 3.3 0.00020076 0 0.00020067999999999998 0 0.00020077999999999999 3.3 0.0002007 3.3 0.0002008 0 0.00020072 0 0.00020082 3.3 0.00020074 3.3 0.00020084 0 0.00020076 0 0.00020086 3.3 0.00020077999999999999 3.3 0.00020088 0 0.0002008 0 0.0002009 3.3 0.00020082 3.3 0.00020092 0 0.00020083999999999998 0 0.00020093999999999998 3.3 0.00020086 3.3 0.00020096 0 0.00020088 0 0.00020098 3.3 0.0002009 3.3 0.000201 0 0.00020092 0 0.00020102 3.3 0.00020093999999999998 3.3 0.00020103999999999999 0 0.00020096 0 0.00020106 3.3 0.00020098 3.3 0.00020108 0 0.000201 0 0.0002011 3.3 0.00020102 3.3 0.00020112 0 0.00020103999999999999 0 0.00020114 3.3 0.00020106 3.3 0.00020116 0 0.00020108 0 0.00020118 3.3 0.00020109999999999998 3.3 0.00020119999999999998 0 0.00020112 0 0.00020122 3.3 0.00020114 3.3 0.00020124 0 0.00020116 0 0.00020126 3.3 0.00020118 3.3 0.00020128 0 0.00020119999999999998 0 0.0002013 3.3 0.00020122 3.3 0.00020132 0 0.00020124 0 0.00020134 3.3 0.00020125999999999998 3.3 0.00020135999999999998 0 0.00020128 0 0.00020138 3.3 0.0002013 3.3 0.0002014 0 0.00020132 0 0.00020142 3.3 0.00020134 3.3 0.00020144 0 0.00020135999999999998 0 0.00020145999999999999 3.3 0.00020138 3.3 0.00020148 0 0.0002014 0 0.0002015 3.3 0.00020142 3.3 0.00020152 0 0.00020144 0 0.00020154 3.3 0.00020145999999999999 3.3 0.00020156 0 0.00020148 0 0.00020158 3.3 0.0002015 3.3 0.0002016 0 0.00020151999999999998 0 0.00020161999999999998 3.3 0.00020154 3.3 0.00020164 0 0.00020156 0 0.00020166 3.3 0.00020158 3.3 0.00020168 0 0.0002016 0 0.0002017 3.3 0.00020161999999999998 3.3 0.00020171999999999999 0 0.00020164 0 0.00020174 3.3 0.00020166 3.3 0.00020176 0 0.00020168 0 0.00020178 3.3 0.0002017 3.3 0.0002018 0 0.00020171999999999999 0 0.00020182 3.3 0.00020174 3.3 0.00020184 0 0.00020176 0 0.00020186 3.3 0.00020177999999999998 3.3 0.00020187999999999998 0 0.0002018 0 0.0002019 3.3 0.00020182 3.3 0.00020192 0 0.00020184 0 0.00020194 3.3 0.00020186 3.3 0.00020196 0 0.00020187999999999998 0 0.00020198 3.3 0.0002019 3.3 0.000202 0 0.00020192 0 0.00020202 3.3 0.00020193999999999998 3.3 0.00020203999999999998 0 0.00020196 0 0.00020206 3.3 0.00020198 3.3 0.00020208 0 0.000202 0 0.0002021 3.3 0.00020202 3.3 0.00020212 0 0.00020203999999999998 0 0.00020213999999999999 3.3 0.00020206 3.3 0.00020216 0 0.00020208 0 0.00020218 3.3 0.0002021 3.3 0.0002022 0 0.00020212 0 0.00020222 3.3 0.00020213999999999999 3.3 0.00020224 0 0.00020216 0 0.00020226 3.3 0.00020218 3.3 0.00020228 0 0.00020219999999999998 0 0.00020229999999999998 3.3 0.00020222 3.3 0.00020232 0 0.00020224 0 0.00020234 3.3 0.00020226 3.3 0.00020236 0 0.00020228 0 0.00020238 3.3 0.00020229999999999998 3.3 0.0002024 0 0.00020232 0 0.00020242 3.3 0.00020234 3.3 0.00020244 0 0.00020235999999999998 0 0.00020245999999999998 3.3 0.00020238 3.3 0.00020248 0 0.0002024 0 0.0002025 3.3 0.00020242 3.3 0.00020252 0 0.00020244 0 0.00020254 3.3 0.00020245999999999998 3.3 0.00020255999999999999 0 0.00020248 0 0.00020258 3.3 0.0002025 3.3 0.0002026 0 0.00020252 0 0.00020262 3.3 0.00020254 3.3 0.00020264 0 0.00020255999999999999 0 0.00020266 3.3 0.00020258 3.3 0.00020268 0 0.0002026 0 0.0002027 3.3 0.00020261999999999998 3.3 0.00020271999999999998 0 0.00020264 0 0.00020274 3.3 0.00020266 3.3 0.00020276 0 0.00020268 0 0.00020278 3.3 0.0002027 3.3 0.0002028 0 0.00020271999999999998 0 0.00020281999999999999 3.3 0.00020274 3.3 0.00020284 0 0.00020276 0 0.00020286 3.3 0.00020278 3.3 0.00020288 0 0.0002028 0 0.0002029 3.3 0.00020281999999999999 3.3 0.00020292 0 0.00020284 0 0.00020294 3.3 0.00020286 3.3 0.00020296 0 0.00020287999999999998 0 0.00020297999999999998 3.3 0.0002029 3.3 0.000203 0 0.00020292 0 0.00020302 3.3 0.00020294 3.3 0.00020304 0 0.00020296 0 0.00020306 3.3 0.00020297999999999998 3.3 0.00020308 0 0.000203 0 0.0002031 3.3 0.00020302 3.3 0.00020312 0 0.00020303999999999998 0 0.00020313999999999998 3.3 0.00020306 3.3 0.00020316 0 0.00020308 0 0.00020318 3.3 0.0002031 3.3 0.0002032 0 0.00020312 0 0.00020322 3.3 0.00020313999999999998 3.3 0.00020323999999999999 0 0.00020316 0 0.00020326 3.3 0.00020318 3.3 0.00020328 0 0.0002032 0 0.0002033 3.3 0.00020322 3.3 0.00020332 0 0.00020323999999999999 0 0.00020334 3.3 0.00020326 3.3 0.00020336 0 0.00020328 0 0.00020338 3.3 0.00020329999999999998 3.3 0.00020339999999999998 0 0.00020332 0 0.00020342 3.3 0.00020334 3.3 0.00020344 0 0.00020336 0 0.00020346 3.3 0.00020338 3.3 0.00020348 0 0.00020339999999999998 0 0.00020349999999999999 3.3 0.00020342 3.3 0.00020352 0 0.00020344 0 0.00020354 3.3 0.00020346 3.3 0.00020356 0 0.00020348 0 0.00020358 3.3 0.00020349999999999999 3.3 0.0002036 0 0.00020352 0 0.00020362 3.3 0.00020354 3.3 0.00020364 0 0.00020355999999999998 0 0.00020365999999999998 3.3 0.00020358 3.3 0.00020368 0 0.0002036 0 0.0002037 3.3 0.00020362 3.3 0.00020372 0 0.00020364 0 0.00020374 3.3 0.00020365999999999998 3.3 0.00020376 0 0.00020368 0 0.00020378 3.3 0.0002037 3.3 0.0002038 0 0.00020371999999999998 0 0.00020381999999999998 3.3 0.00020374 3.3 0.00020384 0 0.00020376 0 0.00020386 3.3 0.00020378 3.3 0.00020388 0 0.0002038 0 0.0002039 3.3 0.00020381999999999998 3.3 0.00020391999999999999 0 0.00020384 0 0.00020394 3.3 0.00020386 3.3 0.00020396 0 0.00020388 0 0.00020398 3.3 0.0002039 3.3 0.000204 0 0.00020391999999999999 0 0.00020402 3.3 0.00020394 3.3 0.00020404 0 0.00020396 0 0.00020406 3.3 0.00020397999999999998 3.3 0.00020407999999999998 0 0.000204 0 0.0002041 3.3 0.00020402 3.3 0.00020412 0 0.00020404 0 0.00020414 3.3 0.00020406 3.3 0.00020416 0 0.00020407999999999998 0 0.00020418 3.3 0.0002041 3.3 0.0002042 0 0.00020412 0 0.00020422 3.3 0.00020413999999999998 3.3 0.00020423999999999998 0 0.00020416 0 0.00020426 3.3 0.00020418 3.3 0.00020428 0 0.0002042 0 0.0002043 3.3 0.00020422 3.3 0.00020432 0 0.00020423999999999998 0 0.00020433999999999998 3.3 0.00020426 3.3 0.00020436 0 0.00020428 0 0.00020438 3.3 0.0002043 3.3 0.0002044 0 0.00020432 0 0.00020442 3.3 0.00020433999999999998 3.3 0.00020444 0 0.00020436 0 0.00020446 3.3 0.00020438 3.3 0.00020448 0 0.00020439999999999998 0 0.00020449999999999998 3.3 0.00020442 3.3 0.00020452 0 0.00020444 0 0.00020454 3.3 0.00020446 3.3 0.00020456 0 0.00020448 0 0.00020458 3.3 0.00020449999999999998 3.3 0.00020459999999999999 0 0.00020452 0 0.00020462 3.3 0.00020454 3.3 0.00020464 0 0.00020456 0 0.00020466 3.3 0.00020458 3.3 0.00020468 0 0.00020459999999999999 0 0.0002047 3.3 0.00020462 3.3 0.00020472 0 0.00020464 0 0.00020474 3.3 0.00020465999999999998 3.3 0.00020475999999999998 0 0.00020468 0 0.00020478 3.3 0.0002047 3.3 0.0002048 0 0.00020472 0 0.00020482 3.3 0.00020474 3.3 0.00020484 0 0.00020475999999999998 0 0.00020486 3.3 0.00020478 3.3 0.00020488 0 0.0002048 0 0.0002049 3.3 0.00020481999999999998 3.3 0.00020491999999999998 0 0.00020484 0 0.00020494 3.3 0.00020486 3.3 0.00020496 0 0.00020488 0 0.00020498 3.3 0.0002049 3.3 0.000205 0 0.00020491999999999998 0 0.00020501999999999999 3.3 0.00020494 3.3 0.00020504 0 0.00020496 0 0.00020506 3.3 0.00020498 3.3 0.00020508 0 0.000205 0 0.0002051 3.3 0.00020501999999999999 3.3 0.00020512 0 0.00020504 0 0.00020514 3.3 0.00020506 3.3 0.00020516 0 0.00020507999999999998 0 0.00020517999999999998 3.3 0.0002051 3.3 0.0002052 0 0.00020512 0 0.00020522 3.3 0.00020514 3.3 0.00020524 0 0.00020516 0 0.00020526 3.3 0.00020517999999999998 3.3 0.00020527999999999999 0 0.0002052 0 0.0002053 3.3 0.00020522 3.3 0.00020532 0 0.00020524 0 0.00020534 3.3 0.00020526 3.3 0.00020536 0 0.00020527999999999999 0 0.00020538 3.3 0.0002053 3.3 0.0002054 0 0.00020532 0 0.00020542 3.3 0.00020533999999999998 3.3 0.00020543999999999998 0 0.00020536 0 0.00020546 3.3 0.00020538 3.3 0.00020548 0 0.0002054 0 0.0002055 3.3 0.00020542 3.3 0.00020552 0 0.00020543999999999998 0 0.00020554 3.3 0.00020546 3.3 0.00020556 0 0.00020548 0 0.00020558 3.3 0.00020549999999999998 3.3 0.00020559999999999998 0 0.00020552 0 0.00020562 3.3 0.00020554 3.3 0.00020564 0 0.00020556 0 0.00020566 3.3 0.00020558 3.3 0.00020568 0 0.00020559999999999998 0 0.00020569999999999999 3.3 0.00020562 3.3 0.00020572 0 0.00020564 0 0.00020574 3.3 0.00020566 3.3 0.00020576 0 0.00020568 0 0.00020578 3.3 0.00020569999999999999 3.3 0.0002058 0 0.00020572 0 0.00020582 3.3 0.00020574 3.3 0.00020584 0 0.00020575999999999998 0 0.00020585999999999998 3.3 0.00020578 3.3 0.00020588 0 0.0002058 0 0.0002059 3.3 0.00020582 3.3 0.00020592 0 0.00020584 0 0.00020594 3.3 0.00020585999999999998 3.3 0.00020595999999999999 0 0.00020588 0 0.00020598 3.3 0.0002059 3.3 0.000206 0 0.00020591999999999998 0 0.00020601999999999998 3.3 0.00020594 3.3 0.00020604 0 0.00020595999999999999 0 0.00020606 3.3 0.00020598 3.3 0.00020608 0 0.000206 0 0.0002061 3.3 0.00020601999999999998 3.3 0.00020611999999999998 0 0.00020604 0 0.00020614 3.3 0.00020606 3.3 0.00020616 0 0.00020608 0 0.00020618 3.3 0.0002061 3.3 0.0002062 0 0.00020611999999999998 0 0.00020622 3.3 0.00020614 3.3 0.00020624 0 0.00020616 0 0.00020626 3.3 0.00020617999999999998 3.3 0.00020627999999999998 0 0.0002062 0 0.0002063 3.3 0.00020622 3.3 0.00020632 0 0.00020624 0 0.00020634 3.3 0.00020626 3.3 0.00020636 0 0.00020627999999999998 0 0.00020637999999999999 3.3 0.0002063 3.3 0.0002064 0 0.00020632 0 0.00020642 3.3 0.00020634 3.3 0.00020644 0 0.00020636 0 0.00020646 3.3 0.00020637999999999999 3.3 0.00020648 0 0.0002064 0 0.0002065 3.3 0.00020642 3.3 0.00020652 0 0.00020643999999999998 0 0.00020653999999999998 3.3 0.00020646 3.3 0.00020656 0 0.00020648 0 0.00020658 3.3 0.0002065 3.3 0.0002066 0 0.00020652 0 0.00020662 3.3 0.00020653999999999998 3.3 0.00020664 0 0.00020656 0 0.00020666 3.3 0.00020658 3.3 0.00020668 0 0.00020659999999999998 0 0.00020669999999999998 3.3 0.00020662 3.3 0.00020672 0 0.00020664 0 0.00020674 3.3 0.00020666 3.3 0.00020676 0 0.00020668 0 0.00020678 3.3 0.00020669999999999998 3.3 0.00020679999999999999 0 0.00020672 0 0.00020682 3.3 0.00020674 3.3 0.00020684 0 0.00020676 0 0.00020686 3.3 0.00020678 3.3 0.00020688 0 0.00020679999999999999 0 0.0002069 3.3 0.00020682 3.3 0.00020692 0 0.00020684 0 0.00020694 3.3 0.00020685999999999998 3.3 0.00020695999999999998 0 0.00020688 0 0.00020698 3.3 0.0002069 3.3 0.000207 0 0.00020692 0 0.00020702 3.3 0.00020694 3.3 0.00020704 0 0.00020695999999999998 0 0.00020705999999999999 3.3 0.00020698 3.3 0.00020708 0 0.000207 0 0.0002071 3.3 0.00020702 3.3 0.00020712 0 0.00020704 0 0.00020714 3.3 0.00020705999999999999 3.3 0.00020716 0 0.00020708 0 0.00020718 3.3 0.0002071 3.3 0.0002072 0 0.00020711999999999998 0 0.00020721999999999998 3.3 0.00020714 3.3 0.00020724 0 0.00020716 0 0.00020726 3.3 0.00020718 3.3 0.00020728 0 0.0002072 0 0.0002073 3.3 0.00020721999999999998 3.3 0.00020732 0 0.00020724 0 0.00020734 3.3 0.00020726 3.3 0.00020736 0 0.00020727999999999998 0 0.00020737999999999998 3.3 0.0002073 3.3 0.0002074 0 0.00020732 0 0.00020742 3.3 0.00020734 3.3 0.00020744 0 0.00020736 0 0.00020746 3.3 0.00020737999999999998 3.3 0.00020747999999999999 0 0.0002074 0 0.0002075 3.3 0.00020742 3.3 0.00020752 0 0.00020744 0 0.00020754 3.3 0.00020746 3.3 0.00020756 0 0.00020747999999999999 0 0.00020758 3.3 0.0002075 3.3 0.0002076 0 0.00020752 0 0.00020762 3.3 0.00020753999999999998 3.3 0.00020763999999999998 0 0.00020756 0 0.00020766 3.3 0.00020758 3.3 0.00020768 0 0.0002076 0 0.0002077 3.3 0.00020762 3.3 0.00020772 0 0.00020763999999999998 0 0.00020773999999999999 3.3 0.00020766 3.3 0.00020776 0 0.00020768 0 0.00020778 3.3 0.00020769999999999998 3.3 0.00020779999999999998 0 0.00020772 0 0.00020782 3.3 0.00020773999999999999 3.3 0.00020784 0 0.00020776 0 0.00020786 3.3 0.00020778 3.3 0.00020788 0 0.00020779999999999998 0 0.00020789999999999998 3.3 0.00020782 3.3 0.00020792 0 0.00020784 0 0.00020794 3.3 0.00020786 3.3 0.00020796 0 0.00020788 0 0.00020798 3.3 0.00020789999999999998 3.3 0.000208 0 0.00020792 0 0.00020802 3.3 0.00020794 3.3 0.00020804 0 0.00020795999999999998 0 0.00020805999999999998 3.3 0.00020798 3.3 0.00020808 0 0.000208 0 0.0002081 3.3 0.00020802 3.3 0.00020812 0 0.00020804 0 0.00020814 3.3 0.00020805999999999998 3.3 0.00020815999999999999 0 0.00020808 0 0.00020818 3.3 0.0002081 3.3 0.0002082 0 0.00020812 0 0.00020822 3.3 0.00020814 3.3 0.00020824 0 0.00020815999999999999 0 0.00020826 3.3 0.00020818 3.3 0.00020828 0 0.0002082 0 0.0002083 3.3 0.00020821999999999998 3.3 0.00020831999999999998 0 0.00020824 0 0.00020834 3.3 0.00020826 3.3 0.00020836 0 0.00020828 0 0.00020838 3.3 0.0002083 3.3 0.0002084 0 0.00020831999999999998 0 0.00020842 3.3 0.00020834 3.3 0.00020844 0 0.00020836 0 0.00020846 3.3 0.00020837999999999998 3.3 0.00020847999999999998 0 0.0002084 0 0.0002085 3.3 0.00020842 3.3 0.00020852 0 0.00020844 0 0.00020854 3.3 0.00020846 3.3 0.00020856 0 0.00020847999999999998 0 0.00020857999999999999 3.3 0.0002085 3.3 0.0002086 0 0.00020852 0 0.00020862 3.3 0.00020854 3.3 0.00020864 0 0.00020856 0 0.00020866 3.3 0.00020857999999999999 3.3 0.00020868 0 0.0002086 0 0.0002087 3.3 0.00020862 3.3 0.00020872 0 0.00020863999999999998 0 0.00020873999999999998 3.3 0.00020866 3.3 0.00020876 0 0.00020868 0 0.00020878 3.3 0.0002087 3.3 0.0002088 0 0.00020872 0 0.00020882 3.3 0.00020873999999999998 3.3 0.00020883999999999999 0 0.00020876 0 0.00020886 3.3 0.00020878 3.3 0.00020888 0 0.0002088 0 0.0002089 3.3 0.00020882 3.3 0.00020892 0 0.00020883999999999999 0 0.00020894 3.3 0.00020886 3.3 0.00020896 0 0.00020888 0 0.00020898 3.3 0.00020889999999999998 3.3 0.00020899999999999998 0 0.00020892 0 0.00020902 3.3 0.00020894 3.3 0.00020904 0 0.00020896 0 0.00020906 3.3 0.00020898 3.3 0.00020908 0 0.00020899999999999998 0 0.0002091 3.3 0.00020902 3.3 0.00020912 0 0.00020904 0 0.00020914 3.3 0.00020905999999999998 3.3 0.00020915999999999998 0 0.00020908 0 0.00020918 3.3 0.0002091 3.3 0.0002092 0 0.00020912 0 0.00020922 3.3 0.00020914 3.3 0.00020924 0 0.00020915999999999998 0 0.00020925999999999999 3.3 0.00020918 3.3 0.00020928 0 0.0002092 0 0.0002093 3.3 0.00020922 3.3 0.00020932 0 0.00020924 0 0.00020934 3.3 0.00020925999999999999 3.3 0.00020936 0 0.00020928 0 0.00020938 3.3 0.0002093 3.3 0.0002094 0 0.00020931999999999998 0 0.00020941999999999998 3.3 0.00020934 3.3 0.00020944 0 0.00020936 0 0.00020946 3.3 0.00020938 3.3 0.00020948 0 0.0002094 0 0.0002095 3.3 0.00020941999999999998 3.3 0.00020951999999999999 0 0.00020944 0 0.00020954 3.3 0.00020946 3.3 0.00020956 0 0.00020947999999999998 0 0.00020957999999999998 3.3 0.0002095 3.3 0.0002096 0 0.00020951999999999999 0 0.00020962 3.3 0.00020954 3.3 0.00020964 0 0.00020956 0 0.00020966 3.3 0.00020957999999999998 3.3 0.00020967999999999998 0 0.0002096 0 0.0002097 3.3 0.00020962 3.3 0.00020972 0 0.00020964 0 0.00020974 3.3 0.00020966 3.3 0.00020976 0 0.00020967999999999998 0 0.00020978 3.3 0.0002097 3.3 0.0002098 0 0.00020972 0 0.00020982 3.3 0.00020973999999999998 3.3 0.00020983999999999998 0 0.00020976 0 0.00020986 3.3 0.00020978 3.3 0.00020988 0 0.0002098 0 0.0002099 3.3 0.00020982 3.3 0.00020992 0 0.00020983999999999998 0 0.00020993999999999999 3.3 0.00020986 3.3 0.00020996 0 0.00020988 0 0.00020998 3.3 0.0002099 3.3 0.00021 0 0.00020992 0 0.00021002 3.3 0.00020993999999999999 3.3 0.00021004 0 0.00020996 0 0.00021006 3.3 0.00020998 3.3 0.00021008 0 0.00020999999999999998 0 0.00021009999999999998 3.3 0.00021002 3.3 0.00021012 0 0.00021004 0 0.00021014 3.3 0.00021006 3.3 0.00021016 0 0.00021008 0 0.00021018 3.3 0.00021009999999999998 3.3 0.0002102 0 0.00021012 0 0.00021022 3.3 0.00021014 3.3 0.00021024 0 0.00021015999999999998 0 0.00021025999999999998 3.3 0.00021018 3.3 0.00021028 0 0.0002102 0 0.0002103 3.3 0.00021022 3.3 0.00021032 0 0.00021024 0 0.00021034 3.3 0.00021025999999999998 3.3 0.00021035999999999998 0 0.00021028 0 0.00021038 3.3 0.0002103 3.3 0.0002104 0 0.00021032 0 0.00021042 3.3 0.00021034 3.3 0.00021044 0 0.00021035999999999998 0 0.00021046 3.3 0.00021038 3.3 0.00021048 0 0.0002104 0 0.0002105 3.3 0.00021041999999999998 3.3 0.00021051999999999998 0 0.00021044 0 0.00021054 3.3 0.00021046 3.3 0.00021056 0 0.00021048 0 0.00021058 3.3 0.0002105 3.3 0.0002106 0 0.00021051999999999998 0 0.00021061999999999999 3.3 0.00021054 3.3 0.00021064 0 0.00021056 0 0.00021066 3.3 0.00021058 3.3 0.00021068 0 0.0002106 0 0.0002107 3.3 0.00021061999999999999 3.3 0.00021072 0 0.00021064 0 0.00021074 3.3 0.00021066 3.3 0.00021076 0 0.00021067999999999998 0 0.00021077999999999998 3.3 0.0002107 3.3 0.0002108 0 0.00021072 0 0.00021082 3.3 0.00021074 3.3 0.00021084 0 0.00021076 0 0.00021086 3.3 0.00021077999999999998 3.3 0.00021088 0 0.0002108 0 0.0002109 3.3 0.00021082 3.3 0.00021092 0 0.00021083999999999998 0 0.00021093999999999998 3.3 0.00021086 3.3 0.00021096 0 0.00021088 0 0.00021098 3.3 0.0002109 3.3 0.000211 0 0.00021092 0 0.00021102 3.3 0.00021093999999999998 3.3 0.00021103999999999999 0 0.00021096 0 0.00021106 3.3 0.00021098 3.3 0.00021108 0 0.000211 0 0.0002111 3.3 0.00021102 3.3 0.00021112 0 0.00021103999999999999 0 0.00021114 3.3 0.00021106 3.3 0.00021116 0 0.00021108 0 0.00021118 3.3 0.00021109999999999998 3.3 0.00021119999999999998 0 0.00021112 0 0.00021122 3.3 0.00021114 3.3 0.00021124 0 0.00021116 0 0.00021126 3.3 0.00021118 3.3 0.00021128 0 0.00021119999999999998 0 0.00021129999999999999 3.3 0.00021122 3.3 0.00021132 0 0.00021124 0 0.00021134 3.3 0.00021126 3.3 0.00021136 0 0.00021128 0 0.00021138 3.3 0.00021129999999999999 3.3 0.0002114 0 0.00021132 0 0.00021142 3.3 0.00021134 3.3 0.00021144 0 0.00021135999999999998 0 0.00021145999999999998 3.3 0.00021138 3.3 0.00021148 0 0.0002114 0 0.0002115 3.3 0.00021142 3.3 0.00021152 0 0.00021144 0 0.00021154 3.3 0.00021145999999999998 3.3 0.00021156 0 0.00021148 0 0.00021158 3.3 0.0002115 3.3 0.0002116 0 0.00021151999999999998 0 0.00021161999999999998 3.3 0.00021154 3.3 0.00021164 0 0.00021156 0 0.00021166 3.3 0.00021158 3.3 0.00021168 0 0.0002116 0 0.0002117 3.3 0.00021161999999999998 3.3 0.00021171999999999999 0 0.00021164 0 0.00021174 3.3 0.00021166 3.3 0.00021176 0 0.00021168 0 0.00021178 3.3 0.0002117 3.3 0.0002118 0 0.00021171999999999999 0 0.00021182 3.3 0.00021174 3.3 0.00021184 0 0.00021176 0 0.00021186 3.3 0.00021177999999999998 3.3 0.00021187999999999998 0 0.0002118 0 0.0002119 3.3 0.00021182 3.3 0.00021192 0 0.00021184 0 0.00021194 3.3 0.00021186 3.3 0.00021196 0 0.00021187999999999998 0 0.00021197999999999999 3.3 0.0002119 3.3 0.000212 0 0.00021192 0 0.00021202 3.3 0.00021193999999999998 3.3 0.00021203999999999998 0 0.00021196 0 0.00021206 3.3 0.00021197999999999999 3.3 0.00021208 0 0.000212 0 0.0002121 3.3 0.00021202 3.3 0.00021212 0 0.00021203999999999998 0 0.00021213999999999998 3.3 0.00021206 3.3 0.00021216 0 0.00021208 0 0.00021218 3.3 0.0002121 3.3 0.0002122 0 0.00021212 0 0.00021222 3.3 0.00021213999999999998 3.3 0.00021224 0 0.00021216 0 0.00021226 3.3 0.00021218 3.3 0.00021228 0 0.00021219999999999998 0 0.00021229999999999998 3.3 0.00021222 3.3 0.00021232 0 0.00021224 0 0.00021234 3.3 0.00021226 3.3 0.00021236 0 0.00021228 0 0.00021238 3.3 0.00021229999999999998 3.3 0.00021239999999999999 0 0.00021232 0 0.00021242 3.3 0.00021234 3.3 0.00021244 0 0.00021236 0 0.00021246 3.3 0.00021238 3.3 0.00021248 0 0.00021239999999999999 0 0.0002125 3.3 0.00021242 3.3 0.00021252 0 0.00021244 0 0.00021254 3.3 0.00021245999999999998 3.3 0.00021255999999999998 0 0.00021248 0 0.00021258 3.3 0.0002125 3.3 0.0002126 0 0.00021252 0 0.00021262 3.3 0.00021254 3.3 0.00021264 0 0.00021255999999999998 0 0.00021266 3.3 0.00021258 3.3 0.00021268 0 0.0002126 0 0.0002127 3.3 0.00021261999999999998 3.3 0.00021271999999999998 0 0.00021264 0 0.00021274 3.3 0.00021266 3.3 0.00021276 0 0.00021268 0 0.00021278 3.3 0.0002127 3.3 0.0002128 0 0.00021271999999999998 0 0.00021281999999999999 3.3 0.00021274 3.3 0.00021284 0 0.00021276 0 0.00021286 3.3 0.00021278 3.3 0.00021288 0 0.0002128 0 0.0002129 3.3 0.00021281999999999999 3.3 0.00021292 0 0.00021284 0 0.00021294 3.3 0.00021286 3.3 0.00021296 0 0.00021287999999999998 0 0.00021297999999999998 3.3 0.0002129 3.3 0.000213 0 0.00021292 0 0.00021302 3.3 0.00021294 3.3 0.00021304 0 0.00021296 0 0.00021306 3.3 0.00021297999999999998 3.3 0.00021307999999999999 0 0.000213 0 0.0002131 3.3 0.00021302 3.3 0.00021312 0 0.00021304 0 0.00021314 3.3 0.00021306 3.3 0.00021316 0 0.00021307999999999999 0 0.00021318 3.3 0.0002131 3.3 0.0002132 0 0.00021312 0 0.00021322 3.3 0.00021313999999999998 3.3 0.00021323999999999998 0 0.00021316 0 0.00021326 3.3 0.00021318 3.3 0.00021328 0 0.0002132 0 0.0002133 3.3 0.00021322 3.3 0.00021332 0 0.00021323999999999998 0 0.00021334 3.3 0.00021326 3.3 0.00021336 0 0.00021328 0 0.00021338 3.3 0.00021329999999999998 3.3 0.00021339999999999998 0 0.00021332 0 0.00021342 3.3 0.00021334 3.3 0.00021344 0 0.00021336 0 0.00021346 3.3 0.00021338 3.3 0.00021348 0 0.00021339999999999998 0 0.00021349999999999999 3.3 0.00021342 3.3 0.00021352 0 0.00021344 0 0.00021354 3.3 0.00021346 3.3 0.00021356 0 0.00021348 0 0.00021358 3.3 0.00021349999999999999 3.3 0.0002136 0 0.00021352 0 0.00021362 3.3 0.00021354 3.3 0.00021364 0 0.00021355999999999998 0 0.00021365999999999998 3.3 0.00021358 3.3 0.00021368 0 0.0002136 0 0.0002137 3.3 0.00021362 3.3 0.00021372 0 0.00021364 0 0.00021374 3.3 0.00021365999999999998 3.3 0.00021375999999999999 0 0.00021368 0 0.00021378 3.3 0.0002137 3.3 0.0002138 0 0.00021371999999999998 0 0.00021381999999999998 3.3 0.00021374 3.3 0.00021384 0 0.00021375999999999999 0 0.00021386 3.3 0.00021378 3.3 0.00021388 0 0.0002138 0 0.0002139 3.3 0.00021381999999999998 3.3 0.00021391999999999998 0 0.00021384 0 0.00021394 3.3 0.00021386 3.3 0.00021396 0 0.00021388 0 0.00021398 3.3 0.0002139 3.3 0.000214 0 0.00021391999999999998 0 0.00021402 3.3 0.00021394 3.3 0.00021404 0 0.00021396 0 0.00021406 3.3 0.00021397999999999998 3.3 0.00021407999999999998 0 0.000214 0 0.0002141 3.3 0.00021402 3.3 0.00021412 0 0.00021404 0 0.00021414 3.3 0.00021406 3.3 0.00021416 0 0.00021407999999999998 0 0.00021417999999999999 3.3 0.0002141 3.3 0.0002142 0 0.00021412 0 0.00021422 3.3 0.00021414 3.3 0.00021424 0 0.00021416 0 0.00021426 3.3 0.00021417999999999999 3.3 0.00021428 0 0.0002142 0 0.0002143 3.3 0.00021422 3.3 0.00021432 0 0.00021423999999999998 0 0.00021433999999999998 3.3 0.00021426 3.3 0.00021436 0 0.00021428 0 0.00021438 3.3 0.0002143 3.3 0.0002144 0 0.00021432 0 0.00021442 3.3 0.00021433999999999998 3.3 0.00021444 0 0.00021436 0 0.00021446 3.3 0.00021438 3.3 0.00021448 0 0.00021439999999999998 0 0.00021449999999999998 3.3 0.00021442 3.3 0.00021452 0 0.00021444 0 0.00021454 3.3 0.00021446 3.3 0.00021456 0 0.00021448 0 0.00021458 3.3 0.00021449999999999998 3.3 0.00021459999999999998 0 0.00021452 0 0.00021462 3.3 0.00021454 3.3 0.00021464 0 0.00021456 0 0.00021466 3.3 0.00021458 3.3 0.00021468 0 0.00021459999999999998 0 0.0002147 3.3 0.00021462 3.3 0.00021472 0 0.00021464 0 0.00021474 3.3 0.00021465999999999998 3.3 0.00021475999999999998 0 0.00021468 0 0.00021478 3.3 0.0002147 3.3 0.0002148 0 0.00021472 0 0.00021482 3.3 0.00021474 3.3 0.00021484 0 0.00021475999999999998 0 0.00021485999999999999 3.3 0.00021478 3.3 0.00021488 0 0.0002148 0 0.0002149 3.3 0.00021482 3.3 0.00021492 0 0.00021484 0 0.00021494 3.3 0.00021485999999999999 3.3 0.00021496 0 0.00021488 0 0.00021498 3.3 0.0002149 3.3 0.000215 0 0.00021491999999999998 0 0.00021501999999999998 3.3 0.00021494 3.3 0.00021504 0 0.00021496 0 0.00021506 3.3 0.00021498 3.3 0.00021508 0 0.000215 0 0.0002151 3.3 0.00021501999999999998 3.3 0.00021512 0 0.00021504 0 0.00021514 3.3 0.00021506 3.3 0.00021516 0 0.00021507999999999998 0 0.00021517999999999998 3.3 0.0002151 3.3 0.0002152 0 0.00021512 0 0.00021522 3.3 0.00021514 3.3 0.00021524 0 0.00021516 0 0.00021526 3.3 0.00021517999999999998 3.3 0.00021527999999999999 0 0.0002152 0 0.0002153 3.3 0.00021522 3.3 0.00021532 0 0.00021524 0 0.00021534 3.3 0.00021526 3.3 0.00021536 0 0.00021527999999999999 0 0.00021538 3.3 0.0002153 3.3 0.0002154 0 0.00021532 0 0.00021542 3.3 0.00021533999999999998 3.3 0.00021543999999999998 0 0.00021536 0 0.00021546 3.3 0.00021538 3.3 0.00021548 0 0.0002154 0 0.0002155 3.3 0.00021542 3.3 0.00021552 0 0.00021543999999999998 0 0.00021553999999999999 3.3 0.00021546 3.3 0.00021556 0 0.00021548 0 0.00021558 3.3 0.00021549999999999998 3.3 0.00021559999999999998 0 0.00021552 0 0.00021562 3.3 0.00021553999999999999 3.3 0.00021564 0 0.00021556 0 0.00021566 3.3 0.00021558 3.3 0.00021568 0 0.00021559999999999998 0 0.00021569999999999998 3.3 0.00021562 3.3 0.00021572 0 0.00021564 0 0.00021574 3.3 0.00021566 3.3 0.00021576 0 0.00021568 0 0.00021578 3.3 0.00021569999999999998 3.3 0.0002158 0 0.00021572 0 0.00021582 3.3 0.00021574 3.3 0.00021584 0 0.00021575999999999998 0 0.00021585999999999998 3.3 0.00021578 3.3 0.00021588 0 0.0002158 0 0.0002159 3.3 0.00021582 3.3 0.00021592 0 0.00021584 0 0.00021594 3.3 0.00021585999999999998 3.3 0.00021595999999999999 0 0.00021588 0 0.00021598 3.3 0.0002159 3.3 0.000216 0 0.00021592 0 0.00021602 3.3 0.00021594 3.3 0.00021604 0 0.00021595999999999999 0 0.00021606 3.3 0.00021598 3.3 0.00021608 0 0.000216 0 0.0002161 3.3 0.00021601999999999998 3.3 0.00021611999999999998 0 0.00021604 0 0.00021614 3.3 0.00021606 3.3 0.00021616 0 0.00021608 0 0.00021618 3.3 0.0002161 3.3 0.0002162 0 0.00021611999999999998 0 0.00021621999999999999 3.3 0.00021614 3.3 0.00021624 0 0.00021616 0 0.00021626 3.3 0.00021617999999999998 3.3 0.00021627999999999998 0 0.0002162 0 0.0002163 3.3 0.00021621999999999999 3.3 0.00021632 0 0.00021624 0 0.00021634 3.3 0.00021626 3.3 0.00021636 0 0.00021627999999999998 0 0.00021637999999999998 3.3 0.0002163 3.3 0.0002164 0 0.00021632 0 0.00021642 3.3 0.00021634 3.3 0.00021644 0 0.00021636 0 0.00021646 3.3 0.00021637999999999998 3.3 0.00021648 0 0.0002164 0 0.0002165 3.3 0.00021642 3.3 0.00021652 0 0.00021643999999999998 0 0.00021653999999999998 3.3 0.00021646 3.3 0.00021656 0 0.00021648 0 0.00021658 3.3 0.0002165 3.3 0.0002166 0 0.00021652 0 0.00021662 3.3 0.00021653999999999998 3.3 0.00021663999999999999 0 0.00021656 0 0.00021666 3.3 0.00021658 3.3 0.00021668 0 0.0002166 0 0.0002167 3.3 0.00021662 3.3 0.00021672 0 0.00021663999999999999 0 0.00021674 3.3 0.00021666 3.3 0.00021676 0 0.00021668 0 0.00021678 3.3 0.00021669999999999998 3.3 0.00021679999999999998 0 0.00021672 0 0.00021682 3.3 0.00021674 3.3 0.00021684 0 0.00021676 0 0.00021686 3.3 0.00021678 3.3 0.00021688 0 0.00021679999999999998 0 0.0002169 3.3 0.00021682 3.3 0.00021692 0 0.00021684 0 0.00021694 3.3 0.00021685999999999998 3.3 0.00021695999999999998 0 0.00021688 0 0.00021698 3.3 0.0002169 3.3 0.000217 0 0.00021692 0 0.00021702 3.3 0.00021694 3.3 0.00021704 0 0.00021695999999999998 0 0.00021705999999999999 3.3 0.00021698 3.3 0.00021708 0 0.000217 0 0.0002171 3.3 0.00021702 3.3 0.00021712 0 0.00021704 0 0.00021714 3.3 0.00021705999999999999 3.3 0.00021716 0 0.00021708 0 0.00021718 3.3 0.0002171 3.3 0.0002172 0 0.00021711999999999998 0 0.00021721999999999998 3.3 0.00021714 3.3 0.00021724 0 0.00021716 0 0.00021726 3.3 0.00021718 3.3 0.00021728 0 0.0002172 0 0.0002173 3.3 0.00021721999999999998 3.3 0.00021731999999999999 0 0.00021724 0 0.00021734 3.3 0.00021726 3.3 0.00021736 0 0.00021727999999999998 0 0.00021737999999999998 3.3 0.0002173 3.3 0.0002174 0 0.00021731999999999999 0 0.00021742 3.3 0.00021734 3.3 0.00021744 0 0.00021736 0 0.00021746 3.3 0.00021737999999999998 3.3 0.00021747999999999998 0 0.0002174 0 0.0002175 3.3 0.00021742 3.3 0.00021752 0 0.00021744 0 0.00021754 3.3 0.00021746 3.3 0.00021756 0 0.00021747999999999998 0 0.00021758 3.3 0.0002175 3.3 0.0002176 0 0.00021752 0 0.00021762 3.3 0.00021753999999999998 3.3 0.00021763999999999998 0 0.00021756 0 0.00021766 3.3 0.00021758 3.3 0.00021768 0 0.0002176 0 0.0002177 3.3 0.00021762 3.3 0.00021772 0 0.00021763999999999998 0 0.00021773999999999999 3.3 0.00021766 3.3 0.00021776 0 0.00021768 0 0.00021778 3.3 0.0002177 3.3 0.0002178 0 0.00021772 0 0.00021782 3.3 0.00021773999999999999 3.3 0.00021784 0 0.00021776 0 0.00021786 3.3 0.00021778 3.3 0.00021788 0 0.00021779999999999998 0 0.00021789999999999998 3.3 0.00021782 3.3 0.00021792 0 0.00021784 0 0.00021794 3.3 0.00021786 3.3 0.00021796 0 0.00021788 0 0.00021798 3.3 0.00021789999999999998 3.3 0.00021799999999999999 0 0.00021792 0 0.00021802 3.3 0.00021794 3.3 0.00021804 0 0.00021795999999999998 0 0.00021805999999999998 3.3 0.00021798 3.3 0.00021808 0 0.00021799999999999999 0 0.0002181 3.3 0.00021802 3.3 0.00021812 0 0.00021804 0 0.00021814 3.3 0.00021805999999999998 3.3 0.00021815999999999998 0 0.00021808 0 0.00021818 3.3 0.0002181 3.3 0.0002182 0 0.00021812 0 0.00021822 3.3 0.00021814 3.3 0.00021824 0 0.00021815999999999998 0 0.00021826 3.3 0.00021818 3.3 0.00021828 0 0.0002182 0 0.0002183 3.3 0.00021821999999999998 3.3 0.00021831999999999998 0 0.00021824 0 0.00021834 3.3 0.00021826 3.3 0.00021836 0 0.00021828 0 0.00021838 3.3 0.0002183 3.3 0.0002184 0 0.00021831999999999998 0 0.00021841999999999999 3.3 0.00021834 3.3 0.00021844 0 0.00021836 0 0.00021846 3.3 0.00021838 3.3 0.00021848 0 0.0002184 0 0.0002185 3.3 0.00021841999999999999 3.3 0.00021852 0 0.00021844 0 0.00021854 3.3 0.00021846 3.3 0.00021856 0 0.00021847999999999998 0 0.00021857999999999998 3.3 0.0002185 3.3 0.0002186 0 0.00021852 0 0.00021862 3.3 0.00021854 3.3 0.00021864 0 0.00021856 0 0.00021866 3.3 0.00021857999999999998 3.3 0.00021868 0 0.0002186 0 0.0002187 3.3 0.00021862 3.3 0.00021872 0 0.00021863999999999998 0 0.00021873999999999998 3.3 0.00021866 3.3 0.00021876 0 0.00021868 0 0.00021878 3.3 0.0002187 3.3 0.0002188 0 0.00021872 0 0.00021882 3.3 0.00021873999999999998 3.3 0.00021883999999999999 0 0.00021876 0 0.00021886 3.3 0.00021878 3.3 0.00021888 0 0.0002188 0 0.0002189 3.3 0.00021882 3.3 0.00021892 0 0.00021883999999999999 0 0.00021894 3.3 0.00021886 3.3 0.00021896 0 0.00021888 0 0.00021898 3.3 0.00021889999999999998 3.3 0.00021899999999999998 0 0.00021892 0 0.00021902 3.3 0.00021894 3.3 0.00021904 0 0.00021896 0 0.00021906 3.3 0.00021898 3.3 0.00021908 0 0.00021899999999999998 0 0.00021909999999999999 3.3 0.00021902 3.3 0.00021912 0 0.00021904 0 0.00021914 3.3 0.00021906 3.3 0.00021916 0 0.00021908 0 0.00021918 3.3 0.00021909999999999999 3.3 0.0002192 0 0.00021912 0 0.00021922 3.3 0.00021914 3.3 0.00021924 0 0.00021915999999999998 0 0.00021925999999999998 3.3 0.00021918 3.3 0.00021928 0 0.0002192 0 0.0002193 3.3 0.00021922 3.3 0.00021932 0 0.00021924 0 0.00021934 3.3 0.00021925999999999998 3.3 0.00021936 0 0.00021928 0 0.00021938 3.3 0.0002193 3.3 0.0002194 0 0.00021931999999999998 0 0.00021941999999999998 3.3 0.00021934 3.3 0.00021944 0 0.00021936 0 0.00021946 3.3 0.00021938 3.3 0.00021948 0 0.0002194 0 0.0002195 3.3 0.00021941999999999998 3.3 0.00021951999999999999 0 0.00021944 0 0.00021954 3.3 0.00021946 3.3 0.00021956 0 0.00021948 0 0.00021958 3.3 0.0002195 3.3 0.0002196 0 0.00021951999999999999 0 0.00021962 3.3 0.00021954 3.3 0.00021964 0 0.00021956 0 0.00021966 3.3 0.00021957999999999998 3.3 0.00021967999999999998 0 0.0002196 0 0.0002197 3.3 0.00021962 3.3 0.00021972 0 0.00021964 0 0.00021974 3.3 0.00021966 3.3 0.00021976 0 0.00021967999999999998 0 0.00021977999999999999 3.3 0.0002197 3.3 0.0002198 0 0.00021972 0 0.00021982 3.3 0.00021973999999999998 3.3 0.00021983999999999998 0 0.00021976 0 0.00021986 3.3 0.00021977999999999999 3.3 0.00021988 0 0.0002198 0 0.0002199 3.3 0.00021982 3.3 0.00021992 0 0.00021983999999999998 0 0.00021993999999999998 3.3 0.00021986 3.3 0.00021996 0 0.00021988 0 0.00021998 3.3 0.0002199 3.3 0.00022 0 0.00021992 0 0.00022002 3.3 0.00021993999999999998 3.3 0.00022004 0 0.00021996 0 0.00022006 3.3 0.00021998 3.3 0.00022008 0 0.00021999999999999998 0 0.00022009999999999998 3.3 0.00022002 3.3 0.00022012 0 0.00022004 0 0.00022014 3.3 0.00022006 3.3 0.00022016 0 0.00022008 0 0.00022018 3.3 0.00022009999999999998 3.3 0.00022019999999999999 0 0.00022012 0 0.00022022 3.3 0.00022014 3.3 0.00022024 0 0.00022016 0 0.00022026 3.3 0.00022018 3.3 0.00022028 0 0.00022019999999999999 0 0.0002203 3.3 0.00022022 3.3 0.00022032 0 0.00022024 0 0.00022034 3.3 0.00022025999999999998 3.3 0.00022035999999999998 0 0.00022028 0 0.00022038 3.3 0.0002203 3.3 0.0002204 0 0.00022032 0 0.00022042 3.3 0.00022034 3.3 0.00022044 0 0.00022035999999999998 0 0.00022046 3.3 0.00022038 3.3 0.00022048 0 0.0002204 0 0.0002205 3.3 0.00022041999999999998 3.3 0.00022051999999999998 0 0.00022044 0 0.00022054 3.3 0.00022046 3.3 0.00022056 0 0.00022048 0 0.00022058 3.3 0.0002205 3.3 0.0002206 0 0.00022051999999999998 0 0.00022061999999999998 3.3 0.00022054 3.3 0.00022064 0 0.00022056 0 0.00022066 3.3 0.00022058 3.3 0.00022068 0 0.0002206 0 0.0002207 3.3 0.00022061999999999998 3.3 0.00022072 0 0.00022064 0 0.00022074 3.3 0.00022066 3.3 0.00022076 0 0.00022067999999999998 0 0.00022077999999999998 3.3 0.0002207 3.3 0.0002208 0 0.00022072 0 0.00022082 3.3 0.00022074 3.3 0.00022084 0 0.00022076 0 0.00022086 3.3 0.00022077999999999998 3.3 0.00022087999999999999 0 0.0002208 0 0.0002209 3.3 0.00022082 3.3 0.00022092 0 0.00022084 0 0.00022094 3.3 0.00022086 3.3 0.00022096 0 0.00022087999999999999 0 0.00022098 3.3 0.0002209 3.3 0.000221 0 0.00022092 0 0.00022102 3.3 0.00022093999999999998 3.3 0.00022103999999999998 0 0.00022096 0 0.00022106 3.3 0.00022098 3.3 0.00022108 0 0.000221 0 0.0002211 3.3 0.00022102 3.3 0.00022112 0 0.00022103999999999998 0 0.00022114 3.3 0.00022106 3.3 0.00022116 0 0.00022108 0 0.00022118 3.3 0.00022109999999999998 3.3 0.00022119999999999998 0 0.00022112 0 0.00022122 3.3 0.00022114 3.3 0.00022124 0 0.00022116 0 0.00022126 3.3 0.00022118 3.3 0.00022128 0 0.00022119999999999998 0 0.00022129999999999999 3.3 0.00022122 3.3 0.00022132 0 0.00022124 0 0.00022134 3.3 0.00022126 3.3 0.00022136 0 0.00022128 0 0.00022138 3.3 0.00022129999999999999 3.3 0.0002214 0 0.00022132 0 0.00022142 3.3 0.00022134 3.3 0.00022144 0 0.00022135999999999998 0 0.00022145999999999998 3.3 0.00022138 3.3 0.00022148 0 0.0002214 0 0.0002215 3.3 0.00022142 3.3 0.00022152 0 0.00022144 0 0.00022154 3.3 0.00022145999999999998 3.3 0.00022155999999999999 0 0.00022148 0 0.00022158 3.3 0.0002215 3.3 0.0002216 0 0.00022151999999999998 0 0.00022161999999999998 3.3 0.00022154 3.3 0.00022164 0 0.00022155999999999999 0 0.00022166 3.3 0.00022158 3.3 0.00022168 0 0.0002216 0 0.0002217 3.3 0.00022161999999999998 3.3 0.00022171999999999998 0 0.00022164 0 0.00022174 3.3 0.00022166 3.3 0.00022176 0 0.00022168 0 0.00022178 3.3 0.0002217 3.3 0.0002218 0 0.00022171999999999998 0 0.00022182 3.3 0.00022174 3.3 0.00022184 0 0.00022176 0 0.00022186 3.3 0.00022177999999999998 3.3 0.00022187999999999998 0 0.0002218 0 0.0002219 3.3 0.00022182 3.3 0.00022192 0 0.00022184 0 0.00022194 3.3 0.00022186 3.3 0.00022196 0 0.00022187999999999998 0 0.00022197999999999999 3.3 0.0002219 3.3 0.000222 0 0.00022192 0 0.00022202 3.3 0.00022194 3.3 0.00022204 0 0.00022196 0 0.00022206 3.3 0.00022197999999999999 3.3 0.00022208 0 0.000222 0 0.0002221 3.3 0.00022202 3.3 0.00022212 0 0.00022203999999999998 0 0.00022213999999999998 3.3 0.00022206 3.3 0.00022216 0 0.00022208 0 0.00022218 3.3 0.0002221 3.3 0.0002222 0 0.00022212 0 0.00022222 3.3 0.00022213999999999998 3.3 0.00022223999999999999 0 0.00022216 0 0.00022226 3.3 0.00022218 3.3 0.00022228 0 0.00022219999999999998 0 0.00022229999999999998 3.3 0.00022222 3.3 0.00022232 0 0.00022223999999999999 0 0.00022234 3.3 0.00022226 3.3 0.00022236 0 0.00022228 0 0.00022238 3.3 0.00022229999999999998 3.3 0.00022239999999999998 0 0.00022232 0 0.00022242 3.3 0.00022234 3.3 0.00022244 0 0.00022236 0 0.00022246 3.3 0.00022238 3.3 0.00022248 0 0.00022239999999999998 0 0.0002225 3.3 0.00022242 3.3 0.00022252 0 0.00022244 0 0.00022254 3.3 0.00022245999999999998 3.3 0.00022255999999999998 0 0.00022248 0 0.00022258 3.3 0.0002225 3.3 0.0002226 0 0.00022252 0 0.00022262 3.3 0.00022254 3.3 0.00022264 0 0.00022255999999999998 0 0.00022265999999999999 3.3 0.00022258 3.3 0.00022268 0 0.0002226 0 0.0002227 3.3 0.00022262 3.3 0.00022272 0 0.00022264 0 0.00022274 3.3 0.00022265999999999999 3.3 0.00022276 0 0.00022268 0 0.00022278 3.3 0.0002227 3.3 0.0002228 0 0.00022271999999999998 0 0.00022281999999999998 3.3 0.00022274 3.3 0.00022284 0 0.00022276 0 0.00022286 3.3 0.00022278 3.3 0.00022288 0 0.0002228 0 0.0002229 3.3 0.00022281999999999998 3.3 0.00022292 0 0.00022284 0 0.00022294 3.3 0.00022286 3.3 0.00022296 0 0.00022287999999999998 0 0.00022297999999999998 3.3 0.0002229 3.3 0.000223 0 0.00022292 0 0.00022302 3.3 0.00022294 3.3 0.00022304 0 0.00022296 0 0.00022306 3.3 0.00022297999999999998 3.3 0.00022307999999999999 0 0.000223 0 0.0002231 3.3 0.00022302 3.3 0.00022312 0 0.00022304 0 0.00022314 3.3 0.00022306 3.3 0.00022316 0 0.00022307999999999999 0 0.00022318 3.3 0.0002231 3.3 0.0002232 0 0.00022312 0 0.00022322 3.3 0.00022313999999999998 3.3 0.00022323999999999998 0 0.00022316 0 0.00022326 3.3 0.00022318 3.3 0.00022328 0 0.0002232 0 0.0002233 3.3 0.00022322 3.3 0.00022332 0 0.00022323999999999998 0 0.00022333999999999999 3.3 0.00022326 3.3 0.00022336 0 0.00022328 0 0.00022338 3.3 0.00022329999999999998 3.3 0.00022339999999999998 0 0.00022332 0 0.00022342 3.3 0.00022333999999999999 3.3 0.00022344 0 0.00022336 0 0.00022346 3.3 0.00022338 3.3 0.00022348 0 0.00022339999999999998 0 0.00022349999999999998 3.3 0.00022342 3.3 0.00022352 0 0.00022344 0 0.00022354 3.3 0.00022346 3.3 0.00022356 0 0.00022348 0 0.00022358 3.3 0.00022349999999999998 3.3 0.0002236 0 0.00022352 0 0.00022362 3.3 0.00022354 3.3 0.00022364 0 0.00022355999999999998 0 0.00022365999999999998 3.3 0.00022358 3.3 0.00022368 0 0.0002236 0 0.0002237 3.3 0.00022362 3.3 0.00022372 0 0.00022364 0 0.00022374 3.3 0.00022365999999999998 3.3 0.00022375999999999999 0 0.00022368 0 0.00022378 3.3 0.0002237 3.3 0.0002238 0 0.00022372 0 0.00022382 3.3 0.00022374 3.3 0.00022384 0 0.00022375999999999999 0 0.00022386 3.3 0.00022378 3.3 0.00022388 0 0.0002238 0 0.0002239 3.3 0.00022381999999999998 3.3 0.00022391999999999998 0 0.00022384 0 0.00022394 3.3 0.00022386 3.3 0.00022396 0 0.00022388 0 0.00022398 3.3 0.0002239 3.3 0.000224 0 0.00022391999999999998 0 0.00022401999999999999 3.3 0.00022394 3.3 0.00022404 0 0.00022396 0 0.00022406 3.3 0.00022397999999999998 3.3 0.00022407999999999998 0 0.000224 0 0.0002241 3.3 0.00022401999999999999 3.3 0.00022412 0 0.00022404 0 0.00022414 3.3 0.00022406 3.3 0.00022416 0 0.00022407999999999998 0 0.00022417999999999998 3.3 0.0002241 3.3 0.0002242 0 0.00022412 0 0.00022422 3.3 0.00022414 3.3 0.00022424 0 0.00022416 0 0.00022426 3.3 0.00022417999999999998 3.3 0.00022428 0 0.0002242 0 0.0002243 3.3 0.00022422 3.3 0.00022432 0 0.00022423999999999998 0 0.00022433999999999998 3.3 0.00022426 3.3 0.00022436 0 0.00022428 0 0.00022438 3.3 0.0002243 3.3 0.0002244 0 0.00022432 0 0.00022442 3.3 0.00022433999999999998 3.3 0.00022443999999999999 0 0.00022436 0 0.00022446 3.3 0.00022438 3.3 0.00022448 0 0.0002244 0 0.0002245 3.3 0.00022442 3.3 0.00022452 0 0.00022443999999999999 0 0.00022454 3.3 0.00022446 3.3 0.00022456 0 0.00022448 0 0.00022458 3.3 0.00022449999999999998 3.3 0.00022459999999999998 0 0.00022452 0 0.00022462 3.3 0.00022454 3.3 0.00022464 0 0.00022456 0 0.00022466 3.3 0.00022458 3.3 0.00022468 0 0.00022459999999999998 0 0.0002247 3.3 0.00022462 3.3 0.00022472 0 0.00022464 0 0.00022474 3.3 0.00022465999999999998 3.3 0.00022475999999999998 0 0.00022468 0 0.00022478 3.3 0.0002247 3.3 0.0002248 0 0.00022472 0 0.00022482 3.3 0.00022474 3.3 0.00022484 0 0.00022475999999999998 0 0.00022485999999999999 3.3 0.00022478 3.3 0.00022488 0 0.0002248 0 0.0002249 3.3 0.00022482 3.3 0.00022492 0 0.00022484 0 0.00022494 3.3 0.00022485999999999999 3.3 0.00022496 0 0.00022488 0 0.00022498 3.3 0.0002249 3.3 0.000225 0 0.00022491999999999998 0 0.00022501999999999998 3.3 0.00022494 3.3 0.00022504 0 0.00022496 0 0.00022506 3.3 0.00022498 3.3 0.00022508 0 0.000225 0 0.0002251 3.3 0.00022501999999999998 3.3 0.00022511999999999999 0 0.00022504 0 0.00022514 3.3 0.00022506 3.3 0.00022516 0 0.00022507999999999998 0 0.00022517999999999998 3.3 0.0002251 3.3 0.0002252 0 0.00022511999999999999 0 0.00022522 3.3 0.00022514 3.3 0.00022524 0 0.00022516 0 0.00022526 3.3 0.00022517999999999998 3.3 0.00022527999999999998 0 0.0002252 0 0.0002253 3.3 0.00022522 3.3 0.00022532 0 0.00022524 0 0.00022534 3.3 0.00022526 3.3 0.00022536 0 0.00022527999999999998 0 0.00022538 3.3 0.0002253 3.3 0.0002254 0 0.00022532 0 0.00022542 3.3 0.00022533999999999998 3.3 0.00022543999999999998 0 0.00022536 0 0.00022546 3.3 0.00022538 3.3 0.00022548 0 0.0002254 0 0.0002255 3.3 0.00022542 3.3 0.00022552 0 0.00022543999999999998 0 0.00022553999999999999 3.3 0.00022546 3.3 0.00022556 0 0.00022548 0 0.00022558 3.3 0.0002255 3.3 0.0002256 0 0.00022552 0 0.00022562 3.3 0.00022553999999999999 3.3 0.00022564 0 0.00022556 0 0.00022566 3.3 0.00022558 3.3 0.00022568 0 0.00022559999999999998 0 0.00022569999999999998 3.3 0.00022562 3.3 0.00022572 0 0.00022564 0 0.00022574 3.3 0.00022566 3.3 0.00022576 0 0.00022568 0 0.00022578 3.3 0.00022569999999999998 3.3 0.00022579999999999999 0 0.00022572 0 0.00022582 3.3 0.00022574 3.3 0.00022584 0 0.00022575999999999998 0 0.00022585999999999998 3.3 0.00022578 3.3 0.00022588 0 0.00022579999999999999 0 0.0002259 3.3 0.00022582 3.3 0.00022592 0 0.00022584 0 0.00022594 3.3 0.00022585999999999998 3.3 0.00022595999999999998 0 0.00022588 0 0.00022598 3.3 0.0002259 3.3 0.000226 0 0.00022592 0 0.00022602 3.3 0.00022594 3.3 0.00022604 0 0.00022595999999999998 0 0.00022606 3.3 0.00022598 3.3 0.00022608 0 0.000226 0 0.0002261 3.3 0.00022601999999999998 3.3 0.00022611999999999998 0 0.00022604 0 0.00022614 3.3 0.00022606 3.3 0.00022616 0 0.00022608 0 0.00022618 3.3 0.0002261 3.3 0.0002262 0 0.00022611999999999998 0 0.00022621999999999999 3.3 0.00022614 3.3 0.00022624 0 0.00022616 0 0.00022626 3.3 0.00022618 3.3 0.00022628 0 0.0002262 0 0.0002263 3.3 0.00022621999999999999 3.3 0.00022632 0 0.00022624 0 0.00022634 3.3 0.00022626 3.3 0.00022636 0 0.00022627999999999998 0 0.00022637999999999998 3.3 0.0002263 3.3 0.0002264 0 0.00022632 0 0.00022642 3.3 0.00022634 3.3 0.00022644 0 0.00022636 0 0.00022646 3.3 0.00022637999999999998 3.3 0.00022648 0 0.0002264 0 0.0002265 3.3 0.00022642 3.3 0.00022652 0 0.00022643999999999998 0 0.00022653999999999998 3.3 0.00022646 3.3 0.00022656 0 0.00022648 0 0.00022658 3.3 0.0002265 3.3 0.0002266 0 0.00022652 0 0.00022662 3.3 0.00022653999999999998 3.3 0.00022663999999999998 0 0.00022656 0 0.00022666 3.3 0.00022658 3.3 0.00022668 0 0.0002266 0 0.0002267 3.3 0.00022662 3.3 0.00022672 0 0.00022663999999999998 0 0.00022674 3.3 0.00022666 3.3 0.00022676 0 0.00022668 0 0.00022678 3.3 0.00022669999999999998 3.3 0.00022679999999999998 0 0.00022672 0 0.00022682 3.3 0.00022674 3.3 0.00022684 0 0.00022676 0 0.00022686 3.3 0.00022678 3.3 0.00022688 0 0.00022679999999999998 0 0.00022689999999999999 3.3 0.00022682 3.3 0.00022692 0 0.00022684 0 0.00022694 3.3 0.00022686 3.3 0.00022696 0 0.00022688 0 0.00022698 3.3 0.00022689999999999999 3.3 0.000227 0 0.00022692 0 0.00022702 3.3 0.00022694 3.3 0.00022704 0 0.00022695999999999998 0 0.00022705999999999998 3.3 0.00022698 3.3 0.00022708 0 0.000227 0 0.0002271 3.3 0.00022702 3.3 0.00022712 0 0.00022704 0 0.00022714 3.3 0.00022705999999999998 3.3 0.00022716 0 0.00022708 0 0.00022718 3.3 0.0002271 3.3 0.0002272 0 0.00022711999999999998 0 0.00022721999999999998 3.3 0.00022714 3.3 0.00022724 0 0.00022716 0 0.00022726 3.3 0.00022718 3.3 0.00022728 0 0.0002272 0 0.0002273 3.3 0.00022721999999999998 3.3 0.00022731999999999999 0 0.00022724 0 0.00022734 3.3 0.00022726 3.3 0.00022736 0 0.00022728 0 0.00022738 3.3 0.0002273 3.3 0.0002274 0 0.00022731999999999999 0 0.00022742 3.3 0.00022734 3.3 0.00022744 0 0.00022736 0 0.00022746 3.3 0.00022737999999999998 3.3 0.00022747999999999998 0 0.0002274 0 0.0002275 3.3 0.00022742 3.3 0.00022752 0 0.00022744 0 0.00022754 3.3 0.00022746 3.3 0.00022756 0 0.00022747999999999998 0 0.00022757999999999999 3.3 0.0002275 3.3 0.0002276 0 0.00022752 0 0.00022762 3.3 0.00022753999999999998 3.3 0.00022763999999999998 0 0.00022756 0 0.00022766 3.3 0.00022757999999999999 3.3 0.00022768 0 0.0002276 0 0.0002277 3.3 0.00022762 3.3 0.00022772 0 0.00022763999999999998 0 0.00022773999999999998 3.3 0.00022766 3.3 0.00022776 0 0.00022768 0 0.00022778 3.3 0.0002277 3.3 0.0002278 0 0.00022772 0 0.00022782 3.3 0.00022773999999999998 3.3 0.00022784 0 0.00022776 0 0.00022786 3.3 0.00022778 3.3 0.00022788 0 0.00022779999999999998 0 0.00022789999999999998 3.3 0.00022782 3.3 0.00022792 0 0.00022784 0 0.00022794 3.3 0.00022786 3.3 0.00022796 0 0.00022788 0 0.00022798 3.3 0.00022789999999999998 3.3 0.00022799999999999999 0 0.00022792 0 0.00022802 3.3 0.00022794 3.3 0.00022804 0 0.00022796 0 0.00022806 3.3 0.00022798 3.3 0.00022808 0 0.00022799999999999999 0 0.0002281 3.3 0.00022802 3.3 0.00022812 0 0.00022804 0 0.00022814 3.3 0.00022805999999999998 3.3 0.00022815999999999998 0 0.00022808 0 0.00022818 3.3 0.0002281 3.3 0.0002282 0 0.00022812 0 0.00022822 3.3 0.00022814 3.3 0.00022824 0 0.00022815999999999998 0 0.00022825999999999999 3.3 0.00022818 3.3 0.00022828 0 0.0002282 0 0.0002283 3.3 0.00022821999999999998 3.3 0.00022831999999999998 0 0.00022824 0 0.00022834 3.3 0.00022825999999999999 3.3 0.00022836 0 0.00022828 0 0.00022838 3.3 0.0002283 3.3 0.0002284 0 0.00022831999999999998 0 0.00022841999999999998 3.3 0.00022834 3.3 0.00022844 0 0.00022836 0 0.00022846 3.3 0.00022838 3.3 0.00022848 0 0.0002284 0 0.0002285 3.3 0.00022841999999999998 3.3 0.00022852 0 0.00022844 0 0.00022854 3.3 0.00022846 3.3 0.00022856 0 0.00022847999999999998 0 0.00022857999999999998 3.3 0.0002285 3.3 0.0002286 0 0.00022852 0 0.00022862 3.3 0.00022854 3.3 0.00022864 0 0.00022856 0 0.00022866 3.3 0.00022857999999999998 3.3 0.00022867999999999999 0 0.0002286 0 0.0002287 3.3 0.00022862 3.3 0.00022872 0 0.00022864 0 0.00022874 3.3 0.00022866 3.3 0.00022876 0 0.00022867999999999999 0 0.00022878 3.3 0.0002287 3.3 0.0002288 0 0.00022872 0 0.00022882 3.3 0.00022873999999999998 3.3 0.00022883999999999998 0 0.00022876 0 0.00022886 3.3 0.00022878 3.3 0.00022888 0 0.0002288 0 0.0002289 3.3 0.00022882 3.3 0.00022892 0 0.00022883999999999998 0 0.00022894 3.3 0.00022886 3.3 0.00022896 0 0.00022888 0 0.00022898 3.3 0.00022889999999999998 3.3 0.00022899999999999998 0 0.00022892 0 0.00022902 3.3 0.00022894 3.3 0.00022904 0 0.00022896 0 0.00022906 3.3 0.00022898 3.3 0.00022908 0 0.00022899999999999998 0 0.00022909999999999999 3.3 0.00022902 3.3 0.00022912 0 0.00022904 0 0.00022914 3.3 0.00022906 3.3 0.00022916 0 0.00022908 0 0.00022918 3.3 0.00022909999999999999 3.3 0.0002292 0 0.00022912 0 0.00022922 3.3 0.00022914 3.3 0.00022924 0 0.00022915999999999998 0 0.00022925999999999998 3.3 0.00022918 3.3 0.00022928 0 0.0002292 0 0.0002293 3.3 0.00022922 3.3 0.00022932 0 0.00022924 0 0.00022934 3.3 0.00022925999999999998 3.3 0.00022935999999999999 0 0.00022928 0 0.00022938 3.3 0.0002293 3.3 0.0002294 0 0.00022931999999999998 0 0.00022941999999999998 3.3 0.00022934 3.3 0.00022944 0 0.00022935999999999999 0 0.00022946 3.3 0.00022938 3.3 0.00022948 0 0.0002294 0 0.0002295 3.3 0.00022941999999999998 3.3 0.00022951999999999998 0 0.00022944 0 0.00022954 3.3 0.00022946 3.3 0.00022956 0 0.00022948 0 0.00022958 3.3 0.0002295 3.3 0.0002296 0 0.00022951999999999998 0 0.00022962 3.3 0.00022954 3.3 0.00022964 0 0.00022956 0 0.00022966 3.3 0.00022957999999999998 3.3 0.00022967999999999998 0 0.0002296 0 0.0002297 3.3 0.00022962 3.3 0.00022972 0 0.00022964 0 0.00022974 3.3 0.00022966 3.3 0.00022976 0 0.00022967999999999998 0 0.00022977999999999999 3.3 0.0002297 3.3 0.0002298 0 0.00022972 0 0.00022982 3.3 0.00022974 3.3 0.00022984 0 0.00022976 0 0.00022986 3.3 0.00022977999999999999 3.3 0.00022988 0 0.0002298 0 0.0002299 3.3 0.00022982 3.3 0.00022992 0 0.00022983999999999998 0 0.00022993999999999998 3.3 0.00022986 3.3 0.00022996 0 0.00022988 0 0.00022998 3.3 0.0002299 3.3 0.00023 0 0.00022992 0 0.00023002 3.3 0.00022993999999999998 3.3 0.00023003999999999999 0 0.00022996 0 0.00023006 3.3 0.00022998 3.3 0.00023008 0 0.00022999999999999998 0 0.00023009999999999998 3.3 0.00023002 3.3 0.00023012 0 0.00023003999999999999 0 0.00023014 3.3 0.00023006 3.3 0.00023016 0 0.00023008 0 0.00023018 3.3 0.00023009999999999998 3.3 0.00023019999999999998 0 0.00023012 0 0.00023022 3.3 0.00023014 3.3 0.00023024 0 0.00023016 0 0.00023026 3.3 0.00023018 3.3 0.00023028 0 0.00023019999999999998 0 0.0002303 3.3 0.00023022 3.3 0.00023032 0 0.00023024 0 0.00023034 3.3 0.00023025999999999998 3.3 0.00023035999999999998 0 0.00023028 0 0.00023038 3.3 0.0002303 3.3 0.0002304 0 0.00023032 0 0.00023042 3.3 0.00023034 3.3 0.00023044 0 0.00023035999999999998 0 0.00023045999999999999 3.3 0.00023038 3.3 0.00023048 0 0.0002304 0 0.0002305 3.3 0.00023042 3.3 0.00023052 0 0.00023044 0 0.00023054 3.3 0.00023045999999999999 3.3 0.00023056 0 0.00023048 0 0.00023058 3.3 0.0002305 3.3 0.0002306 0 0.00023051999999999998 0 0.00023061999999999998 3.3 0.00023054 3.3 0.00023064 0 0.00023056 0 0.00023066 3.3 0.00023058 3.3 0.00023068 0 0.0002306 0 0.0002307 3.3 0.00023061999999999998 3.3 0.00023072 0 0.00023064 0 0.00023074 3.3 0.00023066 3.3 0.00023076 0 0.00023067999999999998 0 0.00023077999999999998 3.3 0.0002307 3.3 0.0002308 0 0.00023072 0 0.00023082 3.3 0.00023074 3.3 0.00023084 0 0.00023076 0 0.00023086 3.3 0.00023077999999999998 3.3 0.00023087999999999998 0 0.0002308 0 0.0002309 3.3 0.00023082 3.3 0.00023092 0 0.00023084 0 0.00023094 3.3 0.00023086 3.3 0.00023096 0 0.00023087999999999998 0 0.00023098 3.3 0.0002309 3.3 0.000231 0 0.00023092 0 0.00023102 3.3 0.00023093999999999998 3.3 0.00023103999999999998 0 0.00023096 0 0.00023106 3.3 0.00023098 3.3 0.00023108 0 0.000231 0 0.0002311 3.3 0.00023102 3.3 0.00023112 0 0.00023103999999999998 0 0.00023113999999999999 3.3 0.00023106 3.3 0.00023116 0 0.00023108 0 0.00023118 3.3 0.00023109999999999998 3.3 0.00023119999999999998 0 0.00023112 0 0.00023122 3.3 0.00023113999999999999 3.3 0.00023124 0 0.00023116 0 0.00023126 3.3 0.00023118 3.3 0.00023128 0 0.00023119999999999998 0 0.00023129999999999998 3.3 0.00023122 3.3 0.00023132 0 0.00023124 0 0.00023134 3.3 0.00023126 3.3 0.00023136 0 0.00023128 0 0.00023138 3.3 0.00023129999999999998 3.3 0.0002314 0 0.00023132 0 0.00023142 3.3 0.00023134 3.3 0.00023144 0 0.00023135999999999998 0 0.00023145999999999998 3.3 0.00023138 3.3 0.00023148 0 0.0002314 0 0.0002315 3.3 0.00023142 3.3 0.00023152 0 0.00023144 0 0.00023154 3.3 0.00023145999999999998 3.3 0.00023155999999999999 0 0.00023148 0 0.00023158 3.3 0.0002315 3.3 0.0002316 0 0.00023152 0 0.00023162 3.3 0.00023154 3.3 0.00023164 0 0.00023155999999999999 0 0.00023166 3.3 0.00023158 3.3 0.00023168 0 0.0002316 0 0.0002317 3.3 0.00023161999999999998 3.3 0.00023171999999999998 0 0.00023164 0 0.00023174 3.3 0.00023166 3.3 0.00023176 0 0.00023168 0 0.00023178 3.3 0.0002317 3.3 0.0002318 0 0.00023171999999999998 0 0.00023181999999999999 3.3 0.00023174 3.3 0.00023184 0 0.00023176 0 0.00023186 3.3 0.00023177999999999998 3.3 0.00023187999999999998 0 0.0002318 0 0.0002319 3.3 0.00023181999999999999 3.3 0.00023192 0 0.00023184 0 0.00023194 3.3 0.00023186 3.3 0.00023196 0 0.00023187999999999998 0 0.00023197999999999998 3.3 0.0002319 3.3 0.000232 0 0.00023192 0 0.00023202 3.3 0.00023194 3.3 0.00023204 0 0.00023196 0 0.00023206 3.3 0.00023197999999999998 3.3 0.00023208 0 0.000232 0 0.0002321 3.3 0.00023202 3.3 0.00023212 0 0.00023203999999999998 0 0.00023213999999999998 3.3 0.00023206 3.3 0.00023216 0 0.00023208 0 0.00023218 3.3 0.0002321 3.3 0.0002322 0 0.00023212 0 0.00023222 3.3 0.00023213999999999998 3.3 0.00023223999999999999 0 0.00023216 0 0.00023226 3.3 0.00023218 3.3 0.00023228 0 0.0002322 0 0.0002323 3.3 0.00023222 3.3 0.00023232 0 0.00023223999999999999 0 0.00023234 3.3 0.00023226 3.3 0.00023236 0 0.00023228 0 0.00023238 3.3 0.00023229999999999998 3.3 0.00023239999999999998 0 0.00023232 0 0.00023242 3.3 0.00023234 3.3 0.00023244 0 0.00023236 0 0.00023246 3.3 0.00023238 3.3 0.00023248 0 0.00023239999999999998 0 0.00023249999999999999 3.3 0.00023242 3.3 0.00023252 0 0.00023244 0 0.00023254 3.3 0.00023245999999999998 3.3 0.00023255999999999998 0 0.00023248 0 0.00023258 3.3 0.00023249999999999999 3.3 0.0002326 0 0.00023252 0 0.00023262 3.3 0.00023254 3.3 0.00023264 0 0.00023255999999999998 0 0.00023265999999999998 3.3 0.00023258 3.3 0.00023268 0 0.0002326 0 0.0002327 3.3 0.00023262 3.3 0.00023272 0 0.00023264 0 0.00023274 3.3 0.00023265999999999998 3.3 0.00023276 0 0.00023268 0 0.00023278 3.3 0.0002327 3.3 0.0002328 0 0.00023271999999999998 0 0.00023281999999999998 3.3 0.00023274 3.3 0.00023284 0 0.00023276 0 0.00023286 3.3 0.00023278 3.3 0.00023288 0 0.0002328 0 0.0002329 3.3 0.00023281999999999998 3.3 0.00023291999999999999 0 0.00023284 0 0.00023294 3.3 0.00023286 3.3 0.00023296 0 0.00023287999999999998 0 0.00023297999999999998 3.3 0.0002329 3.3 0.000233 0 0.00023291999999999999 0 0.00023302 3.3 0.00023294 3.3 0.00023304 0 0.00023296 0 0.00023306 3.3 0.00023297999999999998 3.3 0.00023307999999999998 0 0.000233 0 0.0002331 3.3 0.00023302 3.3 0.00023312 0 0.00023304 0 0.00023314 3.3 0.00023306 3.3 0.00023316 0 0.00023307999999999998 0 0.00023318 3.3 0.0002331 3.3 0.0002332 0 0.00023312 0 0.00023322 3.3 0.00023313999999999998 3.3 0.00023323999999999998 0 0.00023316 0 0.00023326 3.3 0.00023318 3.3 0.00023328 0 0.0002332 0 0.0002333 3.3 0.00023322 3.3 0.00023332 0 0.00023323999999999998 0 0.00023333999999999999 3.3 0.00023326 3.3 0.00023336 0 0.00023328 0 0.00023338 3.3 0.0002333 3.3 0.0002334 0 0.00023332 0 0.00023342 3.3 0.00023333999999999999 3.3 0.00023344 0 0.00023336 0 0.00023346 3.3 0.00023338 3.3 0.00023348 0 0.00023339999999999998 0 0.00023349999999999998 3.3 0.00023342 3.3 0.00023352 0 0.00023344 0 0.00023354 3.3 0.00023346 3.3 0.00023356 0 0.00023348 0 0.00023358 3.3 0.00023349999999999998 3.3 0.00023359999999999999 0 0.00023352 0 0.00023362 3.3 0.00023354 3.3 0.00023364 0 0.00023355999999999998 0 0.00023365999999999998 3.3 0.00023358 3.3 0.00023368 0 0.00023359999999999999 0 0.0002337 3.3 0.00023362 3.3 0.00023372 0 0.00023364 0 0.00023374 3.3 0.00023365999999999998 3.3 0.00023375999999999998 0 0.00023368 0 0.00023378 3.3 0.0002337 3.3 0.0002338 0 0.00023372 0 0.00023382 3.3 0.00023374 3.3 0.00023384 0 0.00023375999999999998 0 0.00023386 3.3 0.00023378 3.3 0.00023388 0 0.0002338 0 0.0002339 3.3 0.00023381999999999998 3.3 0.00023391999999999998 0 0.00023384 0 0.00023394 3.3 0.00023386 3.3 0.00023396 0 0.00023388 0 0.00023398 3.3 0.0002339 3.3 0.000234 0 0.00023391999999999998 0 0.00023401999999999999 3.3 0.00023394 3.3 0.00023404 0 0.00023396 0 0.00023406 3.3 0.00023398 3.3 0.00023408 0 0.000234 0 0.0002341 3.3 0.00023401999999999999 3.3 0.00023412 0 0.00023404 0 0.00023414 3.3 0.00023406 3.3 0.00023416 0 0.00023407999999999998 0 0.00023417999999999998 3.3 0.0002341 3.3 0.0002342 0 0.00023412 0 0.00023422 3.3 0.00023414 3.3 0.00023424 0 0.00023416 0 0.00023426 3.3 0.00023417999999999998 3.3 0.00023427999999999999 0 0.0002342 0 0.0002343 3.3 0.00023422 3.3 0.00023432 0 0.00023423999999999998 0 0.00023433999999999998 3.3 0.00023426 3.3 0.00023436 0 0.00023427999999999999 0 0.00023438 3.3 0.0002343 3.3 0.0002344 0 0.00023432 0 0.00023442 3.3 0.00023433999999999998 3.3 0.00023443999999999998 0 0.00023436 0 0.00023446 3.3 0.00023438 3.3 0.00023448 0 0.0002344 0 0.0002345 3.3 0.00023442 3.3 0.00023452 0 0.00023443999999999998 0 0.00023454 3.3 0.00023446 3.3 0.00023456 0 0.00023448 0 0.00023458 3.3 0.00023449999999999998 3.3 0.00023459999999999998 0 0.00023452 0 0.00023462 3.3 0.00023454 3.3 0.00023464 0 0.00023456 0 0.00023466 3.3 0.00023458 3.3 0.00023468 0 0.00023459999999999998 0 0.00023469999999999999 3.3 0.00023462 3.3 0.00023472 0 0.00023464 0 0.00023474 3.3 0.00023466 3.3 0.00023476 0 0.00023468 0 0.00023478 3.3 0.00023469999999999999 3.3 0.0002348 0 0.00023472 0 0.00023482 3.3 0.00023474 3.3 0.00023484 0 0.00023475999999999998 0 0.00023485999999999998 3.3 0.00023478 3.3 0.00023488 0 0.0002348 0 0.0002349 3.3 0.00023482 3.3 0.00023492 0 0.00023484 0 0.00023494 3.3 0.00023485999999999998 3.3 0.00023496 0 0.00023488 0 0.00023498 3.3 0.0002349 3.3 0.000235 0 0.00023491999999999998 0 0.00023501999999999998 3.3 0.00023494 3.3 0.00023504 0 0.00023496 0 0.00023506 3.3 0.00023498 3.3 0.00023508 0 0.000235 0 0.0002351 3.3 0.00023501999999999998 3.3 0.00023511999999999999 0 0.00023504 0 0.00023514 3.3 0.00023506 3.3 0.00023516 0 0.00023508 0 0.00023518 3.3 0.0002351 3.3 0.0002352 0 0.00023511999999999999 0 0.00023522 3.3 0.00023514 3.3 0.00023524 0 0.00023516 0 0.00023526 3.3 0.00023517999999999998 3.3 0.00023527999999999998 0 0.0002352 0 0.0002353 3.3 0.00023522 3.3 0.00023532 0 0.00023524 0 0.00023534 3.3 0.00023526 3.3 0.00023536 0 0.00023527999999999998 0 0.00023537999999999999 3.3 0.0002353 3.3 0.0002354 0 0.00023532 0 0.00023542 3.3 0.00023533999999999998 3.3 0.00023543999999999998 0 0.00023536 0 0.00023546 3.3 0.00023537999999999999 3.3 0.00023548 0 0.0002354 0 0.0002355 3.3 0.00023542 3.3 0.00023552 0 0.00023543999999999998 0 0.00023553999999999998 3.3 0.00023546 3.3 0.00023556 0 0.00023548 0 0.00023558 3.3 0.0002355 3.3 0.0002356 0 0.00023552 0 0.00023562 3.3 0.00023553999999999998 3.3 0.00023564 0 0.00023556 0 0.00023566 3.3 0.00023558 3.3 0.00023568 0 0.00023559999999999998 0 0.00023569999999999998 3.3 0.00023562 3.3 0.00023572 0 0.00023564 0 0.00023574 3.3 0.00023566 3.3 0.00023576 0 0.00023568 0 0.00023578 3.3 0.00023569999999999998 3.3 0.00023579999999999999 0 0.00023572 0 0.00023582 3.3 0.00023574 3.3 0.00023584 0 0.00023576 0 0.00023586 3.3 0.00023578 3.3 0.00023588 0 0.00023579999999999999 0 0.0002359 3.3 0.00023582 3.3 0.00023592 0 0.00023584 0 0.00023594 3.3 0.00023585999999999998 3.3 0.00023595999999999998 0 0.00023588 0 0.00023598 3.3 0.0002359 3.3 0.000236 0 0.00023592 0 0.00023602 3.3 0.00023594 3.3 0.00023604 0 0.00023595999999999998 0 0.00023605999999999999 3.3 0.00023598 3.3 0.00023608 0 0.000236 0 0.0002361 3.3 0.00023601999999999998 3.3 0.00023611999999999998 0 0.00023604 0 0.00023614 3.3 0.00023605999999999999 3.3 0.00023616 0 0.00023608 0 0.00023618 3.3 0.0002361 3.3 0.0002362 0 0.00023611999999999998 0 0.00023621999999999998 3.3 0.00023614 3.3 0.00023624 0 0.00023616 0 0.00023626 3.3 0.00023618 3.3 0.00023628 0 0.0002362 0 0.0002363 3.3 0.00023621999999999998 3.3 0.00023632 0 0.00023624 0 0.00023634 3.3 0.00023626 3.3 0.00023636 0 0.00023627999999999998 0 0.00023637999999999998 3.3 0.0002363 3.3 0.0002364 0 0.00023632 0 0.00023642 3.3 0.00023634 3.3 0.00023644 0 0.00023636 0 0.00023646 3.3 0.00023637999999999998 3.3 0.00023647999999999999 0 0.0002364 0 0.0002365 3.3 0.00023642 3.3 0.00023652 0 0.00023644 0 0.00023654 3.3 0.00023646 3.3 0.00023656 0 0.00023647999999999999 0 0.00023658 3.3 0.0002365 3.3 0.0002366 0 0.00023652 0 0.00023662 3.3 0.00023653999999999998 3.3 0.00023663999999999998 0 0.00023656 0 0.00023666 3.3 0.00023658 3.3 0.00023668 0 0.0002366 0 0.0002367 3.3 0.00023662 3.3 0.00023672 0 0.00023663999999999998 0 0.00023674 3.3 0.00023666 3.3 0.00023676 0 0.00023668 0 0.00023678 3.3 0.00023669999999999998 3.3 0.00023679999999999998 0 0.00023672 0 0.00023682 3.3 0.00023674 3.3 0.00023684 0 0.00023676 0 0.00023686 3.3 0.00023678 3.3 0.00023688 0 0.00023679999999999998 0 0.00023689999999999998 3.3 0.00023682 3.3 0.00023692 0 0.00023684 0 0.00023694 3.3 0.00023686 3.3 0.00023696 0 0.00023688 0 0.00023698 3.3 0.00023689999999999998 3.3 0.000237 0 0.00023692 0 0.00023702 3.3 0.00023694 3.3 0.00023704 0 0.00023695999999999998 0 0.00023705999999999998 3.3 0.00023698 3.3 0.00023708 0 0.000237 0 0.0002371 3.3 0.00023702 3.3 0.00023712 0 0.00023704 0 0.00023714 3.3 0.00023705999999999998 3.3 0.00023715999999999999 0 0.00023708 0 0.00023718 3.3 0.0002371 3.3 0.0002372 0 0.00023711999999999998 0 0.00023721999999999998 3.3 0.00023714 3.3 0.00023724 0 0.00023715999999999999 0 0.00023726 3.3 0.00023718 3.3 0.00023728 0 0.0002372 0 0.0002373 3.3 0.00023721999999999998 3.3 0.00023731999999999998 0 0.00023724 0 0.00023734 3.3 0.00023726 3.3 0.00023736 0 0.00023728 0 0.00023738 3.3 0.0002373 3.3 0.0002374 0 0.00023731999999999998 0 0.00023742 3.3 0.00023734 3.3 0.00023744 0 0.00023736 0 0.00023746 3.3 0.00023737999999999998 3.3 0.00023747999999999998 0 0.0002374 0 0.0002375 3.3 0.00023742 3.3 0.00023752 0 0.00023744 0 0.00023754 3.3 0.00023746 3.3 0.00023756 0 0.00023747999999999998 0 0.00023757999999999999 3.3 0.0002375 3.3 0.0002376 0 0.00023752 0 0.00023762 3.3 0.00023754 3.3 0.00023764 0 0.00023756 0 0.00023766 3.3 0.00023757999999999999 3.3 0.00023768 0 0.0002376 0 0.0002377 3.3 0.00023762 3.3 0.00023772 0 0.00023763999999999998 0 0.00023773999999999998 3.3 0.00023766 3.3 0.00023776 0 0.00023768 0 0.00023778 3.3 0.0002377 3.3 0.0002378 0 0.00023772 0 0.00023782 3.3 0.00023773999999999998 3.3 0.00023783999999999999 0 0.00023776 0 0.00023786 3.3 0.00023778 3.3 0.00023788 0 0.00023779999999999998 0 0.00023789999999999998 3.3 0.00023782 3.3 0.00023792 0 0.00023783999999999999 0 0.00023794 3.3 0.00023786 3.3 0.00023796 0 0.00023788 0 0.00023798 3.3 0.00023789999999999998 3.3 0.00023799999999999998 0 0.00023792 0 0.00023802 3.3 0.00023794 3.3 0.00023804 0 0.00023796 0 0.00023806 3.3 0.00023798 3.3 0.00023808 0 0.00023799999999999998 0 0.0002381 3.3 0.00023802 3.3 0.00023812 0 0.00023804 0 0.00023814 3.3 0.00023805999999999998 3.3 0.00023815999999999998 0 0.00023808 0 0.00023818 3.3 0.0002381 3.3 0.0002382 0 0.00023812 0 0.00023822 3.3 0.00023814 3.3 0.00023824 0 0.00023815999999999998 0 0.00023825999999999999 3.3 0.00023818 3.3 0.00023828 0 0.0002382 0 0.0002383 3.3 0.00023822 3.3 0.00023832 0 0.00023824 0 0.00023834 3.3 0.00023825999999999999 3.3 0.00023836 0 0.00023828 0 0.00023838 3.3 0.0002383 3.3 0.0002384 0 0.00023831999999999998 0 0.00023841999999999998 3.3 0.00023834 3.3 0.00023844 0 0.00023836 0 0.00023846 3.3 0.00023838 3.3 0.00023848 0 0.0002384 0 0.0002385 3.3 0.00023841999999999998 3.3 0.00023851999999999999 0 0.00023844 0 0.00023854 3.3 0.00023846 3.3 0.00023856 0 0.00023847999999999998 0 0.00023857999999999998 3.3 0.0002385 3.3 0.0002386 0 0.00023851999999999999 0 0.00023862 3.3 0.00023854 3.3 0.00023864 0 0.00023856 0 0.00023866 3.3 0.00023857999999999998 3.3 0.00023867999999999998 0 0.0002386 0 0.0002387 3.3 0.00023862 3.3 0.00023872 0 0.00023864 0 0.00023874 3.3 0.00023866 3.3 0.00023876 0 0.00023867999999999998 0 0.00023878 3.3 0.0002387 3.3 0.0002388 0 0.00023872 0 0.00023882 3.3 0.00023873999999999998 3.3 0.00023883999999999998 0 0.00023876 0 0.00023886 3.3 0.00023878 3.3 0.00023888 0 0.0002388 0 0.0002389 3.3 0.00023882 3.3 0.00023892 0 0.00023883999999999998 0 0.00023893999999999999 3.3 0.00023886 3.3 0.00023896 0 0.00023888 0 0.00023898 3.3 0.00023889999999999998 3.3 0.00023899999999999998 0 0.00023892 0 0.00023902 3.3 0.00023893999999999999 3.3 0.00023904 0 0.00023896 0 0.00023906 3.3 0.00023898 3.3 0.00023908 0 0.00023899999999999998 0 0.00023909999999999998 3.3 0.00023902 3.3 0.00023912 0 0.00023904 0 0.00023914 3.3 0.00023906 3.3 0.00023916 0 0.00023908 0 0.00023918 3.3 0.00023909999999999998 3.3 0.0002392 0 0.00023912 0 0.00023922 3.3 0.00023914 3.3 0.00023924 0 0.00023915999999999998 0 0.00023925999999999998 3.3 0.00023918 3.3 0.00023928 0 0.0002392 0 0.0002393 3.3 0.00023922 3.3 0.00023932 0 0.00023924 0 0.00023934 3.3 0.00023925999999999998 3.3 0.00023935999999999999 0 0.00023928 0 0.00023938 3.3 0.0002393 3.3 0.0002394 0 0.00023932 0 0.00023942 3.3 0.00023934 3.3 0.00023944 0 0.00023935999999999999 0 0.00023946 3.3 0.00023938 3.3 0.00023948 0 0.0002394 0 0.0002395 3.3 0.00023941999999999998 3.3 0.00023951999999999998 0 0.00023944 0 0.00023954 3.3 0.00023946 3.3 0.00023956 0 0.00023948 0 0.00023958 3.3 0.0002395 3.3 0.0002396 0 0.00023951999999999998 0 0.00023961999999999999 3.3 0.00023954 3.3 0.00023964 0 0.00023956 0 0.00023966 3.3 0.00023957999999999998 3.3 0.00023967999999999998 0 0.0002396 0 0.0002397 3.3 0.00023961999999999999 3.3 0.00023972 0 0.00023964 0 0.00023974 3.3 0.00023966 3.3 0.00023976 0 0.00023967999999999998 0 0.00023977999999999998 3.3 0.0002397 3.3 0.0002398 0 0.00023972 0 0.00023982 3.3 0.00023974 3.3 0.00023984 0 0.00023976 0 0.00023986 3.3 0.00023977999999999998 3.3 0.00023988 0 0.0002398 0 0.0002399 3.3 0.00023982 3.3 0.00023992 0 0.00023983999999999998 0 0.00023993999999999998 3.3 0.00023986 3.3 0.00023996 0 0.00023988 0 0.00023998 3.3 0.0002399 3.3 0.00024 0 0.00023992 0 0.00024002 3.3 0.00023993999999999998 3.3 0.00024003999999999999 0 0.00023996 0 0.00024006 3.3 0.00023998 3.3 0.00024008 0 0.00024 0 0.0002401 3.3 0.00024002 3.3 0.00024012 0 0.00024003999999999999 0 0.00024014 3.3 0.00024006 3.3 0.00024016 0 0.00024008 0 0.00024018 3.3 0.00024009999999999998 3.3 0.00024019999999999998 0 0.00024012 0 0.00024022 3.3 0.00024014 3.3 0.00024024 0 0.00024016 0 0.00024026 3.3 0.00024018 3.3 0.00024028 0 0.00024019999999999998 0 0.00024029999999999999 3.3 0.00024022 3.3 0.00024032 0 0.00024024 0 0.00024034 3.3 0.00024025999999999998 3.3 0.00024035999999999998 0 0.00024028 0 0.00024038 3.3 0.00024029999999999999 3.3 0.0002404 0 0.00024032 0 0.00024042 3.3 0.00024034 3.3 0.00024044 0 0.00024035999999999998 0 0.00024045999999999998 3.3 0.00024038 3.3 0.00024048 0 0.0002404 0 0.0002405 3.3 0.00024042 3.3 0.00024052 0 0.00024044 0 0.00024054 3.3 0.00024045999999999998 3.3 0.00024056 0 0.00024048 0 0.00024058 3.3 0.0002405 3.3 0.0002406 0 0.00024051999999999998 0 0.00024061999999999998 3.3 0.00024054 3.3 0.00024064 0 0.00024056 0 0.00024066 3.3 0.00024058 3.3 0.00024068 0 0.0002406 0 0.0002407 3.3 0.00024061999999999998 3.3 0.00024071999999999999 0 0.00024064 0 0.00024074 3.3 0.00024066 3.3 0.00024076 0 0.00024067999999999998 0 0.00024077999999999998 3.3 0.0002407 3.3 0.0002408 0 0.00024071999999999999 0 0.00024082 3.3 0.00024074 3.3 0.00024084 0 0.00024076 0 0.00024086 3.3 0.00024077999999999998 3.3 0.00024087999999999998 0 0.0002408 0 0.0002409 3.3 0.00024082 3.3 0.00024092 0 0.00024084 0 0.00024094 3.3 0.00024086 3.3 0.00024096 0 0.00024087999999999998 0 0.00024098 3.3 0.0002409 3.3 0.000241 0 0.00024092 0 0.00024102 3.3 0.00024093999999999998 3.3 0.00024103999999999998 0 0.00024096 0 0.00024106 3.3 0.00024098 3.3 0.00024108 0 0.000241 0 0.0002411 3.3 0.00024102 3.3 0.00024112 0 0.00024103999999999998 0 0.00024113999999999999 3.3 0.00024106 3.3 0.00024116 0 0.00024108 0 0.00024118 3.3 0.0002411 3.3 0.0002412 0 0.00024112 0 0.00024122 3.3 0.00024113999999999999 3.3 0.00024124 0 0.00024116 0 0.00024126 3.3 0.00024118 3.3 0.00024128 0 0.00024119999999999998 0 0.00024129999999999998 3.3 0.00024122 3.3 0.00024132 0 0.00024124 0 0.00024134 3.3 0.00024126 3.3 0.00024136 0 0.00024128 0 0.00024138 3.3 0.00024129999999999998 3.3 0.00024139999999999999 0 0.00024132 0 0.00024142 3.3 0.00024134 3.3 0.00024144 0 0.00024135999999999998 0 0.00024145999999999998 3.3 0.00024138 3.3 0.00024148 0 0.00024139999999999999 0 0.0002415 3.3 0.00024142 3.3 0.00024152 0 0.00024144 0 0.00024154 3.3 0.00024145999999999998 3.3 0.00024155999999999998 0 0.00024148 0 0.00024158 3.3 0.0002415 3.3 0.0002416 0 0.00024152 0 0.00024162 3.3 0.00024154 3.3 0.00024164 0 0.00024155999999999998 0 0.00024166 3.3 0.00024158 3.3 0.00024168 0 0.0002416 0 0.0002417 3.3 0.00024161999999999998 3.3 0.00024171999999999998 0 0.00024164 0 0.00024174 3.3 0.00024166 3.3 0.00024176 0 0.00024168 0 0.00024178 3.3 0.0002417 3.3 0.0002418 0 0.00024171999999999998 0 0.00024181999999999999 3.3 0.00024174 3.3 0.00024184 0 0.00024176 0 0.00024186 3.3 0.00024178 3.3 0.00024188 0 0.0002418 0 0.0002419 3.3 0.00024181999999999999 3.3 0.00024192 0 0.00024184 0 0.00024194 3.3 0.00024186 3.3 0.00024196 0 0.00024187999999999998 0 0.00024197999999999998 3.3 0.0002419 3.3 0.000242 0 0.00024192 0 0.00024202 3.3 0.00024194 3.3 0.00024204 0 0.00024196 0 0.00024206 3.3 0.00024197999999999998 3.3 0.00024207999999999999 0 0.000242 0 0.0002421 3.3 0.00024202 3.3 0.00024212 0 0.00024203999999999998 0 0.00024213999999999998 3.3 0.00024206 3.3 0.00024216 0 0.00024207999999999999 0 0.00024218 3.3 0.0002421 3.3 0.0002422 0 0.00024212 0 0.00024222 3.3 0.00024213999999999998 3.3 0.00024223999999999998 0 0.00024216 0 0.00024226 3.3 0.00024218 3.3 0.00024228 0 0.0002422 0 0.0002423 3.3 0.00024222 3.3 0.00024232 0 0.00024223999999999998 0 0.00024234 3.3 0.00024226 3.3 0.00024236 0 0.00024228 0 0.00024238 3.3 0.00024229999999999998 3.3 0.00024239999999999998 0 0.00024232 0 0.00024242 3.3 0.00024234 3.3 0.00024244 0 0.00024236 0 0.00024246 3.3 0.00024238 3.3 0.00024248 0 0.00024239999999999998 0 0.00024249999999999999 3.3 0.00024242 3.3 0.00024252 0 0.00024244 0 0.00024254 3.3 0.00024245999999999998 3.3 0.00024255999999999998 0 0.00024248 0 0.00024258 3.3 0.00024249999999999999 3.3 0.0002426 0 0.00024252 0 0.00024262 3.3 0.00024254 3.3 0.00024264 0 0.00024255999999999998 0 0.00024265999999999998 3.3 0.00024258 3.3 0.00024268 0 0.0002426 0 0.0002427 3.3 0.00024262 3.3 0.00024272 0 0.00024264 0 0.00024274 3.3 0.00024265999999999998 3.3 0.00024275999999999999 0 0.00024268 0 0.00024278 3.3 0.0002427 3.3 0.0002428 0 0.00024271999999999998 0 0.00024281999999999998 3.3 0.00024274 3.3 0.00024284 0 0.00024275999999999999 0 0.00024286 3.3 0.00024278 3.3 0.00024288 0 0.0002428 0 0.0002429 3.3 0.00024281999999999998 3.3 0.00024291999999999998 0 0.00024284 0 0.00024294 3.3 0.00024286 3.3 0.00024296 0 0.00024288 0 0.00024298 3.3 0.0002429 3.3 0.000243 0 0.00024291999999999998 0 0.00024302 3.3 0.00024294 3.3 0.00024304 0 0.00024296 0 0.00024306 3.3 0.00024297999999999998 3.3 0.00024307999999999998 0 0.000243 0 0.0002431 3.3 0.00024302 3.3 0.00024312 0 0.00024304 0 0.00024314 3.3 0.00024306 3.3 0.00024316 0 0.00024307999999999998 0 0.00024317999999999999 3.3 0.0002431 3.3 0.0002432 0 0.00024312 0 0.00024322 3.3 0.00024313999999999998 3.3 0.00024323999999999998 0 0.00024316 0 0.00024326 3.3 0.00024317999999999999 3.3 0.00024328 0 0.0002432 0 0.0002433 3.3 0.00024322 3.3 0.00024332 0 0.00024323999999999998 0 0.00024333999999999998 3.3 0.00024326 3.3 0.00024336 0 0.00024328 0 0.00024338 3.3 0.0002433 3.3 0.0002434 0 0.00024332 0 0.00024342 3.3 0.00024333999999999998 3.3 0.00024344 0 0.00024336 0 0.00024346 3.3 0.00024338 3.3 0.00024348 0 0.00024339999999999998 0 0.00024349999999999998 3.3 0.00024342 3.3 0.00024352 0 0.00024344 0 0.00024354 3.3 0.00024346 3.3 0.00024356 0 0.00024348 0 0.00024358 3.3 0.00024349999999999998 3.3 0.00024359999999999999 0 0.00024352 0 0.00024362 3.3 0.00024354 3.3 0.00024364 0 0.00024356 0 0.00024366 3.3 0.00024358 3.3 0.00024368 0 0.00024359999999999999 0 0.0002437 3.3 0.00024362 3.3 0.00024372 0 0.00024364 0 0.00024374 3.3 0.00024365999999999998 3.3 0.00024375999999999998 0 0.00024368 0 0.00024378 3.3 0.0002437 3.3 0.0002438 0 0.00024372 0 0.00024382 3.3 0.00024374 3.3 0.00024384 0 0.00024375999999999998 0 0.00024385999999999999 3.3 0.00024378 3.3 0.00024388 0 0.0002438 0 0.0002439 3.3 0.00024381999999999998 3.3 0.00024391999999999998 0 0.00024384 0 0.00024394 3.3 0.00024385999999999999 3.3 0.00024396 0 0.00024388 0 0.00024398 3.3 0.0002439 3.3 0.000244 0 0.00024391999999999998 0 0.00024401999999999998 3.3 0.00024394 3.3 0.00024404 0 0.00024396 0 0.00024406 3.3 0.00024398 3.3 0.00024408 0 0.000244 0 0.0002441 3.3 0.00024401999999999998 3.3 0.00024412 0 0.00024404 0 0.00024414 3.3 0.00024406 3.3 0.00024416 0 0.00024407999999999998 0 0.00024418 3.3 0.00024409999999999997 3.3 0.00024419999999999997 0 0.00024412000000000001 0 0.00024422 3.3 0.00024414 3.3 0.00024424 0 0.00024416 0 0.00024426 3.3 0.00024418 3.3 0.00024428 0 0.00024419999999999997 0 0.0002443 3.3 0.00024422 3.3 0.00024432 0 0.00024424 0 0.00024434 3.3 0.00024426 3.3 0.00024436 0 0.00024428 0 0.00024438 3.3 0.0002443 3.3 0.0002444 0 0.00024432 0 0.00024442 3.3 0.00024434 3.3 0.00024444 0 0.00024436 0 0.00024446 3.3 0.00024438 3.3 0.00024448 0 0.0002444 0 0.0002445 3.3 0.00024441999999999997 3.3 0.00024451999999999997 0 0.00024444 0 0.00024454 3.3 0.00024446 3.3 0.00024456 0 0.00024448 0 0.00024458 3.3 0.0002445 3.3 0.0002446 0 0.00024451999999999997 0 0.00024461999999999997 3.3 0.00024454 3.3 0.00024464 0 0.00024456 0 0.00024466 3.3 0.00024458 3.3 0.00024468 0 0.0002446 0 0.0002447 3.3 0.00024461999999999997 3.3 0.00024472 0 0.00024464 0 0.00024474 3.3 0.00024466 3.3 0.00024476 0 0.00024468 0 0.00024478 3.3 0.0002447 3.3 0.0002448 0 0.00024472 0 0.00024482 3.3 0.00024474 3.3 0.00024484 0 0.00024476 0 0.00024486 3.3 0.00024478 3.3 0.00024488 0 0.0002448 0 0.0002449 3.3 0.00024482 3.3 0.00024492 0 0.00024483999999999997 0 0.00024493999999999997 3.3 0.00024486 3.3 0.00024496 0 0.00024488 0 0.00024498 3.3 0.0002449 3.3 0.000245 0 0.00024492 0 0.00024502 3.3 0.00024493999999999997 3.3 0.00024503999999999997 0 0.00024496 0 0.00024506 3.3 0.00024498 3.3 0.00024508 0 0.000245 0 0.0002451 3.3 0.00024502 3.3 0.00024512 0 0.00024503999999999997 0 0.00024514 3.3 0.00024506 3.3 0.00024516 0 0.00024508 0 0.00024518 3.3 0.0002451 3.3 0.0002452 0 0.00024512 0 0.00024522 3.3 0.00024514 3.3 0.00024524 0 0.00024516 0 0.00024526 3.3 0.00024518 3.3 0.00024528 0 0.0002452 0 0.0002453 3.3 0.00024522 3.3 0.00024532 0 0.00024524 0 0.00024534 3.3 0.00024525999999999997 3.3 0.00024535999999999997 0 0.00024528 0 0.00024538 3.3 0.0002453 3.3 0.0002454 0 0.00024532 0 0.00024542 3.3 0.00024534 3.3 0.00024544 0 0.00024535999999999997 0 0.00024545999999999997 3.3 0.00024538 3.3 0.00024548 0 0.0002454 0 0.0002455 3.3 0.00024542 3.3 0.00024552 0 0.00024544 0 0.00024554 3.3 0.00024545999999999997 3.3 0.00024556 0 0.00024548 0 0.00024558 3.3 0.0002455 3.3 0.0002456 0 0.00024552 0 0.00024562 3.3 0.00024554 3.3 0.00024564 0 0.00024556 0 0.00024566 3.3 0.00024558 3.3 0.00024568 0 0.0002456 0 0.0002457 3.3 0.00024562 3.3 0.00024572 0 0.00024564 0 0.00024574 3.3 0.00024566 3.3 0.00024576 0 0.00024568 0 0.00024578 3.3 0.0002457 3.3 0.0002458 0 0.00024572 0 0.00024582 3.3 0.00024574 3.3 0.00024584 0 0.00024576 0 0.00024586 3.3 0.00024577999999999997 3.3 0.00024587999999999997 0 0.0002458 0 0.0002459 3.3 0.00024582 3.3 0.00024592 0 0.00024584 0 0.00024594 3.3 0.00024586 3.3 0.00024596 0 0.00024587999999999997 0 0.00024597999999999997 3.3 0.0002459 3.3 0.000246 0 0.00024592 0 0.00024602 3.3 0.00024594 3.3 0.00024604 0 0.00024596 0 0.00024606 3.3 0.00024597999999999997 3.3 0.00024608 0 0.000246 0 0.0002461 3.3 0.00024602 3.3 0.00024612 0 0.00024604 0 0.00024614 3.3 0.00024606 3.3 0.00024616 0 0.00024608 0 0.00024618 3.3 0.0002461 3.3 0.0002462 0 0.00024612 0 0.00024622 3.3 0.00024614 3.3 0.00024624 0 0.00024616 0 0.00024626 3.3 0.00024618 3.3 0.00024628 0 0.00024619999999999997 0 0.00024629999999999997 3.3 0.00024622 3.3 0.00024632 0 0.00024624 0 0.00024634 3.3 0.00024626 3.3 0.00024636 0 0.00024628 0 0.00024638 3.3 0.00024629999999999997 3.3 0.00024639999999999997 0 0.00024632 0 0.00024642 3.3 0.00024634 3.3 0.00024644 0 0.00024636 0 0.00024646 3.3 0.00024638 3.3 0.00024648 0 0.00024639999999999997 0 0.0002465 3.3 0.00024642 3.3 0.00024652 0 0.00024644 0 0.00024654 3.3 0.00024646 3.3 0.00024656 0 0.00024648 0 0.00024658 3.3 0.0002465 3.3 0.0002466 0 0.00024652 0 0.00024662 3.3 0.00024654 3.3 0.00024664 0 0.00024656 0 0.00024666 3.3 0.00024658 3.3 0.00024668 0 0.0002466 0 0.0002467 3.3 0.00024661999999999997 3.3 0.00024671999999999997 0 0.00024664 0 0.00024674 3.3 0.00024666 3.3 0.00024676 0 0.00024668 0 0.00024678 3.3 0.0002467 3.3 0.0002468 0 0.00024671999999999997 0 0.00024681999999999997 3.3 0.00024674 3.3 0.00024684 0 0.00024676 0 0.00024686 3.3 0.00024678 3.3 0.00024688 0 0.0002468 0 0.0002469 3.3 0.00024681999999999997 3.3 0.00024692 0 0.00024684 0 0.00024694 3.3 0.00024686 3.3 0.00024696 0 0.00024688 0 0.00024698 3.3 0.0002469 3.3 0.000247 0 0.00024692 0 0.00024702 3.3 0.00024694 3.3 0.00024704 0 0.00024696 0 0.00024706 3.3 0.00024698 3.3 0.00024708 0 0.000247 0 0.0002471 3.3 0.00024702 3.3 0.00024712 0 0.00024703999999999997 0 0.00024713999999999997 3.3 0.00024706 3.3 0.00024716 0 0.00024708 0 0.00024718 3.3 0.0002471 3.3 0.0002472 0 0.00024712 0 0.00024722 3.3 0.00024713999999999997 3.3 0.00024723999999999997 0 0.00024716 0 0.00024726 3.3 0.00024718 3.3 0.00024728 0 0.0002472 0 0.0002473 3.3 0.00024722 3.3 0.00024732 0 0.00024723999999999997 0 0.00024734 3.3 0.00024726 3.3 0.00024736 0 0.00024728 0 0.00024738 3.3 0.0002473 3.3 0.0002474 0 0.00024732 0 0.00024742 3.3 0.00024734 3.3 0.00024744 0 0.00024736 0 0.00024746 3.3 0.00024738 3.3 0.00024748 0 0.0002474 0 0.0002475 3.3 0.00024742 3.3 0.00024752 0 0.00024744 0 0.00024754 3.3 0.00024746 3.3 0.00024756 0 0.00024748 0 0.00024758 3.3 0.0002475 3.3 0.0002476 0 0.00024752 0 0.00024762 3.3 0.00024754 3.3 0.00024764 0 0.00024755999999999997 0 0.00024765999999999997 3.3 0.00024758 3.3 0.00024768 0 0.0002476 0 0.0002477 3.3 0.00024762 3.3 0.00024772 0 0.00024764 0 0.00024774 3.3 0.00024765999999999997 3.3 0.00024775999999999997 0 0.00024768 0 0.00024778 3.3 0.0002477 3.3 0.0002478 0 0.00024772 0 0.00024782 3.3 0.00024774 3.3 0.00024784 0 0.00024775999999999997 0 0.00024786 3.3 0.00024778 3.3 0.00024788 0 0.0002478 0 0.0002479 3.3 0.00024782 3.3 0.00024792 0 0.00024784 0 0.00024794 3.3 0.00024786 3.3 0.00024796 0 0.00024788 0 0.00024798 3.3 0.0002479 3.3 0.000248 0 0.00024792 0 0.00024802 3.3 0.00024794 3.3 0.00024804 0 0.00024796 0 0.00024806 3.3 0.00024797999999999997 3.3 0.00024807999999999997 0 0.000248 0 0.0002481 3.3 0.00024802 3.3 0.00024812 0 0.00024804 0 0.00024814 3.3 0.00024806 3.3 0.00024816 0 0.00024807999999999997 0 0.00024817999999999997 3.3 0.0002481 3.3 0.0002482 0 0.00024812 0 0.00024822 3.3 0.00024814 3.3 0.00024824 0 0.00024816 0 0.00024826 3.3 0.00024817999999999997 3.3 0.00024828 0 0.0002482 0 0.0002483 3.3 0.00024822 3.3 0.00024832 0 0.00024824 0 0.00024834 3.3 0.00024826 3.3 0.00024836 0 0.00024828 0 0.00024838 3.3 0.0002483 3.3 0.0002484 0 0.00024832 0 0.00024842 3.3 0.00024834 3.3 0.00024844 0 0.00024836 0 0.00024846 3.3 0.00024838 3.3 0.00024848 0 0.00024839999999999997 0 0.00024849999999999997 3.3 0.00024842 3.3 0.00024852 0 0.00024844 0 0.00024854 3.3 0.00024846 3.3 0.00024856 0 0.00024848 0 0.00024858 3.3 0.00024849999999999997 3.3 0.00024859999999999997 0 0.00024852 0 0.00024862 3.3 0.00024854 3.3 0.00024864 0 0.00024856 0 0.00024866 3.3 0.00024858 3.3 0.00024868 0 0.00024859999999999997 0 0.0002487 3.3 0.00024862 3.3 0.00024872 0 0.00024864 0 0.00024874 3.3 0.00024866 3.3 0.00024876 0 0.00024868 0 0.00024878 3.3 0.0002487 3.3 0.0002488 0 0.00024872 0 0.00024882 3.3 0.00024874 3.3 0.00024884 0 0.00024876 0 0.00024886 3.3 0.00024878 3.3 0.00024888 0 0.0002488 0 0.0002489 3.3 0.00024881999999999997 3.3 0.00024891999999999997 0 0.00024884 0 0.00024894 3.3 0.00024886 3.3 0.00024896 0 0.00024888 0 0.00024898 3.3 0.0002489 3.3 0.000249 0 0.00024891999999999997 0 0.00024901999999999997 3.3 0.00024894 3.3 0.00024904 0 0.00024896 0 0.00024906 3.3 0.00024898 3.3 0.00024908 0 0.000249 0 0.0002491 3.3 0.00024901999999999997 3.3 0.00024912 0 0.00024904 0 0.00024914 3.3 0.00024906 3.3 0.00024916 0 0.00024908 0 0.00024918 3.3 0.0002491 3.3 0.0002492 0 0.00024912 0 0.00024922 3.3 0.00024914 3.3 0.00024924 0 0.00024916 0 0.00024926 3.3 0.00024918 3.3 0.00024928 0 0.0002492 0 0.0002493 3.3 0.00024922 3.3 0.00024932 0 0.00024924 0 0.00024934 3.3 0.00024926 3.3 0.00024936 0 0.00024928 0 0.00024938 3.3 0.0002493 3.3 0.0002494 0 0.00024932 0 0.00024942 3.3 0.00024933999999999997 3.3 0.00024943999999999997 0 0.00024936 0 0.00024946 3.3 0.00024938 3.3 0.00024948 0 0.0002494 0 0.0002495 3.3 0.00024942 3.3 0.00024952 0 0.00024943999999999997 0 0.00024953999999999997 3.3 0.00024946 3.3 0.00024956 0 0.00024948 0 0.00024958 3.3 0.0002495 3.3 0.0002496 0 0.00024952 0 0.00024962 3.3 0.00024953999999999997 3.3 0.00024964 0 0.00024956 0 0.00024966 3.3 0.00024958 3.3 0.00024968 0 0.0002496 0 0.0002497 3.3 0.00024962 3.3 0.00024972 0 0.00024964 0 0.00024974 3.3 0.00024966 3.3 0.00024976 0 0.00024968 0 0.00024978 3.3 0.0002497 3.3 0.0002498 0 0.00024972 0 0.00024982 3.3 0.00024974 3.3 0.00024984 0 0.00024975999999999997 0 0.00024985999999999997 3.3 0.00024978 3.3 0.00024988 0 0.0002498 0 0.0002499 3.3 0.00024982 3.3 0.00024992 0 0.00024984 0 0.00024994 3.3 0.00024985999999999997 3.3 0.00024995999999999997 0 0.00024988 0 0.00024998 3.3 0.0002499 3.3 0.00025 0 0.00024992 0 0.00025002 3.3 0.00024994 3.3 0.00025004 0 0.00024995999999999997 0 0.00025006 3.3 0.00024998 3.3 0.00025008 0 0.00025 0 0.0002501 3.3 0.00025002 3.3 0.00025012 0 0.00025004 0 0.00025014 3.3 0.00025006 3.3 0.00025016 0 0.00025008 0 0.00025018 3.3 0.0002501 3.3 0.0002502 0 0.00025012 0 0.00025022 3.3 0.00025014 3.3 0.00025024 0 0.00025016 0 0.00025026 3.3 0.00025017999999999997 3.3 0.00025027999999999997 0 0.0002502 0 0.0002503 3.3 0.00025022 3.3 0.00025032 0 0.00025024 0 0.00025034 3.3 0.00025026 3.3 0.00025036 0 0.00025027999999999997 0 0.00025037999999999997 3.3 0.0002503 3.3 0.0002504 0 0.00025032 0 0.00025042 3.3 0.00025034 3.3 0.00025044 0 0.00025036 0 0.00025046 3.3 0.00025037999999999997 3.3 0.00025048 0 0.0002504 0 0.0002505 3.3 0.00025042 3.3 0.00025052 0 0.00025044 0 0.00025054 3.3 0.00025046 3.3 0.00025056 0 0.00025048 0 0.00025058 3.3 0.0002505 3.3 0.0002506 0 0.00025052 0 0.00025062 3.3 0.00025054 3.3 0.00025064 0 0.00025056 0 0.00025066 3.3 0.00025058 3.3 0.00025068 0 0.00025059999999999997 0 0.00025069999999999997 3.3 0.00025062 3.3 0.00025072 0 0.00025064 0 0.00025074 3.3 0.00025066 3.3 0.00025076 0 0.00025068 0 0.00025078 3.3 0.00025069999999999997 3.3 0.00025079999999999997 0 0.00025072 0 0.00025082 3.3 0.00025074 3.3 0.00025084 0 0.00025076 0 0.00025086 3.3 0.00025078 3.3 0.00025088 0 0.00025079999999999997 0 0.00025089999999999997 3.3 0.00025082 3.3 0.00025092 0 0.00025084 0 0.00025094 3.3 0.00025086 3.3 0.00025096 0 0.00025088 0 0.00025098 3.3 0.00025089999999999997 3.3 0.000251 0 0.00025092 0 0.00025102 3.3 0.00025094 3.3 0.00025104 0 0.00025096 0 0.00025106 3.3 0.00025098 3.3 0.00025108 0 0.000251 0 0.0002511 3.3 0.00025102 3.3 0.00025112 0 0.00025104 0 0.00025114 3.3 0.00025106 3.3 0.00025116 0 0.00025108 0 0.00025118 3.3 0.0002511 3.3 0.0002512 0 0.00025111999999999997 0 0.00025121999999999997 3.3 0.00025114 3.3 0.00025124 0 0.00025116 0 0.00025126 3.3 0.00025118 3.3 0.00025128 0 0.0002512 0 0.0002513 3.3 0.00025121999999999997 3.3 0.00025131999999999997 0 0.00025124 0 0.00025134 3.3 0.00025126 3.3 0.00025136 0 0.00025128 0 0.00025138 3.3 0.0002513 3.3 0.0002514 0 0.00025131999999999997 0 0.00025142 3.3 0.00025134 3.3 0.00025144 0 0.00025136 0 0.00025146 3.3 0.00025138 3.3 0.00025148 0 0.0002514 0 0.0002515 3.3 0.00025142 3.3 0.00025152 0 0.00025144 0 0.00025154 3.3 0.00025146 3.3 0.00025156 0 0.00025148 0 0.00025158 3.3 0.0002515 3.3 0.0002516 0 0.00025152 0 0.00025162 3.3 0.00025153999999999997 3.3 0.00025163999999999997 0 0.00025156 0 0.00025166 3.3 0.00025158 3.3 0.00025168 0 0.0002516 0 0.0002517 3.3 0.00025162 3.3 0.00025172 0 0.00025163999999999997 0 0.00025173999999999997 3.3 0.00025166 3.3 0.00025176 0 0.00025168 0 0.00025178 3.3 0.0002517 3.3 0.0002518 0 0.00025172 0 0.00025182 3.3 0.00025173999999999997 3.3 0.00025184 0 0.00025176 0 0.00025186 3.3 0.00025178 3.3 0.00025188 0 0.0002518 0 0.0002519 3.3 0.00025182 3.3 0.00025192 0 0.00025184 0 0.00025194 3.3 0.00025186 3.3 0.00025196 0 0.00025188 0 0.00025198 3.3 0.0002519 3.3 0.000252 0 0.00025192 0 0.00025202 3.3 0.00025194 3.3 0.00025204 0 0.00025195999999999997 0 0.00025205999999999997 3.3 0.00025198 3.3 0.00025208 0 0.000252 0 0.0002521 3.3 0.00025202 3.3 0.00025212 0 0.00025204 0 0.00025214 3.3 0.00025205999999999997 3.3 0.00025215999999999997 0 0.00025208 0 0.00025218 3.3 0.0002521 3.3 0.0002522 0 0.00025212 0 0.00025222 3.3 0.00025214 3.3 0.00025224 0 0.00025215999999999997 0 0.00025226 3.3 0.00025218 3.3 0.00025228 0 0.0002522 0 0.0002523 3.3 0.00025222 3.3 0.00025232 0 0.00025224 0 0.00025234 3.3 0.00025226 3.3 0.00025236 0 0.00025228 0 0.00025238 3.3 0.0002523 3.3 0.0002524 0 0.00025232 0 0.00025242 3.3 0.00025234 3.3 0.00025244 0 0.00025236 0 0.00025246 3.3 0.00025237999999999997 3.3 0.00025247999999999997 0 0.0002524 0 0.0002525 3.3 0.00025242 3.3 0.00025252 0 0.00025244 0 0.00025254 3.3 0.00025246 3.3 0.00025256 0 0.00025247999999999997 0 0.00025257999999999997 3.3 0.0002525 3.3 0.0002526 0 0.00025252 0 0.00025262 3.3 0.00025254 3.3 0.00025264 0 0.00025256 0 0.00025266 3.3 0.00025257999999999997 3.3 0.00025267999999999997 0 0.0002526 0 0.0002527 3.3 0.00025262 3.3 0.00025272 0 0.00025264 0 0.00025274 3.3 0.00025266 3.3 0.00025276 0 0.00025267999999999997 0 0.00025278 3.3 0.0002527 3.3 0.0002528 0 0.00025272 0 0.00025282 3.3 0.00025274 3.3 0.00025284 0 0.00025276 0 0.00025286 3.3 0.00025278 3.3 0.00025288 0 0.0002528 0 0.0002529 3.3 0.00025282 3.3 0.00025292 0 0.00025284 0 0.00025294 3.3 0.00025286 3.3 0.00025296 0 0.00025288 0 0.00025298 3.3 0.00025289999999999997 3.3 0.00025299999999999997 0 0.00025292 0 0.00025302 3.3 0.00025294 3.3 0.00025304 0 0.00025296 0 0.00025306 3.3 0.00025298 3.3 0.00025308 0 0.00025299999999999997 0 0.00025309999999999997 3.3 0.00025302 3.3 0.00025312 0 0.00025304 0 0.00025314 3.3 0.00025306 3.3 0.00025316 0 0.00025308 0 0.00025318 3.3 0.00025309999999999997 3.3 0.0002532 0 0.00025312 0 0.00025322 3.3 0.00025314 3.3 0.00025324 0 0.00025316 0 0.00025326 3.3 0.00025318 3.3 0.00025328 0 0.0002532 0 0.0002533 3.3 0.00025322 3.3 0.00025332 0 0.00025324 0 0.00025334 3.3 0.00025326 3.3 0.00025336 0 0.00025328 0 0.00025338 3.3 0.0002533 3.3 0.0002534 0 0.00025331999999999997 0 0.00025341999999999997 3.3 0.00025334 3.3 0.00025344 0 0.00025336 0 0.00025346 3.3 0.00025338 3.3 0.00025348 0 0.0002534 0 0.0002535 3.3 0.00025341999999999997 3.3 0.00025351999999999997 0 0.00025344 0 0.00025354 3.3 0.00025346 3.3 0.00025356 0 0.00025348 0 0.00025358 3.3 0.0002535 3.3 0.0002536 0 0.00025351999999999997 0 0.00025362 3.3 0.00025354 3.3 0.00025364 0 0.00025356 0 0.00025366 3.3 0.00025358 3.3 0.00025368 0 0.0002536 0 0.0002537 3.3 0.00025362 3.3 0.00025372 0 0.00025364 0 0.00025374 3.3 0.00025366 3.3 0.00025376 0 0.00025368 0 0.00025378 3.3 0.0002537 3.3 0.0002538 0 0.00025372 0 0.00025382 3.3 0.00025373999999999997 3.3 0.00025383999999999997 0 0.00025376 0 0.00025386 3.3 0.00025378 3.3 0.00025388 0 0.0002538 0 0.0002539 3.3 0.00025382 3.3 0.00025392 0 0.00025383999999999997 0 0.00025393999999999997 3.3 0.00025386 3.3 0.00025396 0 0.00025388 0 0.00025398 3.3 0.0002539 3.3 0.000254 0 0.00025392 0 0.00025402 3.3 0.00025393999999999997 3.3 0.00025404 0 0.00025396 0 0.00025406 3.3 0.00025398 3.3 0.00025408 0 0.000254 0 0.0002541 3.3 0.00025402 3.3 0.00025412 0 0.00025404 0 0.00025414 3.3 0.00025406 3.3 0.00025416 0 0.00025408 0 0.00025418 3.3 0.0002541 3.3 0.0002542 0 0.00025412 0 0.00025422 3.3 0.00025414 3.3 0.00025424 0 0.00025415999999999997 0 0.00025425999999999997 3.3 0.00025418 3.3 0.00025428 0 0.0002542 0 0.0002543 3.3 0.00025422 3.3 0.00025432 0 0.00025424 0 0.00025434 3.3 0.00025425999999999997 3.3 0.00025435999999999997 0 0.00025428 0 0.00025438 3.3 0.0002543 3.3 0.0002544 0 0.00025432 0 0.00025442 3.3 0.00025434 3.3 0.00025444 0 0.00025435999999999997 0 0.00025445999999999997 3.3 0.00025438 3.3 0.00025448 0 0.0002544 0 0.0002545 3.3 0.00025442 3.3 0.00025452 0 0.00025444 0 0.00025454 3.3 0.00025445999999999997 3.3 0.00025456 0 0.00025448 0 0.00025458 3.3 0.0002545 3.3 0.0002546 0 0.00025452 0 0.00025462 3.3 0.00025454 3.3 0.00025464 0 0.00025456 0 0.00025466 3.3 0.00025458 3.3 0.00025468 0 0.0002546 0 0.0002547 3.3 0.00025462 3.3 0.00025472 0 0.00025464 0 0.00025474 3.3 0.00025466 3.3 0.00025476 0 0.00025467999999999997 0 0.00025477999999999997 3.3 0.0002547 3.3 0.0002548 0 0.00025472 0 0.00025482 3.3 0.00025474 3.3 0.00025484 0 0.00025476 0 0.00025486 3.3 0.00025477999999999997 3.3 0.00025487999999999997 0 0.0002548 0 0.0002549 3.3 0.00025482 3.3 0.00025492 0 0.00025484 0 0.00025494 3.3 0.00025486 3.3 0.00025496 0 0.00025487999999999997 0 0.00025498 3.3 0.0002549 3.3 0.000255 0 0.00025492 0 0.00025502 3.3 0.00025494 3.3 0.00025504 0 0.00025496 0 0.00025506 3.3 0.00025498 3.3 0.00025508 0 0.000255 0 0.0002551 3.3 0.00025502 3.3 0.00025512 0 0.00025504 0 0.00025514 3.3 0.00025506 3.3 0.00025516 0 0.00025508 0 0.00025518 3.3 0.00025509999999999997 3.3 0.00025519999999999997 0 0.00025512 0 0.00025522 3.3 0.00025514 3.3 0.00025524 0 0.00025516 0 0.00025526 3.3 0.00025518 3.3 0.00025528 0 0.00025519999999999997 0 0.00025529999999999997 3.3 0.00025522 3.3 0.00025532 0 0.00025524 0 0.00025534 3.3 0.00025526 3.3 0.00025536 0 0.00025528 0 0.00025538 3.3 0.00025529999999999997 3.3 0.0002554 0 0.00025532 0 0.00025542 3.3 0.00025534 3.3 0.00025544 0 0.00025536 0 0.00025546 3.3 0.00025538 3.3 0.00025548 0 0.0002554 0 0.0002555 3.3 0.00025542 3.3 0.00025552 0 0.00025544 0 0.00025554 3.3 0.00025546 3.3 0.00025556 0 0.00025548 0 0.00025558 3.3 0.0002555 3.3 0.0002556 0 0.00025551999999999997 0 0.00025561999999999997 3.3 0.00025554 3.3 0.00025564 0 0.00025556 0 0.00025566 3.3 0.00025558 3.3 0.00025568 0 0.0002556 0 0.0002557 3.3 0.00025561999999999997 3.3 0.00025571999999999997 0 0.00025564 0 0.00025574 3.3 0.00025566 3.3 0.00025576 0 0.00025568 0 0.00025578 3.3 0.0002557 3.3 0.0002558 0 0.00025571999999999997 0 0.00025582 3.3 0.00025574 3.3 0.00025584 0 0.00025576 0 0.00025586 3.3 0.00025578 3.3 0.00025588 0 0.0002558 0 0.0002559 3.3 0.00025582 3.3 0.00025592 0 0.00025584 0 0.00025594 3.3 0.00025586 3.3 0.00025596 0 0.00025588 0 0.00025598 3.3 0.0002559 3.3 0.000256 0 0.00025592 0 0.00025602 3.3 0.00025594 3.3 0.00025604 0 0.00025596 0 0.00025606 3.3 0.00025598 3.3 0.00025608 0 0.000256 0 0.0002561 3.3 0.00025602 3.3 0.00025612 0 0.00025603999999999997 0 0.00025613999999999997 3.3 0.00025606 3.3 0.00025616 0 0.00025608 0 0.00025618 3.3 0.0002561 3.3 0.0002562 0 0.00025612 0 0.00025622 3.3 0.00025613999999999997 3.3 0.00025623999999999997 0 0.00025616 0 0.00025626 3.3 0.00025618 3.3 0.00025628 0 0.0002562 0 0.0002563 3.3 0.00025622 3.3 0.00025632 0 0.00025623999999999997 0 0.00025634 3.3 0.00025626 3.3 0.00025636 0 0.00025628 0 0.00025638 3.3 0.0002563 3.3 0.0002564 0 0.00025632 0 0.00025642 3.3 0.00025634 3.3 0.00025644 0 0.00025636 0 0.00025646 3.3 0.00025638 3.3 0.00025648 0 0.0002564 0 0.0002565 3.3 0.00025642 3.3 0.00025652 0 0.00025644 0 0.00025654 3.3 0.00025645999999999997 3.3 0.00025655999999999997 0 0.00025648 0 0.00025658 3.3 0.0002565 3.3 0.0002566 0 0.00025652 0 0.00025662 3.3 0.00025654 3.3 0.00025664 0 0.00025655999999999997 0 0.00025665999999999997 3.3 0.00025658 3.3 0.00025668 0 0.0002566 0 0.0002567 3.3 0.00025662 3.3 0.00025672 0 0.00025664 0 0.00025674 3.3 0.00025665999999999997 3.3 0.00025676 0 0.00025668 0 0.00025678 3.3 0.0002567 3.3 0.0002568 0 0.00025672 0 0.00025682 3.3 0.00025674 3.3 0.00025684 0 0.00025676 0 0.00025686 3.3 0.00025678 3.3 0.00025688 0 0.0002568 0 0.0002569 3.3 0.00025682 3.3 0.00025692 0 0.00025684 0 0.00025694 3.3 0.00025686 3.3 0.00025696 0 0.00025687999999999997 0 0.00025697999999999997 3.3 0.0002569 3.3 0.000257 0 0.00025692 0 0.00025702 3.3 0.00025694 3.3 0.00025704 0 0.00025696 0 0.00025706 3.3 0.00025697999999999997 3.3 0.00025707999999999997 0 0.000257 0 0.0002571 3.3 0.00025702 3.3 0.00025712 0 0.00025704 0 0.00025714 3.3 0.00025706 3.3 0.00025716 0 0.00025707999999999997 0 0.00025718 3.3 0.0002571 3.3 0.0002572 0 0.00025712 0 0.00025722 3.3 0.00025714 3.3 0.00025724 0 0.00025716 0 0.00025726 3.3 0.00025718 3.3 0.00025728 0 0.0002572 0 0.0002573 3.3 0.00025722 3.3 0.00025732 0 0.00025724 0 0.00025734 3.3 0.00025726 3.3 0.00025736 0 0.00025728 0 0.00025738 3.3 0.00025729999999999997 3.3 0.00025739999999999997 0 0.00025732 0 0.00025742 3.3 0.00025734 3.3 0.00025744 0 0.00025736 0 0.00025746 3.3 0.00025738 3.3 0.00025748 0 0.00025739999999999997 0 0.00025749999999999997 3.3 0.00025742 3.3 0.00025752 0 0.00025744 0 0.00025754 3.3 0.00025746 3.3 0.00025756 0 0.00025748 0 0.00025758 3.3 0.00025749999999999997 3.3 0.0002576 0 0.00025752 0 0.00025762 3.3 0.00025754 3.3 0.00025764 0 0.00025756 0 0.00025766 3.3 0.00025758 3.3 0.00025768 0 0.0002576 0 0.0002577 3.3 0.00025762 3.3 0.00025772 0 0.00025764 0 0.00025774 3.3 0.00025766 3.3 0.00025776 0 0.00025768 0 0.00025778 3.3 0.0002577 3.3 0.0002578 0 0.00025772 0 0.00025782 3.3 0.00025774 3.3 0.00025784 0 0.00025776 0 0.00025786 3.3 0.00025778 3.3 0.00025788 0 0.0002578 0 0.0002579 3.3 0.00025781999999999997 3.3 0.00025791999999999997 0 0.00025784 0 0.00025794 3.3 0.00025786 3.3 0.00025796 0 0.00025788 0 0.00025798 3.3 0.0002579 3.3 0.000258 0 0.00025791999999999997 0 0.00025801999999999997 3.3 0.00025794 3.3 0.00025804 0 0.00025796 0 0.00025806 3.3 0.00025798 3.3 0.00025808 0 0.000258 0 0.0002581 3.3 0.00025801999999999997 3.3 0.00025812 0 0.00025804 0 0.00025814 3.3 0.00025806 3.3 0.00025816 0 0.00025808 0 0.00025818 3.3 0.0002581 3.3 0.0002582 0 0.00025812 0 0.00025822 3.3 0.00025814 3.3 0.00025824 0 0.00025816 0 0.00025826 3.3 0.00025818 3.3 0.00025828 0 0.0002582 0 0.0002583 3.3 0.00025822 3.3 0.00025832 0 0.00025823999999999997 0 0.00025833999999999997 3.3 0.00025826 3.3 0.00025836 0 0.00025828 0 0.00025838 3.3 0.0002583 3.3 0.0002584 0 0.00025832 0 0.00025842 3.3 0.00025833999999999997 3.3 0.00025843999999999997 0 0.00025836 0 0.00025846 3.3 0.00025838 3.3 0.00025848 0 0.0002584 0 0.0002585 3.3 0.00025842 3.3 0.00025852 0 0.00025843999999999997 0 0.00025854 3.3 0.00025846 3.3 0.00025856 0 0.00025848 0 0.00025858 3.3 0.0002585 3.3 0.0002586 0 0.00025852 0 0.00025862 3.3 0.00025854 3.3 0.00025864 0 0.00025856 0 0.00025866 3.3 0.00025858 3.3 0.00025868 0 0.0002586 0 0.0002587 3.3 0.00025862 3.3 0.00025872 0 0.00025864 0 0.00025874 3.3 0.00025865999999999997 3.3 0.00025875999999999997 0 0.00025868 0 0.00025878 3.3 0.0002587 3.3 0.0002588 0 0.00025872 0 0.00025882 3.3 0.00025874 3.3 0.00025884 0 0.00025875999999999997 0 0.00025885999999999997 3.3 0.00025878 3.3 0.00025888 0 0.0002588 0 0.0002589 3.3 0.00025882 3.3 0.00025892 0 0.00025884 0 0.00025894 3.3 0.00025885999999999997 3.3 0.00025896 0 0.00025888 0 0.00025898 3.3 0.0002589 3.3 0.000259 0 0.00025892 0 0.00025902 3.3 0.00025894 3.3 0.00025904 0 0.00025896 0 0.00025906 3.3 0.00025898 3.3 0.00025908 0 0.000259 0 0.0002591 3.3 0.00025902 3.3 0.00025912 0 0.00025904 0 0.00025914 3.3 0.00025906 3.3 0.00025916 0 0.00025907999999999997 0 0.00025917999999999997 3.3 0.0002591 3.3 0.0002592 0 0.00025912 0 0.00025922 3.3 0.00025914 3.3 0.00025924 0 0.00025916 0 0.00025926 3.3 0.00025917999999999997 3.3 0.00025927999999999997 0 0.0002592 0 0.0002593 3.3 0.00025922 3.3 0.00025932 0 0.00025924 0 0.00025934 3.3 0.00025926 3.3 0.00025936 0 0.00025927999999999997 0 0.00025938 3.3 0.0002593 3.3 0.0002594 0 0.00025932 0 0.00025942 3.3 0.00025934 3.3 0.00025944 0 0.00025936 0 0.00025946 3.3 0.00025938 3.3 0.00025948 0 0.0002594 0 0.0002595 3.3 0.00025942 3.3 0.00025952 0 0.00025944 0 0.00025954 3.3 0.00025946 3.3 0.00025956 0 0.00025948 0 0.00025958 3.3 0.0002595 3.3 0.0002596 0 0.00025952 0 0.00025962 3.3 0.00025954 3.3 0.00025964 0 0.00025956 0 0.00025966 3.3 0.00025958 3.3 0.00025968 0 0.00025959999999999997 0 0.00025969999999999997 3.3 0.00025962 3.3 0.00025972 0 0.00025964 0 0.00025974 3.3 0.00025966 3.3 0.00025976 0 0.00025968 0 0.00025978 3.3 0.00025969999999999997 3.3 0.00025979999999999997 0 0.00025972 0 0.00025982 3.3 0.00025974 3.3 0.00025984 0 0.00025976 0 0.00025986 3.3 0.00025978 3.3 0.00025988 0 0.00025979999999999997 0 0.0002599 3.3 0.00025982 3.3 0.00025992 0 0.00025984 0 0.00025994 3.3 0.00025986 3.3 0.00025996 0 0.00025988 0 0.00025998 3.3 0.0002599 3.3 0.00026 0 0.00025992 0 0.00026002 3.3 0.00025994 3.3 0.00026004 0 0.00025996 0 0.00026006 3.3 0.00025998 3.3 0.00026008 0 0.00026 0 0.0002601 3.3 0.00026001999999999997 3.3 0.00026011999999999997 0 0.00026004 0 0.00026014 3.3 0.00026006 3.3 0.00026016 0 0.00026008 0 0.00026018 3.3 0.0002601 3.3 0.0002602 0 0.00026011999999999997 0 0.00026021999999999997 3.3 0.00026014 3.3 0.00026024 0 0.00026016 0 0.00026026 3.3 0.00026018 3.3 0.00026028 0 0.0002602 0 0.0002603 3.3 0.00026021999999999997 3.3 0.00026032 0 0.00026024 0 0.00026034 3.3 0.00026026 3.3 0.00026036 0 0.00026028 0 0.00026038 3.3 0.0002603 3.3 0.0002604 0 0.00026032 0 0.00026042 3.3 0.00026034 3.3 0.00026044 0 0.00026036 0 0.00026046 3.3 0.00026038 3.3 0.00026048 0 0.0002604 0 0.0002605 3.3 0.00026042 3.3 0.00026052 0 0.00026043999999999997 0 0.00026053999999999997 3.3 0.00026046 3.3 0.00026056 0 0.00026048 0 0.00026058 3.3 0.0002605 3.3 0.0002606 0 0.00026052 0 0.00026062 3.3 0.00026053999999999997 3.3 0.00026063999999999997 0 0.00026056 0 0.00026066 3.3 0.00026058 3.3 0.00026068 0 0.0002606 0 0.0002607 3.3 0.00026062 3.3 0.00026072 0 0.00026063999999999997 0 0.00026074 3.3 0.00026066 3.3 0.00026076 0 0.00026068 0 0.00026078 3.3 0.0002607 3.3 0.0002608 0 0.00026072 0 0.00026082 3.3 0.00026074 3.3 0.00026084 0 0.00026076 0 0.00026086 3.3 0.00026078 3.3 0.00026088 0 0.0002608 0 0.0002609 3.3 0.00026082 3.3 0.00026092 0 0.00026084 0 0.00026094 3.3 0.00026085999999999997 3.3 0.00026095999999999997 0 0.00026088 0 0.00026098 3.3 0.0002609 3.3 0.000261 0 0.00026092 0 0.00026102 3.3 0.00026094 3.3 0.00026104 0 0.00026095999999999997 0 0.00026105999999999997 3.3 0.00026098 3.3 0.00026108 0 0.000261 0 0.0002611 3.3 0.00026102 3.3 0.00026112 0 0.00026104 0 0.00026114 3.3 0.00026105999999999997 3.3 0.00026115999999999997 0 0.00026108 0 0.00026118 3.3 0.0002611 3.3 0.0002612 0 0.00026112 0 0.00026122 3.3 0.00026114 3.3 0.00026124 0 0.00026115999999999997 0 0.00026126 3.3 0.00026118 3.3 0.00026128 0 0.0002612 0 0.0002613 3.3 0.00026122 3.3 0.00026132 0 0.00026124 0 0.00026134 3.3 0.00026126 3.3 0.00026136 0 0.00026128 0 0.00026138 3.3 0.0002613 3.3 0.0002614 0 0.00026132 0 0.00026142 3.3 0.00026134 3.3 0.00026144 0 0.00026136 0 0.00026146 3.3 0.00026137999999999997 3.3 0.00026147999999999997 0 0.0002614 0 0.0002615 3.3 0.00026142 3.3 0.00026152 0 0.00026144 0 0.00026154 3.3 0.00026146 3.3 0.00026156 0 0.00026147999999999997 0 0.00026157999999999997 3.3 0.0002615 3.3 0.0002616 0 0.00026152 0 0.00026162 3.3 0.00026154 3.3 0.00026164 0 0.00026156 0 0.00026166 3.3 0.00026157999999999997 3.3 0.00026168 0 0.0002616 0 0.0002617 3.3 0.00026162 3.3 0.00026172 0 0.00026164 0 0.00026174 3.3 0.00026166 3.3 0.00026176 0 0.00026168 0 0.00026178 3.3 0.0002617 3.3 0.0002618 0 0.00026172 0 0.00026182 3.3 0.00026174 3.3 0.00026184 0 0.00026176 0 0.00026186 3.3 0.00026178 3.3 0.00026188 0 0.00026179999999999997 0 0.00026189999999999997 3.3 0.00026182 3.3 0.00026192 0 0.00026184 0 0.00026194 3.3 0.00026186 3.3 0.00026196 0 0.00026188 0 0.00026198 3.3 0.00026189999999999997 3.3 0.00026199999999999997 0 0.00026192 0 0.00026202 3.3 0.00026194 3.3 0.00026204 0 0.00026196 0 0.00026206 3.3 0.00026198 3.3 0.00026208 0 0.00026199999999999997 0 0.0002621 3.3 0.00026202 3.3 0.00026212 0 0.00026204 0 0.00026214 3.3 0.00026206 3.3 0.00026216 0 0.00026208 0 0.00026218 3.3 0.0002621 3.3 0.0002622 0 0.00026212 0 0.00026222 3.3 0.00026214 3.3 0.00026224 0 0.00026216 0 0.00026226 3.3 0.00026218 3.3 0.00026228 0 0.0002622 0 0.0002623 3.3 0.00026221999999999997 3.3 0.00026231999999999997 0 0.00026224 0 0.00026234 3.3 0.00026226 3.3 0.00026236 0 0.00026228 0 0.00026238 3.3 0.0002623 3.3 0.0002624 0 0.00026231999999999997 0 0.00026241999999999997 3.3 0.00026234 3.3 0.00026244 0 0.00026236 0 0.00026246 3.3 0.00026238 3.3 0.00026248 0 0.0002624 0 0.0002625 3.3 0.00026241999999999997 3.3 0.00026252 0 0.00026244 0 0.00026254 3.3 0.00026246 3.3 0.00026256 0 0.00026248 0 0.00026258 3.3 0.0002625 3.3 0.0002626 0 0.00026252 0 0.00026262 3.3 0.00026254 3.3 0.00026264 0 0.00026256 0 0.00026266 3.3 0.00026258 3.3 0.00026268 0 0.0002626 0 0.0002627 3.3 0.00026262 3.3 0.00026272 0 0.00026263999999999997 0 0.00026273999999999997 3.3 0.00026266 3.3 0.00026276 0 0.00026268 0 0.00026278 3.3 0.0002627 3.3 0.0002628 0 0.00026272 0 0.00026282 3.3 0.00026273999999999997 3.3 0.00026283999999999997 0 0.00026276 0 0.00026286 3.3 0.00026278 3.3 0.00026288 0 0.0002628 0 0.0002629 3.3 0.00026282 3.3 0.00026292 0 0.00026283999999999997 0 0.00026293999999999997 3.3 0.00026286 3.3 0.00026296 0 0.00026288 0 0.00026298 3.3 0.0002629 3.3 0.000263 0 0.00026292 0 0.00026302 3.3 0.00026293999999999997 3.3 0.00026304 0 0.00026296 0 0.00026306 3.3 0.00026298 3.3 0.00026308 0 0.000263 0 0.0002631 3.3 0.00026302 3.3 0.00026312 0 0.00026304 0 0.00026314 3.3 0.00026306 3.3 0.00026316 0 0.00026308 0 0.00026318 3.3 0.0002631 3.3 0.0002632 0 0.00026312 0 0.00026322 3.3 0.00026314 3.3 0.00026324 0 0.00026315999999999997 0 0.00026325999999999997 3.3 0.00026318 3.3 0.00026328 0 0.0002632 0 0.0002633 3.3 0.00026322 3.3 0.00026332 0 0.00026324 0 0.00026334 3.3 0.00026325999999999997 3.3 0.00026335999999999997 0 0.00026328 0 0.00026338 3.3 0.0002633 3.3 0.0002634 0 0.00026332 0 0.00026342 3.3 0.00026334 3.3 0.00026344 0 0.00026335999999999997 0 0.00026346 3.3 0.00026338 3.3 0.00026348 0 0.0002634 0 0.0002635 3.3 0.00026342 3.3 0.00026352 0 0.00026344 0 0.00026354 3.3 0.00026346 3.3 0.00026356 0 0.00026348 0 0.00026358 3.3 0.0002635 3.3 0.0002636 0 0.00026352 0 0.00026362 3.3 0.00026354 3.3 0.00026364 0 0.00026356 0 0.00026366 3.3 0.00026357999999999997 3.3 0.00026367999999999997 0 0.0002636 0 0.0002637 3.3 0.00026362 3.3 0.00026372 0 0.00026364 0 0.00026374 3.3 0.00026366 3.3 0.00026376 0 0.00026367999999999997 0 0.00026377999999999997 3.3 0.0002637 3.3 0.0002638 0 0.00026372 0 0.00026382 3.3 0.00026374 3.3 0.00026384 0 0.00026376 0 0.00026386 3.3 0.00026377999999999997 3.3 0.00026388 0 0.0002638 0 0.0002639 3.3 0.00026382 3.3 0.00026392 0 0.00026384 0 0.00026394 3.3 0.00026386 3.3 0.00026396 0 0.00026388 0 0.00026398 3.3 0.0002639 3.3 0.000264 0 0.00026392 0 0.00026402 3.3 0.00026394 3.3 0.00026404 0 0.00026396 0 0.00026406 3.3 0.00026398 3.3 0.00026408 0 0.00026399999999999997 0 0.00026409999999999997 3.3 0.00026402 3.3 0.00026412 0 0.00026404 0 0.00026414 3.3 0.00026406 3.3 0.00026416 0 0.00026408 0 0.00026418 3.3 0.00026409999999999997 3.3 0.00026419999999999997 0 0.00026412 0 0.00026422 3.3 0.00026414 3.3 0.00026424 0 0.00026416 0 0.00026426 3.3 0.00026418 3.3 0.00026428 0 0.00026419999999999997 0 0.0002643 3.3 0.00026422 3.3 0.00026432 0 0.00026424 0 0.00026434 3.3 0.00026426 3.3 0.00026436 0 0.00026428 0 0.00026438 3.3 0.0002643 3.3 0.0002644 0 0.00026432 0 0.00026442 3.3 0.00026434 3.3 0.00026444 0 0.00026436 0 0.00026446 3.3 0.00026438 3.3 0.00026448 0 0.0002644 0 0.0002645 3.3 0.00026441999999999997 3.3 0.00026451999999999997 0 0.00026444 0 0.00026454 3.3 0.00026446 3.3 0.00026456 0 0.00026448 0 0.00026458 3.3 0.0002645 3.3 0.0002646 0 0.00026451999999999997 0 0.00026461999999999997 3.3 0.00026454 3.3 0.00026464 0 0.00026456 0 0.00026466 3.3 0.00026458 3.3 0.00026468 0 0.0002646 0 0.0002647 3.3 0.00026461999999999997 3.3 0.00026471999999999997 0 0.00026464 0 0.00026474 3.3 0.00026466 3.3 0.00026476 0 0.00026468 0 0.00026478 3.3 0.0002647 3.3 0.0002648 0 0.00026471999999999997 0 0.00026482 3.3 0.00026474 3.3 0.00026484 0 0.00026476 0 0.00026486 3.3 0.00026478 3.3 0.00026488 0 0.0002648 0 0.0002649 3.3 0.00026482 3.3 0.00026492 0 0.00026484 0 0.00026494 3.3 0.00026486 3.3 0.00026496 0 0.00026488 0 0.00026498 3.3 0.0002649 3.3 0.000265 0 0.00026492 0 0.00026502 3.3 0.00026493999999999997 3.3 0.00026503999999999997 0 0.00026496 0 0.00026506 3.3 0.00026498 3.3 0.00026508 0 0.000265 0 0.0002651 3.3 0.00026502 3.3 0.00026512 0 0.00026503999999999997 0 0.00026513999999999997 3.3 0.00026506 3.3 0.00026516 0 0.00026508 0 0.00026518 3.3 0.0002651 3.3 0.0002652 0 0.00026512 0 0.00026522 3.3 0.00026513999999999997 3.3 0.00026524 0 0.00026516 0 0.00026526 3.3 0.00026518 3.3 0.00026528 0 0.0002652 0 0.0002653 3.3 0.00026522 3.3 0.00026532 0 0.00026524 0 0.00026534 3.3 0.00026526 3.3 0.00026536 0 0.00026528 0 0.00026538 3.3 0.0002653 3.3 0.0002654 0 0.00026532 0 0.00026542 3.3 0.00026534 3.3 0.00026544 0 0.00026535999999999997 0 0.00026545999999999997 3.3 0.00026538 3.3 0.00026548 0 0.0002654 0 0.0002655 3.3 0.00026542 3.3 0.00026552 0 0.00026544 0 0.00026554 3.3 0.00026545999999999997 3.3 0.00026555999999999997 0 0.00026548 0 0.00026558 3.3 0.0002655 3.3 0.0002656 0 0.00026552 0 0.00026562 3.3 0.00026554 3.3 0.00026564 0 0.00026555999999999997 0 0.00026566 3.3 0.00026558 3.3 0.00026568 0 0.0002656 0 0.0002657 3.3 0.00026562 3.3 0.00026572 0 0.00026564 0 0.00026574 3.3 0.00026566 3.3 0.00026576 0 0.00026568 0 0.00026578 3.3 0.0002657 3.3 0.0002658 0 0.00026572 0 0.00026582 3.3 0.00026574 3.3 0.00026584 0 0.00026576 0 0.00026586 3.3 0.00026577999999999997 3.3 0.00026587999999999997 0 0.0002658 0 0.0002659 3.3 0.00026582 3.3 0.00026592 0 0.00026584 0 0.00026594 3.3 0.00026586 3.3 0.00026596 0 0.00026587999999999997 0 0.00026597999999999997 3.3 0.0002659 3.3 0.000266 0 0.00026592 0 0.00026602 3.3 0.00026594 3.3 0.00026604 0 0.00026596 0 0.00026606 3.3 0.00026597999999999997 3.3 0.00026608 0 0.000266 0 0.0002661 3.3 0.00026602 3.3 0.00026612 0 0.00026604 0 0.00026614 3.3 0.00026606 3.3 0.00026616 0 0.00026608 0 0.00026618 3.3 0.0002661 3.3 0.0002662 0 0.00026612 0 0.00026622 3.3 0.00026614 3.3 0.00026624 0 0.00026616 0 0.00026626 3.3 0.00026618 3.3 0.00026628 0 0.00026619999999999997 0 0.00026629999999999997 3.3 0.00026622 3.3 0.00026632 0 0.00026624 0 0.00026634 3.3 0.00026626 3.3 0.00026636 0 0.00026628 0 0.00026638 3.3 0.00026629999999999997 3.3 0.00026639999999999997 0 0.00026632 0 0.00026642 3.3 0.00026634 3.3 0.00026644 0 0.00026636 0 0.00026646 3.3 0.00026638 3.3 0.00026648 0 0.00026639999999999997 0 0.00026649999999999997 3.3 0.00026642 3.3 0.00026652 0 0.00026644 0 0.00026654 3.3 0.00026646 3.3 0.00026656 0 0.00026648 0 0.00026658 3.3 0.00026649999999999997 3.3 0.0002666 0 0.00026652 0 0.00026662 3.3 0.00026654 3.3 0.00026664 0 0.00026656 0 0.00026666 3.3 0.00026658 3.3 0.00026668 0 0.0002666 0 0.0002667 3.3 0.00026662 3.3 0.00026672 0 0.00026664 0 0.00026674 3.3 0.00026666 3.3 0.00026676 0 0.00026668 0 0.00026678 3.3 0.0002667 3.3 0.0002668 0 0.00026671999999999997 0 0.00026681999999999997 3.3 0.00026674 3.3 0.00026684 0 0.00026676 0 0.00026686 3.3 0.00026678 3.3 0.00026688 0 0.0002668 0 0.0002669 3.3 0.00026681999999999997 3.3 0.00026691999999999997 0 0.00026684 0 0.00026694 3.3 0.00026686 3.3 0.00026696 0 0.00026688 0 0.00026698 3.3 0.0002669 3.3 0.000267 0 0.00026691999999999997 0 0.00026702 3.3 0.00026694 3.3 0.00026704 0 0.00026696 0 0.00026706 3.3 0.00026698 3.3 0.00026708 0 0.000267 0 0.0002671 3.3 0.00026702 3.3 0.00026712 0 0.00026704 0 0.00026714 3.3 0.00026706 3.3 0.00026716 0 0.00026708 0 0.00026718 3.3 0.0002671 3.3 0.0002672 0 0.00026712 0 0.00026722 3.3 0.00026713999999999997 3.3 0.00026723999999999997 0 0.00026716 0 0.00026726 3.3 0.00026718 3.3 0.00026728 0 0.0002672 0 0.0002673 3.3 0.00026722 3.3 0.00026732 0 0.00026723999999999997 0 0.00026733999999999997 3.3 0.00026726 3.3 0.00026736 0 0.00026728 0 0.00026738 3.3 0.0002673 3.3 0.0002674 0 0.00026732 0 0.00026742 3.3 0.00026733999999999997 3.3 0.00026744 0 0.00026736 0 0.00026746 3.3 0.00026738 3.3 0.00026748 0 0.0002674 0 0.0002675 3.3 0.00026742 3.3 0.00026752 0 0.00026744 0 0.00026754 3.3 0.00026746 3.3 0.00026756 0 0.00026748 0 0.00026758 3.3 0.0002675 3.3 0.0002676 0 0.00026752 0 0.00026762 3.3 0.00026754 3.3 0.00026764 0 0.00026755999999999997 0 0.00026765999999999997 3.3 0.00026758 3.3 0.00026768 0 0.0002676 0 0.0002677 3.3 0.00026762 3.3 0.00026772 0 0.00026764 0 0.00026774 3.3 0.00026765999999999997 3.3 0.00026775999999999997 0 0.00026768 0 0.00026778 3.3 0.0002677 3.3 0.0002678 0 0.00026772 0 0.00026782 3.3 0.00026774 3.3 0.00026784 0 0.00026775999999999997 0 0.00026786 3.3 0.00026778 3.3 0.00026788 0 0.0002678 0 0.0002679 3.3 0.00026782 3.3 0.00026792 0 0.00026784 0 0.00026794 3.3 0.00026786 3.3 0.00026796 0 0.00026788 0 0.00026798 3.3 0.0002679 3.3 0.000268 0 0.00026792 0 0.00026802 3.3 0.00026794 3.3 0.00026804 0 0.00026796 0 0.00026806 3.3 0.00026797999999999997 3.3 0.00026807999999999997 0 0.000268 0 0.0002681 3.3 0.00026802 3.3 0.00026812 0 0.00026804 0 0.00026814 3.3 0.00026806 3.3 0.00026816 0 0.00026807999999999997 0 0.00026817999999999997 3.3 0.0002681 3.3 0.0002682 0 0.00026812 0 0.00026822 3.3 0.00026814 3.3 0.00026824 0 0.00026816 0 0.00026826 3.3 0.00026817999999999997 3.3 0.00026827999999999997 0 0.0002682 0 0.0002683 3.3 0.00026822 3.3 0.00026832 0 0.00026824 0 0.00026834 3.3 0.00026826 3.3 0.00026836 0 0.00026827999999999997 0 0.00026838 3.3 0.0002683 3.3 0.0002684 0 0.00026832 0 0.00026842 3.3 0.00026834 3.3 0.00026844 0 0.00026836 0 0.00026846 3.3 0.00026838 3.3 0.00026848 0 0.0002684 0 0.0002685 3.3 0.00026842 3.3 0.00026852 0 0.00026844 0 0.00026854 3.3 0.00026846 3.3 0.00026856 0 0.00026848 0 0.00026858 3.3 0.00026849999999999997 3.3 0.00026859999999999997 0 0.00026852 0 0.00026862 3.3 0.00026854 3.3 0.00026864 0 0.00026856 0 0.00026866 3.3 0.00026858 3.3 0.00026868 0 0.00026859999999999997 0 0.00026869999999999997 3.3 0.00026862 3.3 0.00026872 0 0.00026864 0 0.00026874 3.3 0.00026866 3.3 0.00026876 0 0.00026868 0 0.00026878 3.3 0.00026869999999999997 3.3 0.0002688 0 0.00026872 0 0.00026882 3.3 0.00026874 3.3 0.00026884 0 0.00026876 0 0.00026886 3.3 0.00026878 3.3 0.00026888 0 0.0002688 0 0.0002689 3.3 0.00026882 3.3 0.00026892 0 0.00026884 0 0.00026894 3.3 0.00026886 3.3 0.00026896 0 0.00026888 0 0.00026898 3.3 0.0002689 3.3 0.000269 0 0.00026891999999999997 0 0.00026901999999999997 3.3 0.00026894 3.3 0.00026904 0 0.00026896 0 0.00026906 3.3 0.00026898 3.3 0.00026908 0 0.000269 0 0.0002691 3.3 0.00026901999999999997 3.3 0.00026911999999999997 0 0.00026904 0 0.00026914 3.3 0.00026906 3.3 0.00026916 0 0.00026908 0 0.00026918 3.3 0.0002691 3.3 0.0002692 0 0.00026911999999999997 0 0.00026922 3.3 0.00026914 3.3 0.00026924 0 0.00026916 0 0.00026926 3.3 0.00026918 3.3 0.00026928 0 0.0002692 0 0.0002693 3.3 0.00026922 3.3 0.00026932 0 0.00026924 0 0.00026934 3.3 0.00026926 3.3 0.00026936 0 0.00026928 0 0.00026938 3.3 0.0002693 3.3 0.0002694 0 0.00026932 0 0.00026942 3.3 0.00026933999999999997 3.3 0.00026943999999999997 0 0.00026936 0 0.00026946 3.3 0.00026938 3.3 0.00026948 0 0.0002694 0 0.0002695 3.3 0.00026942 3.3 0.00026952 0 0.00026943999999999997 0 0.00026953999999999997 3.3 0.00026946 3.3 0.00026956 0 0.00026948 0 0.00026958 3.3 0.0002695 3.3 0.0002696 0 0.00026952 0 0.00026962 3.3 0.00026953999999999997 3.3 0.00026964 0 0.00026956 0 0.00026966 3.3 0.00026958 3.3 0.00026968 0 0.0002696 0 0.0002697 3.3 0.00026962 3.3 0.00026972 0 0.00026964 0 0.00026974 3.3 0.00026966 3.3 0.00026976 0 0.00026968 0 0.00026978 3.3 0.0002697 3.3 0.0002698 0 0.00026972 0 0.00026982 3.3 0.00026974 3.3 0.00026984 0 0.00026975999999999997 0 0.00026985999999999997 3.3 0.00026978 3.3 0.00026988 0 0.0002698 0 0.0002699 3.3 0.00026982 3.3 0.00026992 0 0.00026984 0 0.00026994 3.3 0.00026985999999999997 3.3 0.00026995999999999997 0 0.00026988 0 0.00026998 3.3 0.0002699 3.3 0.00027 0 0.00026992 0 0.00027002 3.3 0.00026994 3.3 0.00027004 0 0.00026995999999999997 0 0.00027005999999999997 3.3 0.00026998 3.3 0.00027008 0 0.00027 0 0.0002701 3.3 0.00027002 3.3 0.00027012 0 0.00027004 0 0.00027014 3.3 0.00027005999999999997 3.3 0.00027016 0 0.00027008 0 0.00027018 3.3 0.0002701 3.3 0.0002702 0 0.00027012 0 0.00027022 3.3 0.00027014 3.3 0.00027024 0 0.00027016 0 0.00027026 3.3 0.00027018 3.3 0.00027028 0 0.0002702 0 0.0002703 3.3 0.00027022 3.3 0.00027032 0 0.00027024 0 0.00027034 3.3 0.00027026 3.3 0.00027036 0 0.00027027999999999997 0 0.00027037999999999997 3.3 0.0002703 3.3 0.0002704 0 0.00027032 0 0.00027042 3.3 0.00027034 3.3 0.00027044 0 0.00027036 0 0.00027046 3.3 0.00027037999999999997 3.3 0.00027047999999999997 0 0.0002704 0 0.0002705 3.3 0.00027042 3.3 0.00027052 0 0.00027044 0 0.00027054 3.3 0.00027046 3.3 0.00027056 0 0.00027047999999999997 0 0.00027058 3.3 0.0002705 3.3 0.0002706 0 0.00027052 0 0.00027062 3.3 0.00027054 3.3 0.00027064 0 0.00027056 0 0.00027066 3.3 0.00027058 3.3 0.00027068 0 0.0002706 0 0.0002707 3.3 0.00027062 3.3 0.00027072 0 0.00027064 0 0.00027074 3.3 0.00027066 3.3 0.00027076 0 0.00027068 0 0.00027078 3.3 0.00027069999999999997 3.3 0.00027079999999999997 0 0.00027072 0 0.00027082 3.3 0.00027074 3.3 0.00027084 0 0.00027076 0 0.00027086 3.3 0.00027078 3.3 0.00027088 0 0.00027079999999999997 0 0.00027089999999999997 3.3 0.00027082 3.3 0.00027092 0 0.00027084 0 0.00027094 3.3 0.00027086 3.3 0.00027096 0 0.00027088 0 0.00027098 3.3 0.00027089999999999997 3.3 0.000271 0 0.00027092 0 0.00027102 3.3 0.00027094 3.3 0.00027104 0 0.00027096 0 0.00027106 3.3 0.00027098 3.3 0.00027108 0 0.000271 0 0.0002711 3.3 0.00027102 3.3 0.00027112 0 0.00027104 0 0.00027114 3.3 0.00027106 3.3 0.00027116 0 0.00027108 0 0.00027118 3.3 0.0002711 3.3 0.0002712 0 0.00027111999999999997 0 0.00027121999999999997 3.3 0.00027114 3.3 0.00027124 0 0.00027116 0 0.00027126 3.3 0.00027118 3.3 0.00027128 0 0.0002712 0 0.0002713 3.3 0.00027121999999999997 3.3 0.00027131999999999997 0 0.00027124 0 0.00027134 3.3 0.00027126 3.3 0.00027136 0 0.00027128 0 0.00027138 3.3 0.0002713 3.3 0.0002714 0 0.00027131999999999997 0 0.00027142 3.3 0.00027134 3.3 0.00027144 0 0.00027136 0 0.00027146 3.3 0.00027138 3.3 0.00027148 0 0.0002714 0 0.0002715 3.3 0.00027142 3.3 0.00027152 0 0.00027144 0 0.00027154 3.3 0.00027146 3.3 0.00027156 0 0.00027148 0 0.00027158 3.3 0.0002715 3.3 0.0002716 0 0.00027152 0 0.00027162 3.3 0.00027154 3.3 0.00027164 0 0.00027156 0 0.00027166 3.3 0.00027158 3.3 0.00027168 0 0.0002716 0 0.0002717 3.3 0.00027162 3.3 0.00027172 0 0.00027163999999999997 0 0.00027173999999999997 3.3 0.00027166 3.3 0.00027176 0 0.00027168 0 0.00027178 3.3 0.0002717 3.3 0.0002718 0 0.00027172 0 0.00027182 3.3 0.00027173999999999997 3.3 0.00027183999999999997 0 0.00027176 0 0.00027186 3.3 0.00027178 3.3 0.00027188 0 0.0002718 0 0.0002719 3.3 0.00027182 3.3 0.00027192 0 0.00027183999999999997 0 0.00027194 3.3 0.00027186 3.3 0.00027196 0 0.00027188 0 0.00027198 3.3 0.0002719 3.3 0.000272 0 0.00027192 0 0.00027202 3.3 0.00027194 3.3 0.00027204 0 0.00027196 0 0.00027206 3.3 0.00027198 3.3 0.00027208 0 0.000272 0 0.0002721 3.3 0.00027202 3.3 0.00027212 0 0.00027204 0 0.00027214 3.3 0.00027205999999999997 3.3 0.00027215999999999997 0 0.00027208 0 0.00027218 3.3 0.0002721 3.3 0.0002722 0 0.00027212 0 0.00027222 3.3 0.00027214 3.3 0.00027224 0 0.00027215999999999997 0 0.00027225999999999997 3.3 0.00027218 3.3 0.00027228 0 0.0002722 0 0.0002723 3.3 0.00027222 3.3 0.00027232 0 0.00027224 0 0.00027234 3.3 0.00027225999999999997 3.3 0.00027236 0 0.00027228 0 0.00027238 3.3 0.0002723 3.3 0.0002724 0 0.00027232 0 0.00027242 3.3 0.00027234 3.3 0.00027244 0 0.00027236 0 0.00027246 3.3 0.00027238 3.3 0.00027248 0 0.0002724 0 0.0002725 3.3 0.00027242 3.3 0.00027252 0 0.00027244 0 0.00027254 3.3 0.00027246 3.3 0.00027256 0 0.00027247999999999997 0 0.00027257999999999997 3.3 0.0002725 3.3 0.0002726 0 0.00027252 0 0.00027262 3.3 0.00027254 3.3 0.00027264 0 0.00027256 0 0.00027266 3.3 0.00027257999999999997 3.3 0.00027267999999999997 0 0.0002726 0 0.0002727 3.3 0.00027262 3.3 0.00027272 0 0.00027264 0 0.00027274 3.3 0.00027266 3.3 0.00027276 0 0.00027267999999999997 0 0.00027278 3.3 0.0002727 3.3 0.0002728 0 0.00027272 0 0.00027282 3.3 0.00027274 3.3 0.00027284 0 0.00027276 0 0.00027286 3.3 0.00027278 3.3 0.00027288 0 0.0002728 0 0.0002729 3.3 0.00027282 3.3 0.00027292 0 0.00027284 0 0.00027294 3.3 0.00027286 3.3 0.00027296 0 0.00027288 0 0.00027298 3.3 0.00027289999999999997 3.3 0.00027299999999999997 0 0.00027292 0 0.00027302 3.3 0.00027294 3.3 0.00027304 0 0.00027296 0 0.00027306 3.3 0.00027298 3.3 0.00027308 0 0.00027299999999999997 0 0.00027309999999999997 3.3 0.00027302 3.3 0.00027312 0 0.00027304 0 0.00027314 3.3 0.00027306 3.3 0.00027316 0 0.00027308 0 0.00027318 3.3 0.00027309999999999997 3.3 0.00027319999999999997 0 0.00027312 0 0.00027322 3.3 0.00027314 3.3 0.00027324 0 0.00027316 0 0.00027326 3.3 0.00027318 3.3 0.00027328 0 0.00027319999999999997 0 0.0002733 3.3 0.00027322 3.3 0.00027332 0 0.00027324 0 0.00027334 3.3 0.00027326 3.3 0.00027336 0 0.00027328 0 0.00027338 3.3 0.0002733 3.3 0.0002734 0 0.00027332 0 0.00027342 3.3 0.00027334 3.3 0.00027344 0 0.00027336 0 0.00027346 3.3 0.00027338 3.3 0.00027348 0 0.0002734 0 0.0002735 3.3 0.00027341999999999997 3.3 0.00027351999999999997 0 0.00027344 0 0.00027354 3.3 0.00027346 3.3 0.00027356 0 0.00027348 0 0.00027358 3.3 0.0002735 3.3 0.0002736 0 0.00027351999999999997 0 0.00027361999999999997 3.3 0.00027354 3.3 0.00027364 0 0.00027356 0 0.00027366 3.3 0.00027358 3.3 0.00027368 0 0.0002736 0 0.0002737 3.3 0.00027361999999999997 3.3 0.00027372 0 0.00027364 0 0.00027374 3.3 0.00027366 3.3 0.00027376 0 0.00027368 0 0.00027378 3.3 0.0002737 3.3 0.0002738 0 0.00027372 0 0.00027382 3.3 0.00027374 3.3 0.00027384 0 0.00027376 0 0.00027386 3.3 0.00027378 3.3 0.00027388 0 0.0002738 0 0.0002739 3.3 0.00027382 3.3 0.00027392 0 0.00027383999999999997 0 0.00027393999999999997 3.3 0.00027386 3.3 0.00027396 0 0.00027388 0 0.00027398 3.3 0.0002739 3.3 0.000274 0 0.00027392 0 0.00027402 3.3 0.00027393999999999997 3.3 0.00027403999999999997 0 0.00027396 0 0.00027406 3.3 0.00027398 3.3 0.00027408 0 0.000274 0 0.0002741 3.3 0.00027402 3.3 0.00027412 0 0.00027403999999999997 0 0.00027414 3.3 0.00027406 3.3 0.00027416 0 0.00027408 0 0.00027418 3.3 0.0002741 3.3 0.0002742 0 0.00027412 0 0.00027422 3.3 0.00027414 3.3 0.00027424 0 0.00027416 0 0.00027426 3.3 0.00027418 3.3 0.00027428 0 0.0002742 0 0.0002743 3.3 0.00027422 3.3 0.00027432 0 0.00027424 0 0.00027434 3.3 0.00027425999999999997 3.3 0.00027435999999999997 0 0.00027428 0 0.00027438 3.3 0.0002743 3.3 0.0002744 0 0.00027432 0 0.00027442 3.3 0.00027434 3.3 0.00027444 0 0.00027435999999999997 0 0.00027445999999999997 3.3 0.00027438 3.3 0.00027448 0 0.0002744 0 0.0002745 3.3 0.00027442 3.3 0.00027452 0 0.00027444 0 0.00027454 3.3 0.00027445999999999997 3.3 0.00027456 0 0.00027448 0 0.00027458 3.3 0.0002745 3.3 0.0002746 0 0.00027452 0 0.00027462 3.3 0.00027454 3.3 0.00027464 0 0.00027456 0 0.00027466 3.3 0.00027458 3.3 0.00027468 0 0.0002746 0 0.0002747 3.3 0.00027462 3.3 0.00027472 0 0.00027464 0 0.00027474 3.3 0.00027466 3.3 0.00027476 0 0.00027467999999999997 0 0.00027477999999999997 3.3 0.0002747 3.3 0.0002748 0 0.00027472 0 0.00027482 3.3 0.00027474 3.3 0.00027484 0 0.00027476 0 0.00027486 3.3 0.00027477999999999997 3.3 0.00027487999999999997 0 0.0002748 0 0.0002749 3.3 0.00027482 3.3 0.00027492 0 0.00027484 0 0.00027494 3.3 0.00027486 3.3 0.00027496 0 0.00027487999999999997 0 0.00027497999999999997 3.3 0.0002749 3.3 0.000275 0 0.00027492 0 0.00027502 3.3 0.00027494 3.3 0.00027504 0 0.00027496 0 0.00027506 3.3 0.00027497999999999997 3.3 0.00027508 0 0.000275 0 0.0002751 3.3 0.00027502 3.3 0.00027512 0 0.00027504 0 0.00027514 3.3 0.00027506 3.3 0.00027516 0 0.00027508 0 0.00027518 3.3 0.0002751 3.3 0.0002752 0 0.00027512 0 0.00027522 3.3 0.00027514 3.3 0.00027524 0 0.00027516 0 0.00027526 3.3 0.00027518 3.3 0.00027528 0 0.00027519999999999997 0 0.00027529999999999997 3.3 0.00027522 3.3 0.00027532 0 0.00027524 0 0.00027534 3.3 0.00027526 3.3 0.00027536 0 0.00027528 0 0.00027538 3.3 0.00027529999999999997 3.3 0.00027539999999999997 0 0.00027532 0 0.00027542 3.3 0.00027534 3.3 0.00027544 0 0.00027536 0 0.00027546 3.3 0.00027538 3.3 0.00027548 0 0.00027539999999999997 0 0.0002755 3.3 0.00027542 3.3 0.00027552 0 0.00027544 0 0.00027554 3.3 0.00027546 3.3 0.00027556 0 0.00027548 0 0.00027558 3.3 0.0002755 3.3 0.0002756 0 0.00027552 0 0.00027562 3.3 0.00027554 3.3 0.00027564 0 0.00027556 0 0.00027566 3.3 0.00027558 3.3 0.00027568 0 0.0002756 0 0.0002757 3.3 0.00027561999999999997 3.3 0.00027571999999999997 0 0.00027564 0 0.00027574 3.3 0.00027566 3.3 0.00027576 0 0.00027568 0 0.00027578 3.3 0.0002757 3.3 0.0002758 0 0.00027571999999999997 0 0.00027581999999999997 3.3 0.00027574 3.3 0.00027584 0 0.00027576 0 0.00027586 3.3 0.00027578 3.3 0.00027588 0 0.0002758 0 0.0002759 3.3 0.00027581999999999997 3.3 0.00027592 0 0.00027584 0 0.00027594 3.3 0.00027586 3.3 0.00027596 0 0.00027588 0 0.00027598 3.3 0.0002759 3.3 0.000276 0 0.00027592 0 0.00027602 3.3 0.00027594 3.3 0.00027604 0 0.00027596 0 0.00027606 3.3 0.00027598 3.3 0.00027608 0 0.000276 0 0.0002761 3.3 0.00027602 3.3 0.00027612 0 0.00027603999999999997 0 0.00027613999999999997 3.3 0.00027606 3.3 0.00027616 0 0.00027608 0 0.00027618 3.3 0.0002761 3.3 0.0002762 0 0.00027612 0 0.00027622 3.3 0.00027613999999999997 3.3 0.00027623999999999997 0 0.00027616 0 0.00027626 3.3 0.00027618 3.3 0.00027628 0 0.0002762 0 0.0002763 3.3 0.00027622 3.3 0.00027632 0 0.00027623999999999997 0 0.00027634 3.3 0.00027626 3.3 0.00027636 0 0.00027628 0 0.00027638 3.3 0.0002763 3.3 0.0002764 0 0.00027632 0 0.00027642 3.3 0.00027634 3.3 0.00027644 0 0.00027636 0 0.00027646 3.3 0.00027638 3.3 0.00027648 0 0.0002764 0 0.0002765 3.3 0.00027642 3.3 0.00027652 0 0.00027644 0 0.00027654 3.3 0.00027645999999999997 3.3 0.00027655999999999997 0 0.00027648 0 0.00027658 3.3 0.0002765 3.3 0.0002766 0 0.00027652 0 0.00027662 3.3 0.00027654 3.3 0.00027664 0 0.00027655999999999997 0 0.00027665999999999997 3.3 0.00027658 3.3 0.00027668 0 0.0002766 0 0.0002767 3.3 0.00027662 3.3 0.00027672 0 0.00027664 0 0.00027674 3.3 0.00027665999999999997 3.3 0.00027675999999999997 0 0.00027668 0 0.00027678 3.3 0.0002767 3.3 0.0002768 0 0.00027672 0 0.00027682 3.3 0.00027674 3.3 0.00027684 0 0.00027675999999999997 0 0.00027686 3.3 0.00027678 3.3 0.00027688 0 0.0002768 0 0.0002769 3.3 0.00027682 3.3 0.00027692 0 0.00027684 0 0.00027694 3.3 0.00027686 3.3 0.00027696 0 0.00027688 0 0.00027698 3.3 0.0002769 3.3 0.000277 0 0.00027692 0 0.00027702 3.3 0.00027694 3.3 0.00027704 0 0.00027696 0 0.00027706 3.3 0.00027697999999999997 3.3 0.00027707999999999997 0 0.000277 0 0.0002771 3.3 0.00027702 3.3 0.00027712 0 0.00027704 0 0.00027714 3.3 0.00027706 3.3 0.00027716 0 0.00027707999999999997 0 0.00027717999999999997 3.3 0.0002771 3.3 0.0002772 0 0.00027712 0 0.00027722 3.3 0.00027714 3.3 0.00027724 0 0.00027716 0 0.00027726 3.3 0.00027717999999999997 3.3 0.00027728 0 0.0002772 0 0.0002773 3.3 0.00027722 3.3 0.00027732 0 0.00027724 0 0.00027734 3.3 0.00027726 3.3 0.00027736 0 0.00027728 0 0.00027738 3.3 0.0002773 3.3 0.0002774 0 0.00027732 0 0.00027742 3.3 0.00027734 3.3 0.00027744 0 0.00027736 0 0.00027746 3.3 0.00027738 3.3 0.00027748 0 0.00027739999999999997 0 0.00027749999999999997 3.3 0.00027742 3.3 0.00027752 0 0.00027744 0 0.00027754 3.3 0.00027746 3.3 0.00027756 0 0.00027748 0 0.00027758 3.3 0.00027749999999999997 3.3 0.00027759999999999997 0 0.00027752 0 0.00027762 3.3 0.00027754 3.3 0.00027764 0 0.00027756 0 0.00027766 3.3 0.00027758 3.3 0.00027768 0 0.00027759999999999997 0 0.0002777 3.3 0.00027762 3.3 0.00027772 0 0.00027764 0 0.00027774 3.3 0.00027766 3.3 0.00027776 0 0.00027768 0 0.00027778 3.3 0.0002777 3.3 0.0002778 0 0.00027772 0 0.00027782 3.3 0.00027774 3.3 0.00027784 0 0.00027776 0 0.00027786 3.3 0.00027778 3.3 0.00027788 0 0.0002778 0 0.0002779 3.3 0.00027781999999999997 3.3 0.00027791999999999997 0 0.00027784 0 0.00027794 3.3 0.00027786 3.3 0.00027796 0 0.00027788 0 0.00027798 3.3 0.0002779 3.3 0.000278 0 0.00027791999999999997 0 0.00027801999999999997 3.3 0.00027794 3.3 0.00027804 0 0.00027796 0 0.00027806 3.3 0.00027798 3.3 0.00027808 0 0.000278 0 0.0002781 3.3 0.00027801999999999997 3.3 0.00027812 0 0.00027804 0 0.00027814 3.3 0.00027806 3.3 0.00027816 0 0.00027808 0 0.00027818 3.3 0.0002781 3.3 0.0002782 0 0.00027812 0 0.00027822 3.3 0.00027814 3.3 0.00027824 0 0.00027816 0 0.00027826 3.3 0.00027818 3.3 0.00027828 0 0.0002782 0 0.0002783 3.3 0.00027822 3.3 0.00027832 0 0.00027823999999999997 0 0.00027833999999999997 3.3 0.00027826 3.3 0.00027836 0 0.00027828 0 0.00027838 3.3 0.0002783 3.3 0.0002784 0 0.00027832 0 0.00027842 3.3 0.00027833999999999997 3.3 0.00027843999999999997 0 0.00027836 0 0.00027846 3.3 0.00027838 3.3 0.00027848 0 0.0002784 0 0.0002785 3.3 0.00027842 3.3 0.00027852 0 0.00027843999999999997 0 0.00027853999999999997 3.3 0.00027846 3.3 0.00027856 0 0.00027848 0 0.00027858 3.3 0.0002785 3.3 0.0002786 0 0.00027852 0 0.00027862 3.3 0.00027853999999999997 3.3 0.00027864 0 0.00027856 0 0.00027866 3.3 0.00027858 3.3 0.00027868 0 0.0002786 0 0.0002787 3.3 0.00027862 3.3 0.00027872 0 0.00027864 0 0.00027874 3.3 0.00027866 3.3 0.00027876 0 0.00027868 0 0.00027878 3.3 0.0002787 3.3 0.0002788 0 0.00027872 0 0.00027882 3.3 0.00027874 3.3 0.00027884 0 0.00027875999999999997 0 0.00027885999999999997 3.3 0.00027878 3.3 0.00027888 0 0.0002788 0 0.0002789 3.3 0.00027882 3.3 0.00027892 0 0.00027884 0 0.00027894 3.3 0.00027885999999999997 3.3 0.00027895999999999997 0 0.00027888 0 0.00027898 3.3 0.0002789 3.3 0.000279 0 0.00027892 0 0.00027902 3.3 0.00027894 3.3 0.00027904 0 0.00027895999999999997 0 0.00027906 3.3 0.00027898 3.3 0.00027908 0 0.000279 0 0.0002791 3.3 0.00027902 3.3 0.00027912 0 0.00027904 0 0.00027914 3.3 0.00027906 3.3 0.00027916 0 0.00027908 0 0.00027918 3.3 0.0002791 3.3 0.0002792 0 0.00027912 0 0.00027922 3.3 0.00027914 3.3 0.00027924 0 0.00027916 0 0.00027926 3.3 0.00027917999999999997 3.3 0.00027927999999999997 0 0.0002792 0 0.0002793 3.3 0.00027922 3.3 0.00027932 0 0.00027924 0 0.00027934 3.3 0.00027926 3.3 0.00027936 0 0.00027927999999999997 0 0.00027937999999999997 3.3 0.0002793 3.3 0.0002794 0 0.00027932 0 0.00027942 3.3 0.00027934 3.3 0.00027944 0 0.00027936 0 0.00027946 3.3 0.00027937999999999997 3.3 0.00027948 0 0.0002794 0 0.0002795 3.3 0.00027942 3.3 0.00027952 0 0.00027944 0 0.00027954 3.3 0.00027946 3.3 0.00027956 0 0.00027948 0 0.00027958 3.3 0.0002795 3.3 0.0002796 0 0.00027952 0 0.00027962 3.3 0.00027954 3.3 0.00027964 0 0.00027956 0 0.00027966 3.3 0.00027958 3.3 0.00027968 0 0.00027959999999999997 0 0.00027969999999999997 3.3 0.00027962 3.3 0.00027972 0 0.00027964 0 0.00027974 3.3 0.00027966 3.3 0.00027976 0 0.00027968 0 0.00027978 3.3 0.00027969999999999997 3.3 0.00027979999999999997 0 0.00027972 0 0.00027982 3.3 0.00027974 3.3 0.00027984 0 0.00027976 0 0.00027986 3.3 0.00027978 3.3 0.00027988 0 0.00027979999999999997 0 0.0002799 3.3 0.00027982 3.3 0.00027992 0 0.00027984 0 0.00027994 3.3 0.00027986 3.3 0.00027996 0 0.00027988 0 0.00027998 3.3 0.0002799 3.3 0.00028 0 0.00027992 0 0.00028002 3.3 0.00027994 3.3 0.00028004 0 0.00027996 0 0.00028006 3.3 0.00027998 3.3 0.00028008 0 0.00028 0 0.0002801 3.3 0.00028001999999999997 3.3 0.00028011999999999997 0 0.00028004 0 0.00028014 3.3 0.00028006 3.3 0.00028016 0 0.00028008 0 0.00028018 3.3 0.0002801 3.3 0.0002802 0 0.00028011999999999997 0 0.00028021999999999997 3.3 0.00028014 3.3 0.00028024 0 0.00028016 0 0.00028026 3.3 0.00028018 3.3 0.00028028 0 0.0002802 0 0.0002803 3.3 0.00028021999999999997 3.3 0.00028031999999999997 0 0.00028024 0 0.00028034 3.3 0.00028026 3.3 0.00028036 0 0.00028028 0 0.00028038 3.3 0.0002803 3.3 0.0002804 0 0.00028031999999999997 0 0.00028042 3.3 0.00028034 3.3 0.00028044 0 0.00028036 0 0.00028046 3.3 0.00028038 3.3 0.00028048 0 0.0002804 0 0.0002805 3.3 0.00028042 3.3 0.00028052 0 0.00028044 0 0.00028054 3.3 0.00028046 3.3 0.00028056 0 0.00028048 0 0.00028058 3.3 0.0002805 3.3 0.0002806 0 0.00028052 0 0.00028062 3.3 0.00028053999999999997 3.3 0.00028063999999999997 0 0.00028056 0 0.00028066 3.3 0.00028058 3.3 0.00028068 0 0.0002806 0 0.0002807 3.3 0.00028062 3.3 0.00028072 0 0.00028063999999999997 0 0.00028073999999999997 3.3 0.00028066 3.3 0.00028076 0 0.00028068 0 0.00028078 3.3 0.0002807 3.3 0.0002808 0 0.00028072 0 0.00028082 3.3 0.00028073999999999997 3.3 0.00028084 0 0.00028076 0 0.00028086 3.3 0.00028078 3.3 0.00028088 0 0.0002808 0 0.0002809 3.3 0.00028082 3.3 0.00028092 0 0.00028084 0 0.00028094 3.3 0.00028086 3.3 0.00028096 0 0.00028088 0 0.00028098 3.3 0.0002809 3.3 0.000281 0 0.00028092 0 0.00028102 3.3 0.00028094 3.3 0.00028104 0 0.00028095999999999997 0 0.00028105999999999997 3.3 0.00028098 3.3 0.00028108 0 0.000281 0 0.0002811 3.3 0.00028102 3.3 0.00028112 0 0.00028104 0 0.00028114 3.3 0.00028105999999999997 3.3 0.00028115999999999997 0 0.00028108 0 0.00028118 3.3 0.0002811 3.3 0.0002812 0 0.00028112 0 0.00028122 3.3 0.00028114 3.3 0.00028124 0 0.00028115999999999997 0 0.00028126 3.3 0.00028118 3.3 0.00028128 0 0.0002812 0 0.0002813 3.3 0.00028122 3.3 0.00028132 0 0.00028124 0 0.00028134 3.3 0.00028126 3.3 0.00028136 0 0.00028128 0 0.00028138 3.3 0.0002813 3.3 0.0002814 0 0.00028132 0 0.00028142 3.3 0.00028134 3.3 0.00028144 0 0.00028136 0 0.00028146 3.3 0.00028137999999999997 3.3 0.00028147999999999997 0 0.0002814 0 0.0002815 3.3 0.00028142 3.3 0.00028152 0 0.00028144 0 0.00028154 3.3 0.00028146 3.3 0.00028156 0 0.00028147999999999997 0 0.00028157999999999997 3.3 0.0002815 3.3 0.0002816 0 0.00028152 0 0.00028162 3.3 0.00028154 3.3 0.00028164 0 0.00028156 0 0.00028166 3.3 0.00028157999999999997 3.3 0.00028168 0 0.0002816 0 0.0002817 3.3 0.00028162 3.3 0.00028172 0 0.00028164 0 0.00028174 3.3 0.00028166 3.3 0.00028176 0 0.00028168 0 0.00028178 3.3 0.0002817 3.3 0.0002818 0 0.00028172 0 0.00028182 3.3 0.00028174 3.3 0.00028184 0 0.00028176 0 0.00028186 3.3 0.00028178 3.3 0.00028188 0 0.00028179999999999997 0 0.00028189999999999997 3.3 0.00028182 3.3 0.00028192 0 0.00028184 0 0.00028194 3.3 0.00028186 3.3 0.00028196 0 0.00028188 0 0.00028198 3.3 0.00028189999999999997 3.3 0.00028199999999999997 0 0.00028192 0 0.00028202 3.3 0.00028194 3.3 0.00028204 0 0.00028196 0 0.00028206 3.3 0.00028198 3.3 0.00028208 0 0.00028199999999999997 0 0.00028209999999999997 3.3 0.00028202 3.3 0.00028212 0 0.00028204 0 0.00028214 3.3 0.00028206 3.3 0.00028216 0 0.00028208 0 0.00028218 3.3 0.00028209999999999997 3.3 0.0002822 0 0.00028212 0 0.00028222 3.3 0.00028214 3.3 0.00028224 0 0.00028216 0 0.00028226 3.3 0.00028218 3.3 0.00028228 0 0.0002822 0 0.0002823 3.3 0.00028222 3.3 0.00028232 0 0.00028224 0 0.00028234 3.3 0.00028226 3.3 0.00028236 0 0.00028228 0 0.00028238 3.3 0.0002823 3.3 0.0002824 0 0.00028231999999999997 0 0.00028241999999999997 3.3 0.00028234 3.3 0.00028244 0 0.00028236 0 0.00028246 3.3 0.00028238 3.3 0.00028248 0 0.0002824 0 0.0002825 3.3 0.00028241999999999997 3.3 0.00028251999999999997 0 0.00028244 0 0.00028254 3.3 0.00028246 3.3 0.00028256 0 0.00028248 0 0.00028258 3.3 0.0002825 3.3 0.0002826 0 0.00028251999999999997 0 0.00028262 3.3 0.00028254 3.3 0.00028264 0 0.00028256 0 0.00028266 3.3 0.00028258 3.3 0.00028268 0 0.0002826 0 0.0002827 3.3 0.00028262 3.3 0.00028272 0 0.00028264 0 0.00028274 3.3 0.00028266 3.3 0.00028276 0 0.00028268 0 0.00028278 3.3 0.0002827 3.3 0.0002828 0 0.00028272 0 0.00028282 3.3 0.00028273999999999997 3.3 0.00028283999999999997 0 0.00028276 0 0.00028286 3.3 0.00028278 3.3 0.00028288 0 0.0002828 0 0.0002829 3.3 0.00028282 3.3 0.00028292 0 0.00028283999999999997 0 0.00028293999999999997 3.3 0.00028286 3.3 0.00028296 0 0.00028288 0 0.00028298 3.3 0.0002829 3.3 0.000283 0 0.00028292 0 0.00028302 3.3 0.00028293999999999997 3.3 0.00028304 0 0.00028296 0 0.00028306 3.3 0.00028298 3.3 0.00028308 0 0.000283 0 0.0002831 3.3 0.00028302 3.3 0.00028312 0 0.00028304 0 0.00028314 3.3 0.00028306 3.3 0.00028316 0 0.00028308 0 0.00028318 3.3 0.0002831 3.3 0.0002832 0 0.00028312 0 0.00028322 3.3 0.00028314 3.3 0.00028324 0 0.00028315999999999997 0 0.00028325999999999997 3.3 0.00028318 3.3 0.00028328 0 0.0002832 0 0.0002833 3.3 0.00028322 3.3 0.00028332 0 0.00028324 0 0.00028334 3.3 0.00028325999999999997 3.3 0.00028335999999999997 0 0.00028328 0 0.00028338 3.3 0.0002833 3.3 0.0002834 0 0.00028332 0 0.00028342 3.3 0.00028334 3.3 0.00028344 0 0.00028335999999999997 0 0.00028345999999999997 3.3 0.00028338 3.3 0.00028348 0 0.0002834 0 0.0002835 3.3 0.00028342 3.3 0.00028352 0 0.00028344 0 0.00028354 3.3 0.00028345999999999997 3.3 0.00028356 0 0.00028348 0 0.00028358 3.3 0.0002835 3.3 0.0002836 0 0.00028352 0 0.00028362 3.3 0.00028354 3.3 0.00028364 0 0.00028356 0 0.00028366 3.3 0.00028357999999999996 3.3 0.00028367999999999997 0 0.0002836 0 0.0002837 3.3 0.00028362 3.3 0.00028372 0 0.00028364 0 0.00028374 3.3 0.00028366 3.3 0.00028376 0 0.00028367999999999997 0 0.00028377999999999997 3.3 0.0002837 3.3 0.0002838 0 0.00028372 0 0.00028382 3.3 0.00028374 3.3 0.00028384 0 0.00028376 0 0.00028386 3.3 0.00028377999999999997 3.3 0.00028387999999999997 0 0.0002838 0 0.0002839 3.3 0.00028382 3.3 0.00028392 0 0.00028384 0 0.00028394 3.3 0.00028386 3.3 0.00028396 0 0.00028387999999999997 0 0.00028398 3.3 0.0002839 3.3 0.000284 0 0.00028392 0 0.00028402 3.3 0.00028394 3.3 0.00028404 0 0.00028396 0 0.00028406 3.3 0.00028398 3.3 0.00028408 0 0.000284 0 0.0002841 3.3 0.00028402 3.3 0.00028412 0 0.00028404 0 0.00028414 3.3 0.00028406 3.3 0.00028416 0 0.00028408 0 0.00028418 3.3 0.00028409999999999997 3.3 0.00028419999999999997 0 0.00028412 0 0.00028422 3.3 0.00028414 3.3 0.00028424 0 0.00028416 0 0.00028426 3.3 0.00028418 3.3 0.00028428 0 0.00028419999999999997 0 0.00028429999999999997 3.3 0.00028422 3.3 0.00028432 0 0.00028424 0 0.00028434 3.3 0.00028426 3.3 0.00028436 0 0.00028428 0 0.00028438 3.3 0.00028429999999999997 3.3 0.0002844 0 0.00028432 0 0.00028442 3.3 0.00028434 3.3 0.00028444 0 0.00028436 0 0.00028446 3.3 0.00028438 3.3 0.00028448 0 0.0002844 0 0.0002845 3.3 0.00028442 3.3 0.00028452 0 0.00028444 0 0.00028454 3.3 0.00028446 3.3 0.00028456 0 0.00028448 0 0.00028458 3.3 0.0002845 3.3 0.0002846 0 0.00028451999999999997 0 0.00028461999999999997 3.3 0.00028454 3.3 0.00028464 0 0.00028456 0 0.00028466 3.3 0.00028458 3.3 0.00028468 0 0.0002846 0 0.0002847 3.3 0.00028461999999999997 3.3 0.00028471999999999997 0 0.00028464 0 0.00028474 3.3 0.00028466 3.3 0.00028476 0 0.00028468 0 0.00028478 3.3 0.0002847 3.3 0.0002848 0 0.00028471999999999997 0 0.00028482 3.3 0.00028474 3.3 0.00028484 0 0.00028476 0 0.00028486 3.3 0.00028478 3.3 0.00028488 0 0.0002848 0 0.0002849 3.3 0.00028482 3.3 0.00028492 0 0.00028484 0 0.00028494 3.3 0.00028486 3.3 0.00028496 0 0.00028488 0 0.00028498 3.3 0.0002849 3.3 0.000285 0 0.00028492 0 0.00028502 3.3 0.00028493999999999997 3.3 0.00028503999999999997 0 0.00028496 0 0.00028506 3.3 0.00028498 3.3 0.00028508 0 0.000285 0 0.0002851 3.3 0.00028502 3.3 0.00028512 0 0.00028503999999999997 0 0.00028513999999999997 3.3 0.00028506 3.3 0.00028516 0 0.00028508 0 0.00028518 3.3 0.0002851 3.3 0.0002852 0 0.00028512 0 0.00028522 3.3 0.00028513999999999997 3.3 0.00028523999999999997 0 0.00028516 0 0.00028526 3.3 0.00028518 3.3 0.00028528 0 0.0002852 0 0.0002853 3.3 0.00028522 3.3 0.00028532 0 0.00028523999999999997 0 0.00028534 3.3 0.00028526 3.3 0.00028536 0 0.00028528 0 0.00028538 3.3 0.0002853 3.3 0.0002854 0 0.00028532 0 0.00028542 3.3 0.00028534 3.3 0.00028544 0 0.00028535999999999996 0 0.00028545999999999997 3.3 0.00028538 3.3 0.00028548 0 0.0002854 0 0.0002855 3.3 0.00028542 3.3 0.00028552 0 0.00028544 0 0.00028554 3.3 0.00028545999999999997 3.3 0.00028555999999999997 0 0.00028548 0 0.00028558 3.3 0.0002855 3.3 0.0002856 0 0.00028552 0 0.00028562 3.3 0.00028554 3.3 0.00028564 0 0.00028555999999999997 0 0.00028565999999999997 3.3 0.00028558 3.3 0.00028568 0 0.0002856 0 0.0002857 3.3 0.00028562 3.3 0.00028572 0 0.00028564 0 0.00028574 3.3 0.00028565999999999997 3.3 0.00028576 0 0.00028568 0 0.00028578 3.3 0.0002857 3.3 0.0002858 0 0.00028572 0 0.00028582 3.3 0.00028574 3.3 0.00028584 0 0.00028576 0 0.00028586 3.3 0.00028578 3.3 0.00028588 0 0.0002858 0 0.0002859 3.3 0.00028582 3.3 0.00028592 0 0.00028584 0 0.00028594 3.3 0.00028586 3.3 0.00028596 0 0.00028587999999999997 0 0.00028597999999999997 3.3 0.0002859 3.3 0.000286 0 0.00028592 0 0.00028602 3.3 0.00028594 3.3 0.00028604 0 0.00028596 0 0.00028606 3.3 0.00028597999999999997 3.3 0.00028607999999999997 0 0.000286 0 0.0002861 3.3 0.00028602 3.3 0.00028612 0 0.00028604 0 0.00028614 3.3 0.00028606 3.3 0.00028616 0 0.00028607999999999997 0 0.00028618 3.3 0.0002861 3.3 0.0002862 0 0.00028612 0 0.00028622 3.3 0.00028614 3.3 0.00028624 0 0.00028616 0 0.00028626 3.3 0.00028618 3.3 0.00028628 0 0.0002862 0 0.0002863 3.3 0.00028622 3.3 0.00028632 0 0.00028624 0 0.00028634 3.3 0.00028626 3.3 0.00028636 0 0.00028628 0 0.00028638 3.3 0.00028629999999999997 3.3 0.00028639999999999997 0 0.00028632 0 0.00028642 3.3 0.00028634 3.3 0.00028644 0 0.00028636 0 0.00028646 3.3 0.00028638 3.3 0.00028648 0 0.00028639999999999997 0 0.00028649999999999997 3.3 0.00028642 3.3 0.00028652 0 0.00028644 0 0.00028654 3.3 0.00028646 3.3 0.00028656 0 0.00028648 0 0.00028658 3.3 0.00028649999999999997 3.3 0.0002866 0 0.00028652 0 0.00028662 3.3 0.00028654 3.3 0.00028664 0 0.00028656 0 0.00028666 3.3 0.00028658 3.3 0.00028668 0 0.0002866 0 0.0002867 3.3 0.00028662 3.3 0.00028672 0 0.00028664 0 0.00028674 3.3 0.00028666 3.3 0.00028676 0 0.00028668 0 0.00028678 3.3 0.0002867 3.3 0.0002868 0 0.00028671999999999997 0 0.00028681999999999997 3.3 0.00028674 3.3 0.00028684 0 0.00028676 0 0.00028686 3.3 0.00028678 3.3 0.00028688 0 0.0002868 0 0.0002869 3.3 0.00028681999999999997 3.3 0.00028691999999999997 0 0.00028684 0 0.00028694 3.3 0.00028686 3.3 0.00028696 0 0.00028688 0 0.00028698 3.3 0.0002869 3.3 0.000287 0 0.00028691999999999997 0 0.00028701999999999997 3.3 0.00028694 3.3 0.00028704 0 0.00028696 0 0.00028706 3.3 0.00028698 3.3 0.00028708 0 0.000287 0 0.0002871 3.3 0.00028701999999999997 3.3 0.00028712 0 0.00028704 0 0.00028714 3.3 0.00028706 3.3 0.00028716 0 0.00028708 0 0.00028718 3.3 0.0002871 3.3 0.0002872 0 0.00028712 0 0.00028722 3.3 0.00028713999999999996 3.3 0.00028723999999999997 0 0.00028716 0 0.00028726 3.3 0.00028718 3.3 0.00028728 0 0.0002872 0 0.0002873 3.3 0.00028722 3.3 0.00028732 0 0.00028723999999999997 0 0.00028733999999999997 3.3 0.00028726 3.3 0.00028736 0 0.00028728 0 0.00028738 3.3 0.0002873 3.3 0.0002874 0 0.00028732 0 0.00028742 3.3 0.00028733999999999997 3.3 0.00028743999999999997 0 0.00028736 0 0.00028746 3.3 0.00028738 3.3 0.00028748 0 0.0002874 0 0.0002875 3.3 0.00028742 3.3 0.00028752 0 0.00028743999999999997 0 0.00028754 3.3 0.00028746 3.3 0.00028756 0 0.00028748 0 0.00028758 3.3 0.0002875 3.3 0.0002876 0 0.00028752 0 0.00028762 3.3 0.00028754 3.3 0.00028764 0 0.00028756 0 0.00028766 3.3 0.00028758 3.3 0.00028768 0 0.0002876 0 0.0002877 3.3 0.00028762 3.3 0.00028772 0 0.00028764 0 0.00028774 3.3 0.00028765999999999997 3.3 0.00028775999999999997 0 0.00028768 0 0.00028778 3.3 0.0002877 3.3 0.0002878 0 0.00028772 0 0.00028782 3.3 0.00028774 3.3 0.00028784 0 0.00028775999999999997 0 0.00028785999999999997 3.3 0.00028778 3.3 0.00028788 0 0.0002878 0 0.0002879 3.3 0.00028782 3.3 0.00028792 0 0.00028784 0 0.00028794 3.3 0.00028785999999999997 3.3 0.00028796 0 0.00028788 0 0.00028798 3.3 0.0002879 3.3 0.000288 0 0.00028792 0 0.00028802 3.3 0.00028794 3.3 0.00028804 0 0.00028796 0 0.00028806 3.3 0.00028798 3.3 0.00028808 0 0.000288 0 0.0002881 3.3 0.00028802 3.3 0.00028812 0 0.00028804 0 0.00028814 3.3 0.00028806 3.3 0.00028816 0 0.00028807999999999997 0 0.00028817999999999997 3.3 0.0002881 3.3 0.0002882 0 0.00028812 0 0.00028822 3.3 0.00028814 3.3 0.00028824 0 0.00028816 0 0.00028826 3.3 0.00028817999999999997 3.3 0.00028827999999999997 0 0.0002882 0 0.0002883 3.3 0.00028822 3.3 0.00028832 0 0.00028824 0 0.00028834 3.3 0.00028826 3.3 0.00028836 0 0.00028827999999999997 0 0.00028838 3.3 0.0002883 3.3 0.0002884 0 0.00028832 0 0.00028842 3.3 0.00028834 3.3 0.00028844 0 0.00028836 0 0.00028846 3.3 0.00028838 3.3 0.00028848 0 0.0002884 0 0.0002885 3.3 0.00028842 3.3 0.00028852 0 0.00028844 0 0.00028854 3.3 0.00028846 3.3 0.00028856 0 0.00028848 0 0.00028858 3.3 0.00028849999999999997 3.3 0.00028859999999999997 0 0.00028852 0 0.00028862 3.3 0.00028854 3.3 0.00028864 0 0.00028856 0 0.00028866 3.3 0.00028858 3.3 0.00028868 0 0.00028859999999999997 0 0.00028869999999999997 3.3 0.00028862 3.3 0.00028872 0 0.00028864 0 0.00028874 3.3 0.00028866 3.3 0.00028876 0 0.00028868 0 0.00028878 3.3 0.00028869999999999997 3.3 0.00028879999999999997 0 0.00028872 0 0.00028882 3.3 0.00028874 3.3 0.00028884 0 0.00028876 0 0.00028886 3.3 0.00028878 3.3 0.00028888 0 0.00028879999999999997 0 0.0002889 3.3 0.00028882 3.3 0.00028892 0 0.00028884 0 0.00028894 3.3 0.00028886 3.3 0.00028896 0 0.00028888 0 0.00028898 3.3 0.0002889 3.3 0.000289 0 0.00028892 0 0.00028902 3.3 0.00028894 3.3 0.00028904 0 0.00028896 0 0.00028906 3.3 0.00028898 3.3 0.00028908 0 0.000289 0 0.0002891 3.3 0.00028901999999999997 3.3 0.00028911999999999997 0 0.00028904 0 0.00028914 3.3 0.00028906 3.3 0.00028916 0 0.00028908 0 0.00028918 3.3 0.0002891 3.3 0.0002892 0 0.00028911999999999997 0 0.00028921999999999997 3.3 0.00028914 3.3 0.00028924 0 0.00028916 0 0.00028926 3.3 0.00028918 3.3 0.00028928 0 0.0002892 0 0.0002893 3.3 0.00028921999999999997 3.3 0.00028932 0 0.00028924 0 0.00028934 3.3 0.00028926 3.3 0.00028936 0 0.00028928 0 0.00028938 3.3 0.0002893 3.3 0.0002894 0 0.00028932 0 0.00028942 3.3 0.00028934 3.3 0.00028944 0 0.00028936 0 0.00028946 3.3 0.00028938 3.3 0.00028948 0 0.0002894 0 0.0002895 3.3 0.00028942 3.3 0.00028952 0 0.00028943999999999997 0 0.00028953999999999997 3.3 0.00028946 3.3 0.00028956 0 0.00028948 0 0.00028958 3.3 0.0002895 3.3 0.0002896 0 0.00028952 0 0.00028962 3.3 0.00028953999999999997 3.3 0.00028963999999999997 0 0.00028956 0 0.00028966 3.3 0.00028958 3.3 0.00028968 0 0.0002896 0 0.0002897 3.3 0.00028962 3.3 0.00028972 0 0.00028963999999999997 0 0.00028974 3.3 0.00028966 3.3 0.00028976 0 0.00028968 0 0.00028978 3.3 0.0002897 3.3 0.0002898 0 0.00028972 0 0.00028982 3.3 0.00028974 3.3 0.00028984 0 0.00028976 0 0.00028986 3.3 0.00028978 3.3 0.00028988 0 0.0002898 0 0.0002899 3.3 0.00028982 3.3 0.00028992 0 0.00028984 0 0.00028994 3.3 0.00028985999999999997 3.3 0.00028995999999999997 0 0.00028988 0 0.00028998 3.3 0.0002899 3.3 0.00029 0 0.00028992 0 0.00029002 3.3 0.00028994 3.3 0.00029004 0 0.00028995999999999997 0 0.00029005999999999997 3.3 0.00028998 3.3 0.00029008 0 0.00029 0 0.0002901 3.3 0.00029002 3.3 0.00029012 0 0.00029004 0 0.00029014 3.3 0.00029005999999999997 3.3 0.00029016 0 0.00029008 0 0.00029018 3.3 0.0002901 3.3 0.0002902 0 0.00029012 0 0.00029022 3.3 0.00029014 3.3 0.00029024 0 0.00029016 0 0.00029026 3.3 0.00029018 3.3 0.00029028 0 0.0002902 0 0.0002903 3.3 0.00029022 3.3 0.00029032 0 0.00029024 0 0.00029034 3.3 0.00029026 3.3 0.00029036 0 0.00029027999999999997 0 0.00029037999999999997 3.3 0.0002903 3.3 0.0002904 0 0.00029032 0 0.00029042 3.3 0.00029034 3.3 0.00029044 0 0.00029036 0 0.00029046 3.3 0.00029037999999999997 3.3 0.00029047999999999997 0 0.0002904 0 0.0002905 3.3 0.00029042 3.3 0.00029052 0 0.00029044 0 0.00029054 3.3 0.00029046 3.3 0.00029056 0 0.00029047999999999997 0 0.00029057999999999997 3.3 0.0002905 3.3 0.0002906 0 0.00029052 0 0.00029062 3.3 0.00029054 3.3 0.00029064 0 0.00029056 0 0.00029066 3.3 0.00029057999999999997 3.3 0.00029068 0 0.0002906 0 0.0002907 3.3 0.00029062 3.3 0.00029072 0 0.00029064 0 0.00029074 3.3 0.00029066 3.3 0.00029076 0 0.00029068 0 0.00029078 3.3 0.0002907 3.3 0.0002908 0 0.00029072 0 0.00029082 3.3 0.00029074 3.3 0.00029084 0 0.00029076 0 0.00029086 3.3 0.00029078 3.3 0.00029088 0 0.00029079999999999997 0 0.00029089999999999997 3.3 0.00029082 3.3 0.00029092 0 0.00029084 0 0.00029094 3.3 0.00029086 3.3 0.00029096 0 0.00029088 0 0.00029098 3.3 0.00029089999999999997 3.3 0.00029099999999999997 0 0.00029092 0 0.00029102 3.3 0.00029094 3.3 0.00029104 0 0.00029096 0 0.00029106 3.3 0.00029098 3.3 0.00029108 0 0.00029099999999999997 0 0.0002911 3.3 0.00029102 3.3 0.00029112 0 0.00029104 0 0.00029114 3.3 0.00029106 3.3 0.00029116 0 0.00029108 0 0.00029118 3.3 0.0002911 3.3 0.0002912 0 0.00029112 0 0.00029122 3.3 0.00029114 3.3 0.00029124 0 0.00029116 0 0.00029126 3.3 0.00029118 3.3 0.00029128 0 0.0002912 0 0.0002913 3.3 0.00029121999999999997 3.3 0.00029131999999999997 0 0.00029124 0 0.00029134 3.3 0.00029126 3.3 0.00029136 0 0.00029128 0 0.00029138 3.3 0.0002913 3.3 0.0002914 0 0.00029131999999999997 0 0.00029141999999999997 3.3 0.00029134 3.3 0.00029144 0 0.00029136 0 0.00029146 3.3 0.00029138 3.3 0.00029148 0 0.0002914 0 0.0002915 3.3 0.00029141999999999997 3.3 0.00029152 0 0.00029144 0 0.00029154 3.3 0.00029146 3.3 0.00029156 0 0.00029148 0 0.00029158 3.3 0.0002915 3.3 0.0002916 0 0.00029152 0 0.00029162 3.3 0.00029154 3.3 0.00029164 0 0.00029156 0 0.00029166 3.3 0.00029158 3.3 0.00029168 0 0.0002916 0 0.0002917 3.3 0.00029162 3.3 0.00029172 0 0.00029163999999999997 0 0.00029173999999999997 3.3 0.00029166 3.3 0.00029176 0 0.00029168 0 0.00029178 3.3 0.0002917 3.3 0.0002918 0 0.00029172 0 0.00029182 3.3 0.00029173999999999997 3.3 0.00029183999999999997 0 0.00029176 0 0.00029186 3.3 0.00029178 3.3 0.00029188 0 0.0002918 0 0.0002919 3.3 0.00029182 3.3 0.00029192 0 0.00029183999999999997 0 0.00029194 3.3 0.00029186 3.3 0.00029196 0 0.00029188 0 0.00029198 3.3 0.0002919 3.3 0.000292 0 0.00029192 0 0.00029202 3.3 0.00029194 3.3 0.00029204 0 0.00029196 0 0.00029206 3.3 0.00029198 3.3 0.00029208 0 0.000292 0 0.0002921 3.3 0.00029202 3.3 0.00029212 0 0.00029204 0 0.00029214 3.3 0.00029205999999999997 3.3 0.00029215999999999997 0 0.00029208 0 0.00029218 3.3 0.0002921 3.3 0.0002922 0 0.00029212 0 0.00029222 3.3 0.00029214 3.3 0.00029224 0 0.00029215999999999997 0 0.00029225999999999997 3.3 0.00029218 3.3 0.00029228 0 0.0002922 0 0.0002923 3.3 0.00029222 3.3 0.00029232 0 0.00029224 0 0.00029234 3.3 0.00029225999999999997 3.3 0.00029235999999999997 0 0.00029228 0 0.00029238 3.3 0.0002923 3.3 0.0002924 0 0.00029232 0 0.00029242 3.3 0.00029234 3.3 0.00029244 0 0.00029235999999999997 0 0.00029246 3.3 0.00029238 3.3 0.00029248 0 0.0002924 0 0.0002925 3.3 0.00029242 3.3 0.00029252 0 0.00029244 0 0.00029254 3.3 0.00029246 3.3 0.00029256 0 0.00029248 0 0.00029258 3.3 0.0002925 3.3 0.0002926 0 0.00029252 0 0.00029262 3.3 0.00029254 3.3 0.00029264 0 0.00029256 0 0.00029266 3.3 0.00029257999999999997 3.3 0.00029267999999999997 0 0.0002926 0 0.0002927 3.3 0.00029262 3.3 0.00029272 0 0.00029264 0 0.00029274 3.3 0.00029266 3.3 0.00029276 0 0.00029267999999999997 0 0.00029277999999999997 3.3 0.0002927 3.3 0.0002928 0 0.00029272 0 0.00029282 3.3 0.00029274 3.3 0.00029284 0 0.00029276 0 0.00029286 3.3 0.00029277999999999997 3.3 0.00029288 0 0.0002928 0 0.0002929 3.3 0.00029282 3.3 0.00029292 0 0.00029284 0 0.00029294 3.3 0.00029286 3.3 0.00029296 0 0.00029288 0 0.00029298 3.3 0.0002929 3.3 0.000293 0 0.00029292 0 0.00029302 3.3 0.00029294 3.3 0.00029304 0 0.00029296 0 0.00029306 3.3 0.00029298 3.3 0.00029308 0 0.00029299999999999997 0 0.00029309999999999997 3.3 0.00029302 3.3 0.00029312 0 0.00029304 0 0.00029314 3.3 0.00029306 3.3 0.00029316 0 0.00029308 0 0.00029318 3.3 0.00029309999999999997 3.3 0.00029319999999999997 0 0.00029312 0 0.00029322 3.3 0.00029314 3.3 0.00029324 0 0.00029316 0 0.00029326 3.3 0.00029318 3.3 0.00029328 0 0.00029319999999999997 0 0.0002933 3.3 0.00029322 3.3 0.00029332 0 0.00029324 0 0.00029334 3.3 0.00029326 3.3 0.00029336 0 0.00029328 0 0.00029338 3.3 0.0002933 3.3 0.0002934 0 0.00029332 0 0.00029342 3.3 0.00029334 3.3 0.00029344 0 0.00029336 0 0.00029346 3.3 0.00029338 3.3 0.00029348 0 0.0002934 0 0.0002935 3.3 0.00029341999999999997 3.3 0.00029351999999999997 0 0.00029344 0 0.00029354 3.3 0.00029346 3.3 0.00029356 0 0.00029348 0 0.00029358 3.3 0.0002935 3.3 0.0002936 0 0.00029351999999999997 0 0.00029361999999999997 3.3 0.00029354 3.3 0.00029364 0 0.00029356 0 0.00029366 3.3 0.00029358 3.3 0.00029368 0 0.0002936 0 0.0002937 3.3 0.00029361999999999997 3.3 0.00029371999999999997 0 0.00029364 0 0.00029374 3.3 0.00029366 3.3 0.00029376 0 0.00029368 0 0.00029378 3.3 0.0002937 3.3 0.0002938 0 0.00029371999999999997 0 0.00029382 3.3 0.00029374 3.3 0.00029384 0 0.00029376 0 0.00029386 3.3 0.00029378 3.3 0.00029388 0 0.0002938 0 0.0002939 3.3 0.00029382 3.3 0.00029392 0 0.00029383999999999996 0 0.00029393999999999997 3.3 0.00029386 3.3 0.00029396 0 0.00029388 0 0.00029398 3.3 0.0002939 3.3 0.000294 0 0.00029392 0 0.00029402 3.3 0.00029393999999999997 3.3 0.00029403999999999997 0 0.00029396 0 0.00029406 3.3 0.00029398 3.3 0.00029408 0 0.000294 0 0.0002941 3.3 0.00029402 3.3 0.00029412 0 0.00029403999999999997 0 0.00029413999999999997 3.3 0.00029406 3.3 0.00029416 0 0.00029408 0 0.00029418 3.3 0.0002941 3.3 0.0002942 0 0.00029412 0 0.00029422 3.3 0.00029413999999999997 3.3 0.00029424 0 0.00029416 0 0.00029426 3.3 0.00029418 3.3 0.00029428 0 0.0002942 0 0.0002943 3.3 0.00029422 3.3 0.00029432 0 0.00029424 0 0.00029434 3.3 0.00029426 3.3 0.00029436 0 0.00029428 0 0.00029438 3.3 0.0002943 3.3 0.0002944 0 0.00029432 0 0.00029442 3.3 0.00029434 3.3 0.00029444 0 0.00029435999999999997 0 0.00029445999999999997 3.3 0.00029438 3.3 0.00029448 0 0.0002944 0 0.0002945 3.3 0.00029442 3.3 0.00029452 0 0.00029444 0 0.00029454 3.3 0.00029445999999999997 3.3 0.00029455999999999997 0 0.00029448 0 0.00029458 3.3 0.0002945 3.3 0.0002946 0 0.00029452 0 0.00029462 3.3 0.00029454 3.3 0.00029464 0 0.00029455999999999997 0 0.00029466 3.3 0.00029458 3.3 0.00029468 0 0.0002946 0 0.0002947 3.3 0.00029462 3.3 0.00029472 0 0.00029464 0 0.00029474 3.3 0.00029466 3.3 0.00029476 0 0.00029468 0 0.00029478 3.3 0.0002947 3.3 0.0002948 0 0.00029472 0 0.00029482 3.3 0.00029474 3.3 0.00029484 0 0.00029476 0 0.00029486 3.3 0.00029477999999999997 3.3 0.00029487999999999997 0 0.0002948 0 0.0002949 3.3 0.00029482 3.3 0.00029492 0 0.00029484 0 0.00029494 3.3 0.00029486 3.3 0.00029496 0 0.00029487999999999997 0 0.00029497999999999997 3.3 0.0002949 3.3 0.000295 0 0.00029492 0 0.00029502 3.3 0.00029494 3.3 0.00029504 0 0.00029496 0 0.00029506 3.3 0.00029497999999999997 3.3 0.00029508 0 0.000295 0 0.0002951 3.3 0.00029502 3.3 0.00029512 0 0.00029504 0 0.00029514 3.3 0.00029506 3.3 0.00029516 0 0.00029508 0 0.00029518 3.3 0.0002951 3.3 0.0002952 0 0.00029512 0 0.00029522 3.3 0.00029514 3.3 0.00029524 0 0.00029516 0 0.00029526 3.3 0.00029518 3.3 0.00029528 0 0.00029519999999999997 0 0.00029529999999999997 3.3 0.00029522 3.3 0.00029532 0 0.00029524 0 0.00029534 3.3 0.00029526 3.3 0.00029536 0 0.00029528 0 0.00029538 3.3 0.00029529999999999997 3.3 0.00029539999999999997 0 0.00029532 0 0.00029542 3.3 0.00029534 3.3 0.00029544 0 0.00029536 0 0.00029546 3.3 0.00029538 3.3 0.00029548 0 0.00029539999999999997 0 0.00029549999999999997 3.3 0.00029542 3.3 0.00029552 0 0.00029544 0 0.00029554 3.3 0.00029546 3.3 0.00029556 0 0.00029548 0 0.00029558 3.3 0.00029549999999999997 3.3 0.0002956 0 0.00029552 0 0.00029562 3.3 0.00029554 3.3 0.00029564 0 0.00029556 0 0.00029566 3.3 0.00029558 3.3 0.00029568 0 0.0002956 0 0.0002957 3.3 0.00029561999999999996 3.3 0.00029571999999999997 0 0.00029564 0 0.00029574 3.3 0.00029566 3.3 0.00029576 0 0.00029568 0 0.00029578 3.3 0.0002957 3.3 0.0002958 0 0.00029571999999999997 0 0.00029581999999999997 3.3 0.00029574 3.3 0.00029584 0 0.00029576 0 0.00029586 3.3 0.00029578 3.3 0.00029588 0 0.0002958 0 0.0002959 3.3 0.00029581999999999997 3.3 0.00029591999999999997 0 0.00029584 0 0.00029594 3.3 0.00029586 3.3 0.00029596 0 0.00029588 0 0.00029598 3.3 0.0002959 3.3 0.000296 0 0.00029591999999999997 0 0.00029602 3.3 0.00029594 3.3 0.00029604 0 0.00029596 0 0.00029606 3.3 0.00029598 3.3 0.00029608 0 0.000296 0 0.0002961 3.3 0.00029602 3.3 0.00029612 0 0.00029604 0 0.00029614 3.3 0.00029606 3.3 0.00029616 0 0.00029608 0 0.00029618 3.3 0.0002961 3.3 0.0002962 0 0.00029612 0 0.00029622 3.3 0.00029613999999999997 3.3 0.00029623999999999997 0 0.00029616 0 0.00029626 3.3 0.00029618 3.3 0.00029628 0 0.0002962 0 0.0002963 3.3 0.00029622 3.3 0.00029632 0 0.00029623999999999997 0 0.00029633999999999997 3.3 0.00029626 3.3 0.00029636 0 0.00029628 0 0.00029638 3.3 0.0002963 3.3 0.0002964 0 0.00029632 0 0.00029642 3.3 0.00029633999999999997 3.3 0.00029644 0 0.00029636 0 0.00029646 3.3 0.00029638 3.3 0.00029648 0 0.0002964 0 0.0002965 3.3 0.00029642 3.3 0.00029652 0 0.00029644 0 0.00029654 3.3 0.00029646 3.3 0.00029656 0 0.00029648 0 0.00029658 3.3 0.0002965 3.3 0.0002966 0 0.00029652 0 0.00029662 3.3 0.00029654 3.3 0.00029664 0 0.00029655999999999997 0 0.00029665999999999997 3.3 0.00029658 3.3 0.00029668 0 0.0002966 0 0.0002967 3.3 0.00029662 3.3 0.00029672 0 0.00029664 0 0.00029674 3.3 0.00029665999999999997 3.3 0.00029675999999999997 0 0.00029668 0 0.00029678 3.3 0.0002967 3.3 0.0002968 0 0.00029672 0 0.00029682 3.3 0.00029674 3.3 0.00029684 0 0.00029675999999999997 0 0.00029686 3.3 0.00029678 3.3 0.00029688 0 0.0002968 0 0.0002969 3.3 0.00029682 3.3 0.00029692 0 0.00029684 0 0.00029694 3.3 0.00029686 3.3 0.00029696 0 0.00029688 0 0.00029698 3.3 0.0002969 3.3 0.000297 0 0.00029692 0 0.00029702 3.3 0.00029694 3.3 0.00029704 0 0.00029696 0 0.00029706 3.3 0.00029697999999999997 3.3 0.00029707999999999997 0 0.000297 0 0.0002971 3.3 0.00029702 3.3 0.00029712 0 0.00029704 0 0.00029714 3.3 0.00029706 3.3 0.00029716 0 0.00029707999999999997 0 0.00029717999999999997 3.3 0.0002971 3.3 0.0002972 0 0.00029712 0 0.00029722 3.3 0.00029714 3.3 0.00029724 0 0.00029716 0 0.00029726 3.3 0.00029717999999999997 3.3 0.00029727999999999997 0 0.0002972 0 0.0002973 3.3 0.00029722 3.3 0.00029732 0 0.00029724 0 0.00029734 3.3 0.00029726 3.3 0.00029736 0 0.00029727999999999997 0 0.00029738 3.3 0.0002973 3.3 0.0002974 0 0.00029732 0 0.00029742 3.3 0.00029734 3.3 0.00029744 0 0.00029736 0 0.00029746 3.3 0.00029738 3.3 0.00029748 0 0.00029739999999999996 0 0.00029749999999999997 3.3 0.00029742 3.3 0.00029752 0 0.00029744 0 0.00029754 3.3 0.00029746 3.3 0.00029756 0 0.00029748 0 0.00029758 3.3 0.00029749999999999997 3.3 0.00029759999999999997 0 0.00029752 0 0.00029762 3.3 0.00029754 3.3 0.00029764 0 0.00029756 0 0.00029766 3.3 0.00029758 3.3 0.00029768 0 0.00029759999999999997 0 0.00029769999999999997 3.3 0.00029762 3.3 0.00029772 0 0.00029764 0 0.00029774 3.3 0.00029766 3.3 0.00029776 0 0.00029768 0 0.00029778 3.3 0.00029769999999999997 3.3 0.0002978 0 0.00029772 0 0.00029782 3.3 0.00029774 3.3 0.00029784 0 0.00029776 0 0.00029786 3.3 0.00029778 3.3 0.00029788 0 0.0002978 0 0.0002979 3.3 0.00029782 3.3 0.00029792 0 0.00029784 0 0.00029794 3.3 0.00029786 3.3 0.00029796 0 0.00029788 0 0.00029798 3.3 0.0002979 3.3 0.000298 0 0.00029791999999999997 0 0.00029801999999999997 3.3 0.00029794 3.3 0.00029804 0 0.00029796 0 0.00029806 3.3 0.00029798 3.3 0.00029808 0 0.000298 0 0.0002981 3.3 0.00029801999999999997 3.3 0.00029811999999999997 0 0.00029804 0 0.00029814 3.3 0.00029806 3.3 0.00029816 0 0.00029808 0 0.00029818 3.3 0.0002981 3.3 0.0002982 0 0.00029811999999999997 0 0.00029822 3.3 0.00029814 3.3 0.00029824 0 0.00029816 0 0.00029826 3.3 0.00029818 3.3 0.00029828 0 0.0002982 0 0.0002983 3.3 0.00029822 3.3 0.00029832 0 0.00029824 0 0.00029834 3.3 0.00029826 3.3 0.00029836 0 0.00029828 0 0.00029838 3.3 0.0002983 3.3 0.0002984 0 0.00029832 0 0.00029842 3.3 0.00029833999999999997 3.3 0.00029843999999999997 0 0.00029836 0 0.00029846 3.3 0.00029838 3.3 0.00029848 0 0.0002984 0 0.0002985 3.3 0.00029842 3.3 0.00029852 0 0.00029843999999999997 0 0.00029853999999999997 3.3 0.00029846 3.3 0.00029856 0 0.00029848 0 0.00029858 3.3 0.0002985 3.3 0.0002986 0 0.00029852 0 0.00029862 3.3 0.00029853999999999997 3.3 0.00029864 0 0.00029856 0 0.00029866 3.3 0.00029858 3.3 0.00029868 0 0.0002986 0 0.0002987 3.3 0.00029862 3.3 0.00029872 0 0.00029864 0 0.00029874 3.3 0.00029866 3.3 0.00029876 0 0.00029868 0 0.00029878 3.3 0.0002987 3.3 0.0002988 0 0.00029872 0 0.00029882 3.3 0.00029874 3.3 0.00029884 0 0.00029875999999999997 0 0.00029885999999999997 3.3 0.00029878 3.3 0.00029888 0 0.0002988 0 0.0002989 3.3 0.00029882 3.3 0.00029892 0 0.00029884 0 0.00029894 3.3 0.00029885999999999997 3.3 0.00029895999999999997 0 0.00029888 0 0.00029898 3.3 0.0002989 3.3 0.000299 0 0.00029892 0 0.00029902 3.3 0.00029894 3.3 0.00029904 0 0.00029895999999999997 0 0.00029905999999999997 3.3 0.00029898 3.3 0.00029908 0 0.000299 0 0.0002991 3.3 0.00029902 3.3 0.00029912 0 0.00029904 0 0.00029914 3.3 0.00029905999999999997 3.3 0.00029916 0 0.00029908 0 0.00029918 3.3 0.0002991 3.3 0.0002992 0 0.00029912 0 0.00029922 3.3 0.00029914 3.3 0.00029924 0 0.00029916 0 0.00029926 3.3 0.00029917999999999996 3.3 0.00029927999999999997 0 0.0002992 0 0.0002993 3.3 0.00029922 3.3 0.00029932 0 0.00029924 0 0.00029934 3.3 0.00029926 3.3 0.00029936 0 0.00029927999999999997 0 0.00029937999999999997 3.3 0.0002993 3.3 0.0002994 0 0.00029932 0 0.00029942 3.3 0.00029934 3.3 0.00029944 0 0.00029936 0 0.00029946 3.3 0.00029937999999999997 3.3 0.00029947999999999997 0 0.0002994 0 0.0002995 3.3 0.00029942 3.3 0.00029952 0 0.00029944 0 0.00029954 3.3 0.00029946 3.3 0.00029956 0 0.00029947999999999997 0 0.00029958 3.3 0.0002995 3.3 0.0002996 0 0.00029952 0 0.00029962 3.3 0.00029954 3.3 0.00029964 0 0.00029956 0 0.00029966 3.3 0.00029958 3.3 0.00029968 0 0.0002996 0 0.0002997 3.3 0.00029962 3.3 0.00029972 0 0.00029964 0 0.00029974 3.3 0.00029966 3.3 0.00029976 0 0.00029968 0 0.00029978 3.3 0.00029969999999999997 3.3 0.00029979999999999997 0 0.00029972 0 0.00029982 3.3 0.00029974 3.3 0.00029984 0 0.00029976 0 0.00029986 3.3 0.00029978 3.3 0.00029988 0 0.00029979999999999997 0 0.00029989999999999997 3.3 0.00029982 3.3 0.00029992 0 0.00029984 0 0.00029994 3.3 0.00029986 3.3 0.00029996 0 0.00029988 0 0.00029998 3.3 0.00029989999999999997 3.3 0.0003 0 0.00029992 0 0.00030002 3.3 0.00029994 3.3 0.00030004 0 0.00029996 0 0.00030006 3.3 0.00029998 3.3 0.00030008 0 0.0003 0 0.0003001 3.3 0.00030002 3.3 0.00030012 0 0.00030004 0 0.00030014 3.3 0.00030006 3.3 0.00030016 0 0.00030008 0 0.00030018 3.3 0.0003001 3.3 0.0003002 0 0.00030011999999999997 0 0.00030021999999999997 3.3 0.00030014 3.3 0.00030024 0 0.00030016 0 0.00030026 3.3 0.00030018 3.3 0.00030028 0 0.0003002 0 0.0003003 3.3 0.00030021999999999997 3.3 0.00030031999999999997 0 0.00030024 0 0.00030034 3.3 0.00030026 3.3 0.00030036 0 0.00030028 0 0.00030038 3.3 0.0003003 3.3 0.0003004 0 0.00030031999999999997 0 0.00030042 3.3 0.00030034 3.3 0.00030044 0 0.00030036 0 0.00030046 3.3 0.00030038 3.3 0.00030048 0 0.0003004 0 0.0003005 3.3 0.00030042 3.3 0.00030052 0 0.00030044 0 0.00030054 3.3 0.00030046 3.3 0.00030056 0 0.00030048 0 0.00030058 3.3 0.0003005 3.3 0.0003006 0 0.00030052 0 0.00030062 3.3 0.00030053999999999997 3.3 0.00030063999999999997 0 0.00030056 0 0.00030066 3.3 0.00030058 3.3 0.00030068 0 0.0003006 0 0.0003007 3.3 0.00030062 3.3 0.00030072 0 0.00030063999999999997 0 0.00030073999999999997 3.3 0.00030066 3.3 0.00030076 0 0.00030068 0 0.00030078 3.3 0.0003007 3.3 0.0003008 0 0.00030072 0 0.00030082 3.3 0.00030073999999999997 3.3 0.00030083999999999997 0 0.00030076 0 0.00030086 3.3 0.00030078 3.3 0.00030088 0 0.0003008 0 0.0003009 3.3 0.00030082 3.3 0.00030092 0 0.00030083999999999997 0 0.00030094 3.3 0.00030086 3.3 0.00030096 0 0.00030088 0 0.00030098 3.3 0.0003009 3.3 0.000301 0 0.00030092 0 0.00030102 3.3 0.00030094 3.3 0.00030104 0 0.00030095999999999996 0 0.00030105999999999997 3.3 0.00030098 3.3 0.00030108 0 0.000301 0 0.0003011 3.3 0.00030102 3.3 0.00030112 0 0.00030104 0 0.00030114 3.3 0.00030105999999999997 3.3 0.00030115999999999997 0 0.00030108 0 0.00030118 3.3 0.0003011 3.3 0.0003012 0 0.00030112 0 0.00030122 3.3 0.00030114 3.3 0.00030124 0 0.00030115999999999997 0 0.00030125999999999997 3.3 0.00030118 3.3 0.00030128 0 0.0003012 0 0.0003013 3.3 0.00030122 3.3 0.00030132 0 0.00030124 0 0.00030134 3.3 0.00030125999999999997 3.3 0.00030136 0 0.00030128 0 0.00030138 3.3 0.0003013 3.3 0.0003014 0 0.00030132 0 0.00030142 3.3 0.00030134 3.3 0.00030144 0 0.00030136 0 0.00030146 3.3 0.00030138 3.3 0.00030148 0 0.0003014 0 0.0003015 3.3 0.00030142 3.3 0.00030152 0 0.00030144 0 0.00030154 3.3 0.00030146 3.3 0.00030156 0 0.00030147999999999997 0 0.00030157999999999997 3.3 0.0003015 3.3 0.0003016 0 0.00030152 0 0.00030162 3.3 0.00030154 3.3 0.00030164 0 0.00030156 0 0.00030166 3.3 0.00030157999999999997 3.3 0.00030167999999999997 0 0.0003016 0 0.0003017 3.3 0.00030162 3.3 0.00030172 0 0.00030164 0 0.00030174 3.3 0.00030166 3.3 0.00030176 0 0.00030167999999999997 0 0.00030178 3.3 0.0003017 3.3 0.0003018 0 0.00030172 0 0.00030182 3.3 0.00030174 3.3 0.00030184 0 0.00030176 0 0.00030186 3.3 0.00030178 3.3 0.00030188 0 0.0003018 0 0.0003019 3.3 0.00030182 3.3 0.00030192 0 0.00030184 0 0.00030194 3.3 0.00030186 3.3 0.00030196 0 0.00030188 0 0.00030198 3.3 0.00030189999999999997 3.3 0.00030199999999999997 0 0.00030192 0 0.00030202 3.3 0.00030194 3.3 0.00030204 0 0.00030196 0 0.00030206 3.3 0.00030198 3.3 0.00030208 0 0.00030199999999999997 0 0.00030209999999999997 3.3 0.00030202 3.3 0.00030212 0 0.00030204 0 0.00030214 3.3 0.00030206 3.3 0.00030216 0 0.00030208 0 0.00030218 3.3 0.00030209999999999997 3.3 0.0003022 0 0.00030212 0 0.00030222 3.3 0.00030214 3.3 0.00030224 0 0.00030216 0 0.00030226 3.3 0.00030218 3.3 0.00030228 0 0.0003022 0 0.0003023 3.3 0.00030222 3.3 0.00030232 0 0.00030224 0 0.00030234 3.3 0.00030226 3.3 0.00030236 0 0.00030228 0 0.00030238 3.3 0.0003023 3.3 0.0003024 0 0.00030231999999999997 0 0.00030241999999999997 3.3 0.00030234 3.3 0.00030244 0 0.00030236 0 0.00030246 3.3 0.00030238 3.3 0.00030248 0 0.0003024 0 0.0003025 3.3 0.00030241999999999997 3.3 0.00030251999999999997 0 0.00030244 0 0.00030254 3.3 0.00030246 3.3 0.00030256 0 0.00030248 0 0.00030258 3.3 0.0003025 3.3 0.0003026 0 0.00030251999999999997 0 0.00030261999999999997 3.3 0.00030254 3.3 0.00030264 0 0.00030256 0 0.00030266 3.3 0.00030258 3.3 0.00030268 0 0.0003026 0 0.0003027 3.3 0.00030261999999999997 3.3 0.00030272 0 0.00030264 0 0.00030274 3.3 0.00030266 3.3 0.00030276 0 0.00030268 0 0.00030278 3.3 0.0003027 3.3 0.0003028 0 0.00030272 0 0.00030282 3.3 0.00030273999999999996 3.3 0.00030283999999999997 0 0.00030276 0 0.00030286 3.3 0.00030278 3.3 0.00030288 0 0.0003028 0 0.0003029 3.3 0.00030282 3.3 0.00030292 0 0.00030283999999999997 0 0.00030293999999999997 3.3 0.00030286 3.3 0.00030296 0 0.00030288 0 0.00030298 3.3 0.0003029 3.3 0.000303 0 0.00030292 0 0.00030302 3.3 0.00030293999999999997 3.3 0.00030303999999999997 0 0.00030296 0 0.00030306 3.3 0.00030298 3.3 0.00030308 0 0.000303 0 0.0003031 3.3 0.00030302 3.3 0.00030312 0 0.00030303999999999997 0 0.00030314 3.3 0.00030306 3.3 0.00030316 0 0.00030308 0 0.00030318 3.3 0.0003031 3.3 0.0003032 0 0.00030312 0 0.00030322 3.3 0.00030314 3.3 0.00030324 0 0.00030316 0 0.00030326 3.3 0.00030318 3.3 0.00030328 0 0.0003032 0 0.0003033 3.3 0.00030322 3.3 0.00030332 0 0.00030324 0 0.00030334 3.3 0.00030325999999999997 3.3 0.00030335999999999997 0 0.00030328 0 0.00030338 3.3 0.0003033 3.3 0.0003034 0 0.00030332 0 0.00030342 3.3 0.00030334 3.3 0.00030344 0 0.00030335999999999997 0 0.00030345999999999997 3.3 0.00030338 3.3 0.00030348 0 0.0003034 0 0.0003035 3.3 0.00030342 3.3 0.00030352 0 0.00030344 0 0.00030354 3.3 0.00030345999999999997 3.3 0.00030356 0 0.00030348 0 0.00030358 3.3 0.0003035 3.3 0.0003036 0 0.00030352 0 0.00030362 3.3 0.00030354 3.3 0.00030364 0 0.00030356 0 0.00030366 3.3 0.00030358 3.3 0.00030368 0 0.0003036 0 0.0003037 3.3 0.00030362 3.3 0.00030372 0 0.00030364 0 0.00030374 3.3 0.00030366 3.3 0.00030376 0 0.00030367999999999997 0 0.00030377999999999997 3.3 0.0003037 3.3 0.0003038 0 0.00030372 0 0.00030382 3.3 0.00030374 3.3 0.00030384 0 0.00030376 0 0.00030386 3.3 0.00030377999999999997 3.3 0.00030387999999999997 0 0.0003038 0 0.0003039 3.3 0.00030382 3.3 0.00030392 0 0.00030384 0 0.00030394 3.3 0.00030386 3.3 0.00030396 0 0.00030387999999999997 0 0.00030397999999999997 3.3 0.0003039 3.3 0.000304 0 0.00030392 0 0.00030402 3.3 0.00030394 3.3 0.00030404 0 0.00030396 0 0.00030406 3.3 0.00030397999999999997 3.3 0.00030408 0 0.000304 0 0.0003041 3.3 0.00030402 3.3 0.00030412 0 0.00030404 0 0.00030414 3.3 0.00030406 3.3 0.00030416 0 0.00030408 0 0.00030418 3.3 0.00030409999999999996 3.3 0.00030419999999999997 0 0.00030412 0 0.00030422 3.3 0.00030414 3.3 0.00030424 0 0.00030416 0 0.00030426 3.3 0.00030418 3.3 0.00030428 0 0.00030419999999999997 0 0.00030429999999999997 3.3 0.00030422 3.3 0.00030432 0 0.00030424 0 0.00030434 3.3 0.00030426 3.3 0.00030436 0 0.00030428 0 0.00030438 3.3 0.00030429999999999997 3.3 0.00030439999999999997 0 0.00030432 0 0.00030442 3.3 0.00030434 3.3 0.00030444 0 0.00030436 0 0.00030446 3.3 0.00030438 3.3 0.00030448 0 0.00030439999999999997 0 0.0003045 3.3 0.00030442 3.3 0.00030452 0 0.00030444 0 0.00030454 3.3 0.00030446 3.3 0.00030456 0 0.00030448 0 0.00030458 3.3 0.0003045 3.3 0.0003046 0 0.00030452 0 0.00030462 3.3 0.00030454 3.3 0.00030464 0 0.00030456 0 0.00030466 3.3 0.00030458 3.3 0.00030468 0 0.0003046 0 0.0003047 3.3 0.00030461999999999997 3.3 0.00030471999999999997 0 0.00030464 0 0.00030474 3.3 0.00030466 3.3 0.00030476 0 0.00030468 0 0.00030478 3.3 0.0003047 3.3 0.0003048 0 0.00030471999999999997 0 0.00030481999999999997 3.3 0.00030474 3.3 0.00030484 0 0.00030476 0 0.00030486 3.3 0.00030478 3.3 0.00030488 0 0.0003048 0 0.0003049 3.3 0.00030481999999999997 3.3 0.00030492 0 0.00030484 0 0.00030494 3.3 0.00030486 3.3 0.00030496 0 0.00030488 0 0.00030498 3.3 0.0003049 3.3 0.000305 0 0.00030492 0 0.00030502 3.3 0.00030494 3.3 0.00030504 0 0.00030496 0 0.00030506 3.3 0.00030498 3.3 0.00030508 0 0.000305 0 0.0003051 3.3 0.00030502 3.3 0.00030512 0 0.00030503999999999997 0 0.00030513999999999997 3.3 0.00030506 3.3 0.00030516 0 0.00030508 0 0.00030518 3.3 0.0003051 3.3 0.0003052 0 0.00030512 0 0.00030522 3.3 0.00030513999999999997 3.3 0.00030523999999999997 0 0.00030516 0 0.00030526 3.3 0.00030518 3.3 0.00030528 0 0.0003052 0 0.0003053 3.3 0.00030522 3.3 0.00030532 0 0.00030523999999999997 0 0.00030534 3.3 0.00030526 3.3 0.00030536 0 0.00030528 0 0.00030538 3.3 0.0003053 3.3 0.0003054 0 0.00030532 0 0.00030542 3.3 0.00030534 3.3 0.00030544 0 0.00030536 0 0.00030546 3.3 0.00030538 3.3 0.00030548 0 0.0003054 0 0.0003055 3.3 0.00030542 3.3 0.00030552 0 0.00030544 0 0.00030554 3.3 0.00030545999999999997 3.3 0.00030555999999999997 0 0.00030548 0 0.00030558 3.3 0.0003055 3.3 0.0003056 0 0.00030552 0 0.00030562 3.3 0.00030554 3.3 0.00030564 0 0.00030555999999999997 0 0.00030565999999999997 3.3 0.00030558 3.3 0.00030568 0 0.0003056 0 0.0003057 3.3 0.00030562 3.3 0.00030572 0 0.00030564 0 0.00030574 3.3 0.00030565999999999997 3.3 0.00030575999999999997 0 0.00030568 0 0.00030578 3.3 0.0003057 3.3 0.0003058 0 0.00030572 0 0.00030582 3.3 0.00030574 3.3 0.00030584 0 0.00030575999999999997 0 0.00030586 3.3 0.00030578 3.3 0.00030588 0 0.0003058 0 0.0003059 3.3 0.00030582 3.3 0.00030592 0 0.00030584 0 0.00030594 3.3 0.00030586 3.3 0.00030596 0 0.00030587999999999996 0 0.00030597999999999997 3.3 0.0003059 3.3 0.000306 0 0.00030592 0 0.00030602 3.3 0.00030594 3.3 0.00030604 0 0.00030596 0 0.00030606 3.3 0.00030597999999999997 3.3 0.00030607999999999997 0 0.000306 0 0.0003061 3.3 0.00030602 3.3 0.00030612 0 0.00030604 0 0.00030614 3.3 0.00030606 3.3 0.00030616 0 0.00030607999999999997 0 0.00030617999999999997 3.3 0.0003061 3.3 0.0003062 0 0.00030612 0 0.00030622 3.3 0.00030614 3.3 0.00030624 0 0.00030616 0 0.00030626 3.3 0.00030617999999999997 3.3 0.00030628 0 0.0003062 0 0.0003063 3.3 0.00030622 3.3 0.00030632 0 0.00030624 0 0.00030634 3.3 0.00030626 3.3 0.00030636 0 0.00030628 0 0.00030638 3.3 0.0003063 3.3 0.0003064 0 0.00030632 0 0.00030642 3.3 0.00030634 3.3 0.00030644 0 0.00030636 0 0.00030646 3.3 0.00030638 3.3 0.00030648 0 0.00030639999999999997 0 0.00030649999999999997 3.3 0.00030642 3.3 0.00030652 0 0.00030644 0 0.00030654 3.3 0.00030646 3.3 0.00030656 0 0.00030648 0 0.00030658 3.3 0.00030649999999999997 3.3 0.00030659999999999997 0 0.00030652 0 0.00030662 3.3 0.00030654 3.3 0.00030664 0 0.00030656 0 0.00030666 3.3 0.00030658 3.3 0.00030668 0 0.00030659999999999997 0 0.0003067 3.3 0.00030662 3.3 0.00030672 0 0.00030664 0 0.00030674 3.3 0.00030666 3.3 0.00030676 0 0.00030668 0 0.00030678 3.3 0.0003067 3.3 0.0003068 0 0.00030672 0 0.00030682 3.3 0.00030674 3.3 0.00030684 0 0.00030676 0 0.00030686 3.3 0.00030678 3.3 0.00030688 0 0.0003068 0 0.0003069 3.3 0.00030681999999999997 3.3 0.00030691999999999997 0 0.00030684 0 0.00030694 3.3 0.00030686 3.3 0.00030696 0 0.00030688 0 0.00030698 3.3 0.0003069 3.3 0.000307 0 0.00030691999999999997 0 0.00030701999999999997 3.3 0.00030694 3.3 0.00030704 0 0.00030696 0 0.00030706 3.3 0.00030698 3.3 0.00030708 0 0.000307 0 0.0003071 3.3 0.00030701999999999997 3.3 0.00030712 0 0.00030704 0 0.00030714 3.3 0.00030706 3.3 0.00030716 0 0.00030708 0 0.00030718 3.3 0.0003071 3.3 0.0003072 0 0.00030712 0 0.00030722 3.3 0.00030714 3.3 0.00030724 0 0.00030716 0 0.00030726 3.3 0.00030718 3.3 0.00030728 0 0.0003072 0 0.0003073 3.3 0.00030722 3.3 0.00030732 0 0.00030723999999999997 0 0.00030733999999999997 3.3 0.00030726 3.3 0.00030736 0 0.00030728 0 0.00030738 3.3 0.0003073 3.3 0.0003074 0 0.00030732 0 0.00030742 3.3 0.00030733999999999997 3.3 0.00030743999999999997 0 0.00030736 0 0.00030746 3.3 0.00030738 3.3 0.00030748 0 0.0003074 0 0.0003075 3.3 0.00030742 3.3 0.00030752 0 0.00030743999999999997 0 0.00030753999999999997 3.3 0.00030746 3.3 0.00030756 0 0.00030748 0 0.00030758 3.3 0.0003075 3.3 0.0003076 0 0.00030752 0 0.00030762 3.3 0.00030753999999999997 3.3 0.00030764 0 0.00030756 0 0.00030766 3.3 0.00030758 3.3 0.00030768 0 0.0003076 0 0.0003077 3.3 0.00030762 3.3 0.00030772 0 0.00030764 0 0.00030774 3.3 0.00030765999999999996 3.3 0.00030775999999999997 0 0.00030768 0 0.00030778 3.3 0.0003077 3.3 0.0003078 0 0.00030772 0 0.00030782 3.3 0.00030774 3.3 0.00030784 0 0.00030775999999999997 0 0.00030785999999999997 3.3 0.00030778 3.3 0.00030788 0 0.0003078 0 0.0003079 3.3 0.00030782 3.3 0.00030792 0 0.00030784 0 0.00030794 3.3 0.00030785999999999997 3.3 0.00030795999999999997 0 0.00030788 0 0.00030798 3.3 0.0003079 3.3 0.000308 0 0.00030792 0 0.00030802 3.3 0.00030794 3.3 0.00030804 0 0.00030795999999999997 0 0.00030806 3.3 0.00030798 3.3 0.00030808 0 0.000308 0 0.0003081 3.3 0.00030802 3.3 0.00030812 0 0.00030804 0 0.00030814 3.3 0.00030806 3.3 0.00030816 0 0.00030808 0 0.00030818 3.3 0.0003081 3.3 0.0003082 0 0.00030812 0 0.00030822 3.3 0.00030814 3.3 0.00030824 0 0.00030816 0 0.00030826 3.3 0.00030817999999999997 3.3 0.00030827999999999997 0 0.0003082 0 0.0003083 3.3 0.00030822 3.3 0.00030832 0 0.00030824 0 0.00030834 3.3 0.00030826 3.3 0.00030836 0 0.00030827999999999997 0 0.00030837999999999997 3.3 0.0003083 3.3 0.0003084 0 0.00030832 0 0.00030842 3.3 0.00030834 3.3 0.00030844 0 0.00030836 0 0.00030846 3.3 0.00030837999999999997 3.3 0.00030848 0 0.0003084 0 0.0003085 3.3 0.00030842 3.3 0.00030852 0 0.00030844 0 0.00030854 3.3 0.00030846 3.3 0.00030856 0 0.00030848 0 0.00030858 3.3 0.0003085 3.3 0.0003086 0 0.00030852 0 0.00030862 3.3 0.00030854 3.3 0.00030864 0 0.00030856 0 0.00030866 3.3 0.00030858 3.3 0.00030868 0 0.00030859999999999997 0 0.00030869999999999997 3.3 0.00030862 3.3 0.00030872 0 0.00030864 0 0.00030874 3.3 0.00030866 3.3 0.00030876 0 0.00030868 0 0.00030878 3.3 0.00030869999999999997 3.3 0.00030879999999999997 0 0.00030872 0 0.00030882 3.3 0.00030874 3.3 0.00030884 0 0.00030876 0 0.00030886 3.3 0.00030878 3.3 0.00030888 0 0.00030879999999999997 0 0.0003089 3.3 0.00030882 3.3 0.00030892 0 0.00030884 0 0.00030894 3.3 0.00030886 3.3 0.00030896 0 0.00030888 0 0.00030898 3.3 0.0003089 3.3 0.000309 0 0.00030892 0 0.00030902 3.3 0.00030894 3.3 0.00030904 0 0.00030896 0 0.00030906 3.3 0.00030898 3.3 0.00030908 0 0.000309 0 0.0003091 3.3 0.00030901999999999997 3.3 0.00030911999999999997 0 0.00030904 0 0.00030914 3.3 0.00030906 3.3 0.00030916 0 0.00030908 0 0.00030918 3.3 0.0003091 3.3 0.0003092 0 0.00030911999999999997 0 0.00030921999999999997 3.3 0.00030914 3.3 0.00030924 0 0.00030916 0 0.00030926 3.3 0.00030918 3.3 0.00030928 0 0.0003092 0 0.0003093 3.3 0.00030921999999999997 3.3 0.00030931999999999997 0 0.00030924 0 0.00030934 3.3 0.00030926 3.3 0.00030936 0 0.00030928 0 0.00030938 3.3 0.0003093 3.3 0.0003094 0 0.00030931999999999997 0 0.00030942 3.3 0.00030934 3.3 0.00030944 0 0.00030936 0 0.00030946 3.3 0.00030938 3.3 0.00030948 0 0.0003094 0 0.0003095 3.3 0.00030942 3.3 0.00030952 0 0.00030943999999999996 0 0.00030953999999999997 3.3 0.00030946 3.3 0.00030956 0 0.00030948 0 0.00030958 3.3 0.0003095 3.3 0.0003096 0 0.00030952 0 0.00030962 3.3 0.00030953999999999997 3.3 0.00030963999999999997 0 0.00030956 0 0.00030966 3.3 0.00030958 3.3 0.00030968 0 0.0003096 0 0.0003097 3.3 0.00030962 3.3 0.00030972 0 0.00030963999999999997 0 0.00030973999999999997 3.3 0.00030966 3.3 0.00030976 0 0.00030968 0 0.00030978 3.3 0.0003097 3.3 0.0003098 0 0.00030972 0 0.00030982 3.3 0.00030973999999999997 3.3 0.00030984 0 0.00030976 0 0.00030986 3.3 0.00030978 3.3 0.00030988 0 0.0003098 0 0.0003099 3.3 0.00030982 3.3 0.00030992 0 0.00030984 0 0.00030994 3.3 0.00030986 3.3 0.00030996 0 0.00030988 0 0.00030998 3.3 0.0003099 3.3 0.00031 0 0.00030992 0 0.00031002 3.3 0.00030994 3.3 0.00031004 0 0.00030995999999999997 0 0.00031005999999999997 3.3 0.00030998 3.3 0.00031008 0 0.00031 0 0.0003101 3.3 0.00031002 3.3 0.00031012 0 0.00031004 0 0.00031014 3.3 0.00031005999999999997 3.3 0.00031015999999999997 0 0.00031008 0 0.00031018 3.3 0.0003101 3.3 0.0003102 0 0.00031012 0 0.00031022 3.3 0.00031014 3.3 0.00031024 0 0.00031015999999999997 0 0.00031026 3.3 0.00031018 3.3 0.00031028 0 0.0003102 0 0.0003103 3.3 0.00031022 3.3 0.00031032 0 0.00031024 0 0.00031034 3.3 0.00031026 3.3 0.00031036 0 0.00031028 0 0.00031038 3.3 0.0003103 3.3 0.0003104 0 0.00031032 0 0.00031042 3.3 0.00031034 3.3 0.00031044 0 0.00031036 0 0.00031046 3.3 0.00031037999999999997 3.3 0.00031047999999999997 0 0.0003104 0 0.0003105 3.3 0.00031042 3.3 0.00031052 0 0.00031044 0 0.00031054 3.3 0.00031046 3.3 0.00031056 0 0.00031047999999999997 0 0.00031057999999999997 3.3 0.0003105 3.3 0.0003106 0 0.00031052 0 0.00031062 3.3 0.00031054 3.3 0.00031064 0 0.00031056 0 0.00031066 3.3 0.00031057999999999997 3.3 0.00031068 0 0.0003106 0 0.0003107 3.3 0.00031062 3.3 0.00031072 0 0.00031064 0 0.00031074 3.3 0.00031066 3.3 0.00031076 0 0.00031068 0 0.00031078 3.3 0.0003107 3.3 0.0003108 0 0.00031072 0 0.00031082 3.3 0.00031074 3.3 0.00031084 0 0.00031076 0 0.00031086 3.3 0.00031078 3.3 0.00031088 0 0.00031079999999999997 0 0.00031089999999999997 3.3 0.00031082 3.3 0.00031092 0 0.00031084 0 0.00031094 3.3 0.00031086 3.3 0.00031096 0 0.00031088 0 0.00031098 3.3 0.00031089999999999997 3.3 0.00031099999999999997 0 0.00031092 0 0.00031102 3.3 0.00031094 3.3 0.00031104 0 0.00031096 0 0.00031106 3.3 0.00031098 3.3 0.00031108 0 0.00031099999999999997 0 0.00031109999999999997 3.3 0.00031102 3.3 0.00031112 0 0.00031104 0 0.00031114 3.3 0.00031106 3.3 0.00031116 0 0.00031108 0 0.00031118 3.3 0.00031109999999999997 3.3 0.0003112 0 0.00031112 0 0.00031122 3.3 0.00031114 3.3 0.00031124 0 0.00031116 0 0.00031126 3.3 0.00031118 3.3 0.00031128 0 0.0003112 0 0.0003113 3.3 0.00031121999999999996 3.3 0.00031131999999999997 0 0.00031124 0 0.00031134 3.3 0.00031126 3.3 0.00031136 0 0.00031128 0 0.00031138 3.3 0.0003113 3.3 0.0003114 0 0.00031131999999999997 0 0.00031141999999999997 3.3 0.00031134 3.3 0.00031144 0 0.00031136 0 0.00031146 3.3 0.00031138 3.3 0.00031148 0 0.0003114 0 0.0003115 3.3 0.00031141999999999997 3.3 0.00031151999999999997 0 0.00031144 0 0.00031154 3.3 0.00031146 3.3 0.00031156 0 0.00031148 0 0.00031158 3.3 0.0003115 3.3 0.0003116 0 0.00031151999999999997 0 0.00031162 3.3 0.00031154 3.3 0.00031164 0 0.00031156 0 0.00031166 3.3 0.00031158 3.3 0.00031168 0 0.0003116 0 0.0003117 3.3 0.00031162 3.3 0.00031172 0 0.00031164 0 0.00031174 3.3 0.00031166 3.3 0.00031176 0 0.00031168 0 0.00031178 3.3 0.0003117 3.3 0.0003118 0 0.00031172 0 0.00031182 3.3 0.00031173999999999997 3.3 0.00031183999999999997 0 0.00031176 0 0.00031186 3.3 0.00031178 3.3 0.00031188 0 0.0003118 0 0.0003119 3.3 0.00031182 3.3 0.00031192 0 0.00031183999999999997 0 0.00031193999999999997 3.3 0.00031186 3.3 0.00031196 0 0.00031188 0 0.00031198 3.3 0.0003119 3.3 0.000312 0 0.00031192 0 0.00031202 3.3 0.00031193999999999997 3.3 0.00031204 0 0.00031196 0 0.00031206 3.3 0.00031198 3.3 0.00031208 0 0.000312 0 0.0003121 3.3 0.00031202 3.3 0.00031212 0 0.00031204 0 0.00031214 3.3 0.00031206 3.3 0.00031216 0 0.00031208 0 0.00031218 3.3 0.0003121 3.3 0.0003122 0 0.00031212 0 0.00031222 3.3 0.00031214 3.3 0.00031224 0 0.00031215999999999997 0 0.00031225999999999997 3.3 0.00031218 3.3 0.00031228 0 0.0003122 0 0.0003123 3.3 0.00031222 3.3 0.00031232 0 0.00031224 0 0.00031234 3.3 0.00031225999999999997 3.3 0.00031235999999999997 0 0.00031228 0 0.00031238 3.3 0.0003123 3.3 0.0003124 0 0.00031232 0 0.00031242 3.3 0.00031234 3.3 0.00031244 0 0.00031235999999999997 0 0.00031246 3.3 0.00031238 3.3 0.00031248 0 0.0003124 0 0.0003125 3.3 0.00031242 3.3 0.00031252 0 0.00031244 0 0.00031254 3.3 0.00031246 3.3 0.00031256 0 0.00031248 0 0.00031258 3.3 0.0003125 3.3 0.0003126 0 0.00031252 0 0.00031262 3.3 0.00031254 3.3 0.00031264 0 0.00031256 0 0.00031266 3.3 0.00031257999999999997 3.3 0.00031267999999999997 0 0.0003126 0 0.0003127 3.3 0.00031262 3.3 0.00031272 0 0.00031264 0 0.00031274 3.3 0.00031266 3.3 0.00031276 0 0.00031267999999999997 0 0.00031277999999999997 3.3 0.0003127 3.3 0.0003128 0 0.00031272 0 0.00031282 3.3 0.00031274 3.3 0.00031284 0 0.00031276 0 0.00031286 3.3 0.00031277999999999997 3.3 0.00031287999999999997 0 0.0003128 0 0.0003129 3.3 0.00031282 3.3 0.00031292 0 0.00031284 0 0.00031294 3.3 0.00031286 3.3 0.00031296 0 0.00031287999999999997 0 0.00031298 3.3 0.0003129 3.3 0.000313 0 0.00031292 0 0.00031302 3.3 0.00031294 3.3 0.00031304 0 0.00031296 0 0.00031306 3.3 0.00031298 3.3 0.00031308 0 0.00031299999999999996 0 0.00031309999999999997 3.3 0.00031302 3.3 0.00031312 0 0.00031304 0 0.00031314 3.3 0.00031306 3.3 0.00031316 0 0.00031308 0 0.00031318 3.3 0.00031309999999999997 3.3 0.00031319999999999997 0 0.00031312 0 0.00031322 3.3 0.00031314 3.3 0.00031324 0 0.00031316 0 0.00031326 3.3 0.00031318 3.3 0.00031328 0 0.00031319999999999997 0 0.00031329999999999997 3.3 0.00031322 3.3 0.00031332 0 0.00031324 0 0.00031334 3.3 0.00031326 3.3 0.00031336 0 0.00031328 0 0.00031338 3.3 0.00031329999999999997 3.3 0.0003134 0 0.00031332 0 0.00031342 3.3 0.00031334 3.3 0.00031344 0 0.00031336 0 0.00031346 3.3 0.00031338 3.3 0.00031348 0 0.0003134 0 0.0003135 3.3 0.00031342 3.3 0.00031352 0 0.00031344 0 0.00031354 3.3 0.00031346 3.3 0.00031356 0 0.00031348 0 0.00031358 3.3 0.0003135 3.3 0.0003136 0 0.00031351999999999997 0 0.00031361999999999997 3.3 0.00031354 3.3 0.00031364 0 0.00031356 0 0.00031366 3.3 0.00031358 3.3 0.00031368 0 0.0003136 0 0.0003137 3.3 0.00031361999999999997 3.3 0.00031371999999999997 0 0.00031364 0 0.00031374 3.3 0.00031366 3.3 0.00031376 0 0.00031368 0 0.00031378 3.3 0.0003137 3.3 0.0003138 0 0.00031371999999999997 0 0.00031382 3.3 0.00031374 3.3 0.00031384 0 0.00031376 0 0.00031386 3.3 0.00031378 3.3 0.00031388 0 0.0003138 0 0.0003139 3.3 0.00031382 3.3 0.00031392 0 0.00031384 0 0.00031394 3.3 0.00031386 3.3 0.00031396 0 0.00031388 0 0.00031398 3.3 0.0003139 3.3 0.000314 0 0.00031392 0 0.00031402 3.3 0.00031393999999999997 3.3 0.00031403999999999997 0 0.00031396 0 0.00031406 3.3 0.00031398 3.3 0.00031408 0 0.000314 0 0.0003141 3.3 0.00031402 3.3 0.00031412 0 0.00031403999999999997 0 0.00031413999999999997 3.3 0.00031406 3.3 0.00031416 0 0.00031408 0 0.00031418 3.3 0.0003141 3.3 0.0003142 0 0.00031412 0 0.00031422 3.3 0.00031413999999999997 3.3 0.00031424 0 0.00031416 0 0.00031426 3.3 0.00031418 3.3 0.00031428 0 0.0003142 0 0.0003143 3.3 0.00031422 3.3 0.00031432 0 0.00031424 0 0.00031434 3.3 0.00031426 3.3 0.00031436 0 0.00031428 0 0.00031438 3.3 0.0003143 3.3 0.0003144 0 0.00031432 0 0.00031442 3.3 0.00031434 3.3 0.00031444 0 0.00031435999999999996 0 0.00031445999999999997 3.3 0.00031438 3.3 0.00031448 0 0.0003144 0 0.0003145 3.3 0.00031442 3.3 0.00031452 0 0.00031444 0 0.00031454 3.3 0.00031445999999999997 3.3 0.00031455999999999997 0 0.00031448 0 0.00031458 3.3 0.0003145 3.3 0.0003146 0 0.00031452 0 0.00031462 3.3 0.00031454 3.3 0.00031464 0 0.00031455999999999997 0 0.00031465999999999997 3.3 0.00031458 3.3 0.00031468 0 0.0003146 0 0.0003147 3.3 0.00031462 3.3 0.00031472 0 0.00031464 0 0.00031474 3.3 0.00031465999999999997 3.3 0.00031476 0 0.00031468 0 0.00031478 3.3 0.0003147 3.3 0.0003148 0 0.00031472 0 0.00031482 3.3 0.00031474 3.3 0.00031484 0 0.00031476 0 0.00031486 3.3 0.00031477999999999996 3.3 0.00031487999999999997 0 0.0003148 0 0.0003149 3.3 0.00031482 3.3 0.00031492 0 0.00031484 0 0.00031494 3.3 0.00031486 3.3 0.00031496 0 0.00031487999999999997 0 0.00031497999999999997 3.3 0.0003149 3.3 0.000315 0 0.00031492 0 0.00031502 3.3 0.00031494 3.3 0.00031504 0 0.00031496 0 0.00031506 3.3 0.00031497999999999997 3.3 0.00031507999999999997 0 0.000315 0 0.0003151 3.3 0.00031502 3.3 0.00031512 0 0.00031504 0 0.00031514 3.3 0.00031506 3.3 0.00031516 0 0.00031507999999999997 0 0.00031518 3.3 0.0003151 3.3 0.0003152 0 0.00031512 0 0.00031522 3.3 0.00031514 3.3 0.00031524 0 0.00031516 0 0.00031526 3.3 0.00031518 3.3 0.00031528 0 0.0003152 0 0.0003153 3.3 0.00031522 3.3 0.00031532 0 0.00031524 0 0.00031534 3.3 0.00031526 3.3 0.00031536 0 0.00031528 0 0.00031538 3.3 0.00031529999999999997 3.3 0.00031539999999999997 0 0.00031532 0 0.00031542 3.3 0.00031534 3.3 0.00031544 0 0.00031536 0 0.00031546 3.3 0.00031538 3.3 0.00031548 0 0.00031539999999999997 0 0.00031549999999999997 3.3 0.00031542 3.3 0.00031552 0 0.00031544 0 0.00031554 3.3 0.00031546 3.3 0.00031556 0 0.00031548 0 0.00031558 3.3 0.00031549999999999997 3.3 0.0003156 0 0.00031552 0 0.00031562 3.3 0.00031554 3.3 0.00031564 0 0.00031556 0 0.00031566 3.3 0.00031558 3.3 0.00031568 0 0.0003156 0 0.0003157 3.3 0.00031562 3.3 0.00031572 0 0.00031564 0 0.00031574 3.3 0.00031566 3.3 0.00031576 0 0.00031568 0 0.00031578 3.3 0.0003157 3.3 0.0003158 0 0.00031571999999999997 0 0.00031581999999999997 3.3 0.00031574 3.3 0.00031584 0 0.00031576 0 0.00031586 3.3 0.00031578 3.3 0.00031588 0 0.0003158 0 0.0003159 3.3 0.00031581999999999997 3.3 0.00031591999999999997 0 0.00031584 0 0.00031594 3.3 0.00031586 3.3 0.00031596 0 0.00031588 0 0.00031598 3.3 0.0003159 3.3 0.000316 0 0.00031591999999999997 0 0.00031601999999999997 3.3 0.00031594 3.3 0.00031604 0 0.00031596 0 0.00031606 3.3 0.00031598 3.3 0.00031608 0 0.000316 0 0.0003161 3.3 0.00031601999999999997 3.3 0.00031612 0 0.00031604 0 0.00031614 3.3 0.00031606 3.3 0.00031616 0 0.00031608 0 0.00031618 3.3 0.0003161 3.3 0.0003162 0 0.00031612 0 0.00031622 3.3 0.00031613999999999996 3.3 0.00031623999999999997 0 0.00031616 0 0.00031626 3.3 0.00031618 3.3 0.00031628 0 0.0003162 0 0.0003163 3.3 0.00031622 3.3 0.00031632 0 0.00031623999999999997 0 0.00031633999999999997 3.3 0.00031626 3.3 0.00031636 0 0.00031628 0 0.00031638 3.3 0.0003163 3.3 0.0003164 0 0.00031632 0 0.00031642 3.3 0.00031633999999999997 3.3 0.00031643999999999997 0 0.00031636 0 0.00031646 3.3 0.00031638 3.3 0.00031648 0 0.0003164 0 0.0003165 3.3 0.00031642 3.3 0.00031652 0 0.00031643999999999997 0 0.00031654 3.3 0.00031646 3.3 0.00031656 0 0.00031648 0 0.00031658 3.3 0.0003165 3.3 0.0003166 0 0.00031652 0 0.00031662 3.3 0.00031654 3.3 0.00031664 0 0.00031655999999999996 0 0.00031665999999999997 3.3 0.00031658 3.3 0.00031668 0 0.0003166 0 0.0003167 3.3 0.00031662 3.3 0.00031672 0 0.00031664 0 0.00031674 3.3 0.00031665999999999997 3.3 0.00031675999999999997 0 0.00031668 0 0.00031678 3.3 0.0003167 3.3 0.0003168 0 0.00031672 0 0.00031682 3.3 0.00031674 3.3 0.00031684 0 0.00031675999999999997 0 0.00031685999999999997 3.3 0.00031678 3.3 0.00031688 0 0.0003168 0 0.0003169 3.3 0.00031682 3.3 0.00031692 0 0.00031684 0 0.00031694 3.3 0.00031685999999999997 3.3 0.00031696 0 0.00031688 0 0.00031698 3.3 0.0003169 3.3 0.000317 0 0.00031692 0 0.00031702 3.3 0.00031694 3.3 0.00031704 0 0.00031696 0 0.00031706 3.3 0.00031698 3.3 0.00031708 0 0.000317 0 0.0003171 3.3 0.00031702 3.3 0.00031712 0 0.00031704 0 0.00031714 3.3 0.00031706 3.3 0.00031716 0 0.00031707999999999997 0 0.00031717999999999997 3.3 0.0003171 3.3 0.0003172 0 0.00031712 0 0.00031722 3.3 0.00031714 3.3 0.00031724 0 0.00031716 0 0.00031726 3.3 0.00031717999999999997 3.3 0.00031727999999999997 0 0.0003172 0 0.0003173 3.3 0.00031722 3.3 0.00031732 0 0.00031724 0 0.00031734 3.3 0.00031726 3.3 0.00031736 0 0.00031727999999999997 0 0.00031738 3.3 0.0003173 3.3 0.0003174 0 0.00031732 0 0.00031742 3.3 0.00031734 3.3 0.00031744 0 0.00031736 0 0.00031746 3.3 0.00031738 3.3 0.00031748 0 0.0003174 0 0.0003175 3.3 0.00031742 3.3 0.00031752 0 0.00031744 0 0.00031754 3.3 0.00031746 3.3 0.00031756 0 0.00031748 0 0.00031758 3.3 0.00031749999999999997 3.3 0.00031759999999999997 0 0.00031752 0 0.00031762 3.3 0.00031754 3.3 0.00031764 0 0.00031756 0 0.00031766 3.3 0.00031758 3.3 0.00031768 0 0.00031759999999999997 0 0.00031769999999999997 3.3 0.00031762 3.3 0.00031772 0 0.00031764 0 0.00031774 3.3 0.00031766 3.3 0.00031776 0 0.00031768 0 0.00031778 3.3 0.00031769999999999997 3.3 0.00031779999999999997 0 0.00031772 0 0.00031782 3.3 0.00031774 3.3 0.00031784 0 0.00031776 0 0.00031786 3.3 0.00031778 3.3 0.00031788 0 0.00031779999999999997 0 0.0003179 3.3 0.00031782 3.3 0.00031792 0 0.00031784 0 0.00031794 3.3 0.00031786 3.3 0.00031796 0 0.00031788 0 0.00031798 3.3 0.0003179 3.3 0.000318 0 0.00031791999999999996 0 0.00031801999999999997 3.3 0.00031794 3.3 0.00031804 0 0.00031796 0 0.00031806 3.3 0.00031798 3.3 0.00031808 0 0.000318 0 0.0003181 3.3 0.00031801999999999997 3.3 0.00031811999999999997 0 0.00031804 0 0.00031814 3.3 0.00031806 3.3 0.00031816 0 0.00031808 0 0.00031818 3.3 0.0003181 3.3 0.0003182 0 0.00031811999999999997 0 0.00031821999999999997 3.3 0.00031814 3.3 0.00031824 0 0.00031816 0 0.00031826 3.3 0.00031818 3.3 0.00031828 0 0.0003182 0 0.0003183 3.3 0.00031821999999999997 3.3 0.00031832 0 0.00031824 0 0.00031834 3.3 0.00031826 3.3 0.00031836 0 0.00031828 0 0.00031838 3.3 0.0003183 3.3 0.0003184 0 0.00031832 0 0.00031842 3.3 0.00031833999999999996 3.3 0.00031843999999999997 0 0.00031836 0 0.00031846 3.3 0.00031838 3.3 0.00031848 0 0.0003184 0 0.0003185 3.3 0.00031842 3.3 0.00031852 0 0.00031843999999999997 0 0.00031853999999999997 3.3 0.00031846 3.3 0.00031856 0 0.00031848 0 0.00031858 3.3 0.0003185 3.3 0.0003186 0 0.00031852 0 0.00031862 3.3 0.00031853999999999997 3.3 0.00031863999999999997 0 0.00031856 0 0.00031866 3.3 0.00031858 3.3 0.00031868 0 0.0003186 0 0.0003187 3.3 0.00031862 3.3 0.00031872 0 0.00031863999999999997 0 0.00031874 3.3 0.00031866 3.3 0.00031876 0 0.00031868 0 0.00031878 3.3 0.0003187 3.3 0.0003188 0 0.00031872 0 0.00031882 3.3 0.00031874 3.3 0.00031884 0 0.00031876 0 0.00031886 3.3 0.00031878 3.3 0.00031888 0 0.0003188 0 0.0003189 3.3 0.00031882 3.3 0.00031892 0 0.00031884 0 0.00031894 3.3 0.00031885999999999997 3.3 0.00031895999999999997 0 0.00031888 0 0.00031898 3.3 0.0003189 3.3 0.000319 0 0.00031892 0 0.00031902 3.3 0.00031894 3.3 0.00031904 0 0.00031895999999999997 0 0.00031905999999999997 3.3 0.00031898 3.3 0.00031908 0 0.000319 0 0.0003191 3.3 0.00031902 3.3 0.00031912 0 0.00031904 0 0.00031914 3.3 0.00031905999999999997 3.3 0.00031916 0 0.00031908 0 0.00031918 3.3 0.0003191 3.3 0.0003192 0 0.00031912 0 0.00031922 3.3 0.00031914 3.3 0.00031924 0 0.00031916 0 0.00031926 3.3 0.00031918 3.3 0.00031928 0 0.0003192 0 0.0003193 3.3 0.00031922 3.3 0.00031932 0 0.00031924 0 0.00031934 3.3 0.00031926 3.3 0.00031936 0 0.00031927999999999997 0 0.00031937999999999997 3.3 0.0003193 3.3 0.0003194 0 0.00031932 0 0.00031942 3.3 0.00031934 3.3 0.00031944 0 0.00031936 0 0.00031946 3.3 0.00031937999999999997 3.3 0.00031947999999999997 0 0.0003194 0 0.0003195 3.3 0.00031942 3.3 0.00031952 0 0.00031944 0 0.00031954 3.3 0.00031946 3.3 0.00031956 0 0.00031947999999999997 0 0.00031957999999999997 3.3 0.0003195 3.3 0.0003196 0 0.00031952 0 0.00031962 3.3 0.00031954 3.3 0.00031964 0 0.00031956 0 0.00031966 3.3 0.00031957999999999997 3.3 0.00031968 0 0.0003196 0 0.0003197 3.3 0.00031962 3.3 0.00031972 0 0.00031964 0 0.00031974 3.3 0.00031966 3.3 0.00031976 0 0.00031968 0 0.00031978 3.3 0.00031969999999999996 3.3 0.00031979999999999997 0 0.00031972 0 0.00031982 3.3 0.00031974 3.3 0.00031984 0 0.00031976 0 0.00031986 3.3 0.00031978 3.3 0.00031988 0 0.00031979999999999997 0 0.00031989999999999997 3.3 0.00031982 3.3 0.00031992 0 0.00031984 0 0.00031994 3.3 0.00031986 3.3 0.00031996 0 0.00031988 0 0.00031998 3.3 0.00031989999999999997 3.3 0.00031999999999999997 0 0.00031992 0 0.00032002 3.3 0.00031994 3.3 0.00032004 0 0.00031996 0 0.00032006 3.3 0.00031998 3.3 0.00032008 0 0.00031999999999999997 0 0.0003201 3.3 0.00032002 3.3 0.00032012 0 0.00032004 0 0.00032014 3.3 0.00032006 3.3 0.00032016 0 0.00032008 0 0.00032018 3.3 0.0003201 3.3 0.0003202 0 0.00032011999999999996 0 0.00032021999999999997 3.3 0.00032014 3.3 0.00032024 0 0.00032016 0 0.00032026 3.3 0.00032018 3.3 0.00032028 0 0.0003202 0 0.0003203 3.3 0.00032021999999999997 3.3 0.00032031999999999997 0 0.00032024 0 0.00032034 3.3 0.00032026 3.3 0.00032036 0 0.00032028 0 0.00032038 3.3 0.0003203 3.3 0.0003204 0 0.00032031999999999997 0 0.00032041999999999997 3.3 0.00032034 3.3 0.00032044 0 0.00032036 0 0.00032046 3.3 0.00032038 3.3 0.00032048 0 0.0003204 0 0.0003205 3.3 0.00032041999999999997 3.3 0.00032052 0 0.00032044 0 0.00032054 3.3 0.00032046 3.3 0.00032056 0 0.00032048 0 0.00032058 3.3 0.0003205 3.3 0.0003206 0 0.00032052 0 0.00032062 3.3 0.00032054 3.3 0.00032064 0 0.00032056 0 0.00032066 3.3 0.00032058 3.3 0.00032068 0 0.0003206 0 0.0003207 3.3 0.00032062 3.3 0.00032072 0 0.00032063999999999997 0 0.00032073999999999997 3.3 0.00032066 3.3 0.00032076 0 0.00032068 0 0.00032078 3.3 0.0003207 3.3 0.0003208 0 0.00032072 0 0.00032082 3.3 0.00032073999999999997 3.3 0.00032083999999999997 0 0.00032076 0 0.00032086 3.3 0.00032078 3.3 0.00032088 0 0.0003208 0 0.0003209 3.3 0.00032082 3.3 0.00032092 0 0.00032083999999999997 0 0.00032094 3.3 0.00032086 3.3 0.00032096 0 0.00032088 0 0.00032098 3.3 0.0003209 3.3 0.000321 0 0.00032092 0 0.00032102 3.3 0.00032094 3.3 0.00032104 0 0.00032096 0 0.00032106 3.3 0.00032098 3.3 0.00032108 0 0.000321 0 0.0003211 3.3 0.00032102 3.3 0.00032112 0 0.00032104 0 0.00032114 3.3 0.00032105999999999997 3.3 0.00032115999999999997 0 0.00032108 0 0.00032118 3.3 0.0003211 3.3 0.0003212 0 0.00032112 0 0.00032122 3.3 0.00032114 3.3 0.00032124 0 0.00032115999999999997 0 0.00032125999999999997 3.3 0.00032118 3.3 0.00032128 0 0.0003212 0 0.0003213 3.3 0.00032122 3.3 0.00032132 0 0.00032124 0 0.00032134 3.3 0.00032125999999999997 3.3 0.00032135999999999997 0 0.00032128 0 0.00032138 3.3 0.0003213 3.3 0.0003214 0 0.00032132 0 0.00032142 3.3 0.00032134 3.3 0.00032144 0 0.00032135999999999997 0 0.00032146 3.3 0.00032138 3.3 0.00032148 0 0.0003214 0 0.0003215 3.3 0.00032142 3.3 0.00032152 0 0.00032144 0 0.00032154 3.3 0.00032146 3.3 0.00032156 0 0.00032147999999999996 0 0.00032157999999999997 3.3 0.0003215 3.3 0.0003216 0 0.00032152 0 0.00032162 3.3 0.00032154 3.3 0.00032164 0 0.00032156 0 0.00032166 3.3 0.00032157999999999997 3.3 0.00032167999999999997 0 0.0003216 0 0.0003217 3.3 0.00032162 3.3 0.00032172 0 0.00032164 0 0.00032174 3.3 0.00032166 3.3 0.00032176 0 0.00032167999999999997 0 0.00032177999999999997 3.3 0.0003217 3.3 0.0003218 0 0.00032172 0 0.00032182 3.3 0.00032174 3.3 0.00032184 0 0.00032176 0 0.00032186 3.3 0.00032177999999999997 3.3 0.00032188 0 0.0003218 0 0.0003219 3.3 0.00032182 3.3 0.00032192 0 0.00032184 0 0.00032194 3.3 0.00032186 3.3 0.00032196 0 0.00032188 0 0.00032198 3.3 0.0003219 3.3 0.000322 0 0.00032192 0 0.00032202 3.3 0.00032194 3.3 0.00032204 0 0.00032196 0 0.00032206 3.3 0.00032198 3.3 0.00032208 0 0.00032199999999999997 0 0.00032209999999999997 3.3 0.00032202 3.3 0.00032212 0 0.00032204 0 0.00032214 3.3 0.00032206 3.3 0.00032216 0 0.00032208 0 0.00032218 3.3 0.00032209999999999997 3.3 0.00032219999999999997 0 0.00032212 0 0.00032222 3.3 0.00032214 3.3 0.00032224 0 0.00032216 0 0.00032226 3.3 0.00032218 3.3 0.00032228 0 0.00032219999999999997 0 0.0003223 3.3 0.00032222 3.3 0.00032232 0 0.00032224 0 0.00032234 3.3 0.00032226 3.3 0.00032236 0 0.00032228 0 0.00032238 3.3 0.0003223 3.3 0.0003224 0 0.00032232 0 0.00032242 3.3 0.00032234 3.3 0.00032244 0 0.00032236 0 0.00032246 3.3 0.00032238 3.3 0.00032248 0 0.0003224 0 0.0003225 3.3 0.00032241999999999997 3.3 0.00032251999999999997 0 0.00032244 0 0.00032254 3.3 0.00032246 3.3 0.00032256 0 0.00032248 0 0.00032258 3.3 0.0003225 3.3 0.0003226 0 0.00032251999999999997 0 0.00032261999999999997 3.3 0.00032254 3.3 0.00032264 0 0.00032256 0 0.00032266 3.3 0.00032258 3.3 0.00032268 0 0.0003226 0 0.0003227 3.3 0.00032261999999999997 3.3 0.00032272 0 0.00032264 0 0.00032274 3.3 0.00032266 3.3 0.00032276 0 0.00032268 0 0.00032278 3.3 0.0003227 3.3 0.0003228 0 0.00032272 0 0.00032282 3.3 0.00032274 3.3 0.00032284 0 0.00032276 0 0.00032286 3.3 0.00032278 3.3 0.00032288 0 0.0003228 0 0.0003229 3.3 0.00032282 3.3 0.00032292 0 0.00032283999999999997 0 0.00032293999999999997 3.3 0.00032286 3.3 0.00032296 0 0.00032288 0 0.00032298 3.3 0.0003229 3.3 0.000323 0 0.00032292 0 0.00032302 3.3 0.00032293999999999997 3.3 0.00032303999999999997 0 0.00032296 0 0.00032306 3.3 0.00032298 3.3 0.00032308 0 0.000323 0 0.0003231 3.3 0.00032302 3.3 0.00032312 0 0.00032303999999999997 0 0.00032313999999999997 3.3 0.00032306 3.3 0.00032316 0 0.00032308 0 0.00032318 3.3 0.0003231 3.3 0.0003232 0 0.00032312 0 0.00032322 3.3 0.00032313999999999997 3.3 0.00032324 0 0.00032316 0 0.00032326 3.3 0.00032318 3.3 0.00032328 0 0.0003232 0 0.0003233 3.3 0.00032322 3.3 0.00032332 0 0.00032324 0 0.00032334 3.3 0.00032325999999999996 3.3 0.00032335999999999997 0 0.00032328 0 0.00032338 3.3 0.0003233 3.3 0.0003234 0 0.00032332 0 0.00032342 3.3 0.00032334 3.3 0.00032344 0 0.00032335999999999997 0 0.00032345999999999997 3.3 0.00032338 3.3 0.00032348 0 0.0003234 0 0.0003235 3.3 0.00032342 3.3 0.00032352 0 0.00032344 0 0.00032354 3.3 0.00032345999999999997 3.3 0.00032355999999999997 0 0.00032348 0 0.00032358 3.3 0.0003235 3.3 0.0003236 0 0.00032352 0 0.00032362 3.3 0.00032354 3.3 0.00032364 0 0.00032355999999999997 0 0.00032366 3.3 0.00032358 3.3 0.00032368 0 0.0003236 0 0.0003237 3.3 0.00032362 3.3 0.00032372 0 0.00032364 0 0.00032374 3.3 0.00032366 3.3 0.00032376 0 0.00032368 0 0.00032378 3.3 0.0003237 3.3 0.0003238 0 0.00032372 0 0.00032382 3.3 0.00032374 3.3 0.00032384 0 0.00032376 0 0.00032386 3.3 0.00032377999999999997 3.3 0.00032387999999999997 0 0.0003238 0 0.0003239 3.3 0.00032382 3.3 0.00032392 0 0.00032384 0 0.00032394 3.3 0.00032386 3.3 0.00032396 0 0.00032387999999999997 0 0.00032397999999999997 3.3 0.0003239 3.3 0.000324 0 0.00032392 0 0.00032402 3.3 0.00032394 3.3 0.00032404 0 0.00032396 0 0.00032406 3.3 0.00032397999999999997 3.3 0.00032408 0 0.000324 0 0.0003241 3.3 0.00032402 3.3 0.00032412 0 0.00032404 0 0.00032414 3.3 0.00032406 3.3 0.00032416 0 0.00032408 0 0.00032418 3.3 0.0003241 3.3 0.0003242 0 0.00032412 0 0.00032422 3.3 0.00032414 3.3 0.00032424 0 0.00032416 0 0.00032426 3.3 0.00032418 3.3 0.00032428 0 0.00032419999999999997 0 0.00032429999999999997 3.3 0.00032422 3.3 0.00032432 0 0.00032424 0 0.00032434 3.3 0.00032426 3.3 0.00032436 0 0.00032428 0 0.00032438 3.3 0.00032429999999999997 3.3 0.00032439999999999997 0 0.00032432 0 0.00032442 3.3 0.00032434 3.3 0.00032444 0 0.00032436 0 0.00032446 3.3 0.00032438 3.3 0.00032448 0 0.00032439999999999997 0 0.0003245 3.3 0.00032442 3.3 0.00032452 0 0.00032444 0 0.00032454 3.3 0.00032446 3.3 0.00032456 0 0.00032448 0 0.00032458 3.3 0.0003245 3.3 0.0003246 0 0.00032452 0 0.00032462 3.3 0.00032454 3.3 0.00032464 0 0.00032456 0 0.00032466 3.3 0.00032458 3.3 0.00032468 0 0.0003246 0 0.0003247 3.3 0.00032461999999999997 3.3 0.00032471999999999997 0 0.00032464 0 0.00032474 3.3 0.00032466 3.3 0.00032476 0 0.00032468 0 0.00032478 3.3 0.0003247 3.3 0.0003248 0 0.00032471999999999997 0 0.00032481999999999997 3.3 0.00032474 3.3 0.00032484 0 0.00032476 0 0.00032486 3.3 0.00032478 3.3 0.00032488 0 0.0003248 0 0.0003249 3.3 0.00032481999999999997 3.3 0.00032491999999999997 0 0.00032484 0 0.00032494 3.3 0.00032486 3.3 0.00032496 0 0.00032488 0 0.00032498 3.3 0.0003249 3.3 0.000325 0 0.00032491999999999997 0 0.00032502 3.3 0.00032494 3.3 0.00032504 0 0.00032496 0 0.00032506 3.3 0.00032498 3.3 0.00032508 0 0.000325 0 0.0003251 3.3 0.00032502 3.3 0.00032512 0 0.00032503999999999996 0 0.00032513999999999997 3.3 0.00032506 3.3 0.00032516 0 0.00032508 0 0.00032518 3.3 0.0003251 3.3 0.0003252 0 0.00032512 0 0.00032522 3.3 0.00032513999999999997 3.3 0.00032523999999999997 0 0.00032516 0 0.00032526 3.3 0.00032518 3.3 0.00032528 0 0.0003252 0 0.0003253 3.3 0.00032522 3.3 0.00032532 0 0.00032523999999999997 0 0.00032533999999999997 3.3 0.00032526 3.3 0.00032536 0 0.00032528 0 0.00032538 3.3 0.0003253 3.3 0.0003254 0 0.00032532 0 0.00032542 3.3 0.00032533999999999997 3.3 0.00032544 0 0.00032536 0 0.00032546 3.3 0.00032538 3.3 0.00032548 0 0.0003254 0 0.0003255 3.3 0.00032542 3.3 0.00032552 0 0.00032544 0 0.00032554 3.3 0.00032546 3.3 0.00032556 0 0.00032548 0 0.00032558 3.3 0.0003255 3.3 0.0003256 0 0.00032552 0 0.00032562 3.3 0.00032554 3.3 0.00032564 0 0.00032555999999999997 0 0.00032565999999999997 3.3 0.00032558 3.3 0.00032568 0 0.0003256 0 0.0003257 3.3 0.00032562 3.3 0.00032572 0 0.00032564 0 0.00032574 3.3 0.00032565999999999997 3.3 0.00032575999999999997 0 0.00032568 0 0.00032578 3.3 0.0003257 3.3 0.0003258 0 0.00032572 0 0.00032582 3.3 0.00032574 3.3 0.00032584 0 0.00032575999999999997 0 0.00032586 3.3 0.00032578 3.3 0.00032588 0 0.0003258 0 0.0003259 3.3 0.00032582 3.3 0.00032592 0 0.00032584 0 0.00032594 3.3 0.00032586 3.3 0.00032596 0 0.00032588 0 0.00032598 3.3 0.0003259 3.3 0.000326 0 0.00032592 0 0.00032602 3.3 0.00032594 3.3 0.00032604 0 0.00032596 0 0.00032606 3.3 0.00032597999999999997 3.3 0.00032607999999999997 0 0.000326 0 0.0003261 3.3 0.00032602 3.3 0.00032612 0 0.00032604 0 0.00032614 3.3 0.00032606 3.3 0.00032616 0 0.00032607999999999997 0 0.00032617999999999997 3.3 0.0003261 3.3 0.0003262 0 0.00032612 0 0.00032622 3.3 0.00032614 3.3 0.00032624 0 0.00032616 0 0.00032626 3.3 0.00032617999999999997 3.3 0.00032627999999999997 0 0.0003262 0 0.0003263 3.3 0.00032622 3.3 0.00032632 0 0.00032624 0 0.00032634 3.3 0.00032626 3.3 0.00032636 0 0.00032627999999999997 0 0.00032638 3.3 0.0003263 3.3 0.0003264 0 0.00032632 0 0.00032642 3.3 0.00032634 3.3 0.00032644 0 0.00032636 0 0.00032646 3.3 0.00032638 3.3 0.00032648 0 0.00032639999999999996 0 0.00032649999999999997 3.3 0.00032642 3.3 0.00032652 0 0.00032644 0 0.00032654 3.3 0.00032646 3.3 0.00032656 0 0.00032648 0 0.00032658 3.3 0.00032649999999999997 3.3 0.00032659999999999997 0 0.00032652 0 0.00032662 3.3 0.00032654 3.3 0.00032664 0 0.00032656 0 0.00032666 3.3 0.00032658 3.3 0.00032668 0 0.00032659999999999997 0 0.00032669999999999997 3.3 0.00032662 3.3 0.00032672 0 0.00032664 0 0.00032674 3.3 0.00032666 3.3 0.00032676 0 0.00032668 0 0.00032678 3.3 0.00032669999999999997 3.3 0.0003268 0 0.00032672 0 0.00032682 3.3 0.00032674 3.3 0.00032684 0 0.00032676 0 0.00032686 3.3 0.00032678 3.3 0.00032688 0 0.0003268 0 0.0003269 3.3 0.00032681999999999996 3.3 0.00032691999999999997 0 0.00032684 0 0.00032694 3.3 0.00032686 3.3 0.00032696 0 0.00032688 0 0.00032698 3.3 0.0003269 3.3 0.000327 0 0.00032691999999999997 0 0.00032701999999999997 3.3 0.00032694 3.3 0.00032704 0 0.00032696 0 0.00032706 3.3 0.00032698 3.3 0.00032708 0 0.000327 0 0.0003271 3.3 0.00032701999999999997 3.3 0.00032711999999999997 0 0.00032704 0 0.00032714 3.3 0.00032706 3.3 0.00032716 0 0.00032708 0 0.00032718 3.3 0.0003271 3.3 0.0003272 0 0.00032711999999999997 0 0.00032722 3.3 0.00032714 3.3 0.00032724 0 0.00032716 0 0.00032726 3.3 0.00032718 3.3 0.00032728 0 0.0003272 0 0.0003273 3.3 0.00032722 3.3 0.00032732 0 0.00032724 0 0.00032734 3.3 0.00032726 3.3 0.00032736 0 0.00032728 0 0.00032738 3.3 0.0003273 3.3 0.0003274 0 0.00032732 0 0.00032742 3.3 0.00032733999999999997 3.3 0.00032743999999999997 0 0.00032736 0 0.00032746 3.3 0.00032738 3.3 0.00032748 0 0.0003274 0 0.0003275 3.3 0.00032742 3.3 0.00032752 0 0.00032743999999999997 0 0.00032753999999999997 3.3 0.00032746 3.3 0.00032756 0 0.00032748 0 0.00032758 3.3 0.0003275 3.3 0.0003276 0 0.00032752 0 0.00032762 3.3 0.00032753999999999997 3.3 0.00032764 0 0.00032756 0 0.00032766 3.3 0.00032758 3.3 0.00032768 0 0.0003276 0 0.0003277 3.3 0.00032762 3.3 0.00032772 0 0.00032764 0 0.00032774 3.3 0.00032766 3.3 0.00032776 0 0.00032768 0 0.00032778 3.3 0.0003277 3.3 0.0003278 0 0.00032772 0 0.00032782 3.3 0.00032774 3.3 0.00032784 0 0.00032775999999999997 0 0.00032785999999999997 3.3 0.00032778 3.3 0.00032788 0 0.0003278 0 0.0003279 3.3 0.00032782 3.3 0.00032792 0 0.00032784 0 0.00032794 3.3 0.00032785999999999997 3.3 0.00032795999999999997 0 0.00032788 0 0.00032798 3.3 0.0003279 3.3 0.000328 0 0.00032792 0 0.00032802 3.3 0.00032794 3.3 0.00032804 0 0.00032795999999999997 0 0.00032805999999999997 3.3 0.00032798 3.3 0.00032808 0 0.000328 0 0.0003281 3.3 0.00032802 3.3 0.00032812 0 0.00032804 0 0.00032814 3.3 0.00032805999999999997 3.3 0.00032816 0 0.00032808 0 0.00032818 3.3 0.0003281 3.3 0.0003282 0 0.00032812 0 0.00032822 3.3 0.00032814 3.3 0.00032824 0 0.00032816 0 0.00032826 3.3 0.00032817999999999996 3.3 0.00032827999999999997 0 0.0003282 0 0.0003283 3.3 0.00032822 3.3 0.00032832 0 0.00032824 0 0.00032834 3.3 0.00032826 3.3 0.00032836 0 0.00032827999999999997 0 0.00032837999999999997 3.3 0.0003283 3.3 0.0003284 0 0.00032832 0 0.00032842 3.3 0.00032834 3.3 0.00032844 0 0.00032836 0 0.00032846 3.3 0.00032837999999999997 3.3 0.00032847999999999997 0 0.0003284 0 0.0003285 3.3 0.00032842 3.3 0.00032852 0 0.00032844 0 0.00032854 3.3 0.00032846 3.3 0.00032856 0 0.00032847999999999997 0 0.00032858 3.3 0.0003285 3.3 0.0003286 0 0.00032852 0 0.00032862 3.3 0.00032854 3.3 0.00032864 0 0.00032856 0 0.00032866 3.3 0.00032858 3.3 0.00032868 0 0.00032859999999999996 0 0.00032869999999999997 3.3 0.00032862 3.3 0.00032872 0 0.00032864 0 0.00032874 3.3 0.00032866 3.3 0.00032876 0 0.00032868 0 0.00032878 3.3 0.00032869999999999997 3.3 0.00032879999999999997 0 0.00032872 0 0.00032882 3.3 0.00032874 3.3 0.00032884 0 0.00032876 0 0.00032886 3.3 0.00032878 3.3 0.00032888 0 0.00032879999999999997 0 0.00032889999999999997 3.3 0.00032882 3.3 0.00032892 0 0.00032884 0 0.00032894 3.3 0.00032886 3.3 0.00032896 0 0.00032888 0 0.00032898 3.3 0.00032889999999999997 3.3 0.000329 0 0.00032892 0 0.00032902 3.3 0.00032894 3.3 0.00032904 0 0.00032896 0 0.00032906 3.3 0.00032898 3.3 0.00032908 0 0.000329 0 0.0003291 3.3 0.00032902 3.3 0.00032912 0 0.00032904 0 0.00032914 3.3 0.00032906 3.3 0.00032916 0 0.00032908 0 0.00032918 3.3 0.0003291 3.3 0.0003292 0 0.00032911999999999997 0 0.00032921999999999997 3.3 0.00032914 3.3 0.00032924 0 0.00032916 0 0.00032926 3.3 0.00032918 3.3 0.00032928 0 0.0003292 0 0.0003293 3.3 0.00032921999999999997 3.3 0.00032931999999999997 0 0.00032924 0 0.00032934 3.3 0.00032926 3.3 0.00032936 0 0.00032928 0 0.00032938 3.3 0.0003293 3.3 0.0003294 0 0.00032931999999999997 0 0.00032942 3.3 0.00032934 3.3 0.00032944 0 0.00032936 0 0.00032946 3.3 0.00032938 3.3 0.00032948 0 0.0003294 0 0.0003295 3.3 0.00032942 3.3 0.00032952 0 0.00032944 0 0.00032954 3.3 0.00032946 3.3 0.00032956 0 0.00032948 0 0.00032958 3.3 0.0003295 3.3 0.0003296 0 0.00032952 0 0.00032962 3.3 0.00032953999999999997 3.3 0.00032963999999999997 0 0.00032956 0 0.00032966 3.3 0.00032958 3.3 0.00032968 0 0.0003296 0 0.0003297 3.3 0.00032962 3.3 0.00032972 0 0.00032963999999999997 0 0.00032973999999999997 3.3 0.00032966 3.3 0.00032976 0 0.00032968 0 0.00032978 3.3 0.0003297 3.3 0.0003298 0 0.00032972 0 0.00032982 3.3 0.00032973999999999997 3.3 0.00032983999999999997 0 0.00032976 0 0.00032986 3.3 0.00032978 3.3 0.00032988 0 0.0003298 0 0.0003299 3.3 0.00032982 3.3 0.00032992 0 0.00032983999999999997 0 0.00032994 3.3 0.00032986 3.3 0.00032996 0 0.00032988 0 0.00032998 3.3 0.0003299 3.3 0.00033 0 0.00032992 0 0.00033002 3.3 0.00032994 3.3 0.00033004 0 0.00032995999999999996 0 0.00033005999999999997 3.3 0.00032998 3.3 0.00033008 0 0.00033 0 0.0003301 3.3 0.00033002 3.3 0.00033012 0 0.00033004 0 0.00033014 3.3 0.00033005999999999997 3.3 0.00033015999999999997 0 0.00033008 0 0.00033018 3.3 0.0003301 3.3 0.0003302 0 0.00033012 0 0.00033022 3.3 0.00033014 3.3 0.00033024 0 0.00033015999999999997 0 0.00033025999999999997 3.3 0.00033018 3.3 0.00033028 0 0.0003302 0 0.0003303 3.3 0.00033022 3.3 0.00033032 0 0.00033024 0 0.00033034 3.3 0.00033025999999999997 3.3 0.00033036 0 0.00033028 0 0.00033038 3.3 0.0003303 3.3 0.0003304 0 0.00033032 0 0.00033042 3.3 0.00033034 3.3 0.00033044 0 0.00033036 0 0.00033046 3.3 0.00033037999999999996 3.3 0.00033047999999999997 0 0.0003304 0 0.0003305 3.3 0.00033042 3.3 0.00033052 0 0.00033044 0 0.00033054 3.3 0.00033046 3.3 0.00033056 0 0.00033047999999999997 0 0.00033057999999999997 3.3 0.0003305 3.3 0.0003306 0 0.00033052 0 0.00033062 3.3 0.00033054 3.3 0.00033064 0 0.00033056 0 0.00033066 3.3 0.00033057999999999997 3.3 0.00033067999999999997 0 0.0003306 0 0.0003307 3.3 0.00033062 3.3 0.00033072 0 0.00033064 0 0.00033074 3.3 0.00033066 3.3 0.00033076 0 0.00033067999999999997 0 0.00033078 3.3 0.0003307 3.3 0.0003308 0 0.00033072 0 0.00033082 3.3 0.00033074 3.3 0.00033084 0 0.00033076 0 0.00033086 3.3 0.00033078 3.3 0.00033088 0 0.0003308 0 0.0003309 3.3 0.00033082 3.3 0.00033092 0 0.00033084 0 0.00033094 3.3 0.00033086 3.3 0.00033096 0 0.00033088 0 0.00033098 3.3 0.00033089999999999997 3.3 0.00033099999999999997 0 0.00033092 0 0.00033102 3.3 0.00033094 3.3 0.00033104 0 0.00033096 0 0.00033106 3.3 0.00033098 3.3 0.00033108 0 0.00033099999999999997 0 0.00033109999999999997 3.3 0.00033102 3.3 0.00033112 0 0.00033104 0 0.00033114 3.3 0.00033106 3.3 0.00033116 0 0.00033108 0 0.00033118 3.3 0.00033109999999999997 3.3 0.0003312 0 0.00033112 0 0.00033122 3.3 0.00033114 3.3 0.00033124 0 0.00033116 0 0.00033126 3.3 0.00033118 3.3 0.00033128 0 0.0003312 0 0.0003313 3.3 0.00033122 3.3 0.00033132 0 0.00033124 0 0.00033134 3.3 0.00033126 3.3 0.00033136 0 0.00033128 0 0.00033138 3.3 0.0003313 3.3 0.0003314 0 0.00033131999999999997 0 0.00033141999999999997 3.3 0.00033134 3.3 0.00033144 0 0.00033136 0 0.00033146 3.3 0.00033138 3.3 0.00033148 0 0.0003314 0 0.0003315 3.3 0.00033141999999999997 3.3 0.00033151999999999997 0 0.00033144 0 0.00033154 3.3 0.00033146 3.3 0.00033156 0 0.00033148 0 0.00033158 3.3 0.0003315 3.3 0.0003316 0 0.00033151999999999997 0 0.00033161999999999997 3.3 0.00033154 3.3 0.00033164 0 0.00033156 0 0.00033166 3.3 0.00033158 3.3 0.00033168 0 0.0003316 0 0.0003317 3.3 0.00033161999999999997 3.3 0.00033172 0 0.00033164 0 0.00033174 3.3 0.00033166 3.3 0.00033176 0 0.00033168 0 0.00033178 3.3 0.0003317 3.3 0.0003318 0 0.00033172 0 0.00033182 3.3 0.00033173999999999996 3.3 0.00033183999999999997 0 0.00033176 0 0.00033186 3.3 0.00033178 3.3 0.00033188 0 0.0003318 0 0.0003319 3.3 0.00033182 3.3 0.00033192 0 0.00033183999999999997 0 0.00033193999999999997 3.3 0.00033186 3.3 0.00033196 0 0.00033188 0 0.00033198 3.3 0.0003319 3.3 0.000332 0 0.00033192 0 0.00033202 3.3 0.00033193999999999997 3.3 0.00033203999999999997 0 0.00033196 0 0.00033206 3.3 0.00033198 3.3 0.00033208 0 0.000332 0 0.0003321 3.3 0.00033202 3.3 0.00033212 0 0.00033203999999999997 0 0.00033214 3.3 0.00033206 3.3 0.00033216 0 0.00033208 0 0.00033218 3.3 0.0003321 3.3 0.0003322 0 0.00033212 0 0.00033222 3.3 0.00033214 3.3 0.00033224 0 0.00033215999999999996 0 0.00033225999999999997 3.3 0.00033218 3.3 0.00033228 0 0.0003322 0 0.0003323 3.3 0.00033222 3.3 0.00033232 0 0.00033224 0 0.00033234 3.3 0.00033225999999999997 3.3 0.00033235999999999997 0 0.00033228 0 0.00033238 3.3 0.0003323 3.3 0.0003324 0 0.00033232 0 0.00033242 3.3 0.00033234 3.3 0.00033244 0 0.00033235999999999997 0 0.00033245999999999997 3.3 0.00033238 3.3 0.00033248 0 0.0003324 0 0.0003325 3.3 0.00033242 3.3 0.00033252 0 0.00033244 0 0.00033254 3.3 0.00033245999999999997 3.3 0.00033256 0 0.00033248 0 0.00033258 3.3 0.0003325 3.3 0.0003326 0 0.00033252 0 0.00033262 3.3 0.00033254 3.3 0.00033264 0 0.00033256 0 0.00033266 3.3 0.00033258 3.3 0.00033268 0 0.0003326 0 0.0003327 3.3 0.00033262 3.3 0.00033272 0 0.00033264 0 0.00033274 3.3 0.00033266 3.3 0.00033276 0 0.00033267999999999997 0 0.00033277999999999997 3.3 0.0003327 3.3 0.0003328 0 0.00033272 0 0.00033282 3.3 0.00033274 3.3 0.00033284 0 0.00033276 0 0.00033286 3.3 0.00033277999999999997 3.3 0.00033287999999999997 0 0.0003328 0 0.0003329 3.3 0.00033282 3.3 0.00033292 0 0.00033284 0 0.00033294 3.3 0.00033286 3.3 0.00033296 0 0.00033287999999999997 0 0.00033298 3.3 0.0003329 3.3 0.000333 0 0.00033292 0 0.00033302 3.3 0.00033294 3.3 0.00033304 0 0.00033296 0 0.00033306 3.3 0.00033298 3.3 0.00033308 0 0.000333 0 0.0003331 3.3 0.00033302 3.3 0.00033312 0 0.00033304 0 0.00033314 3.3 0.00033306 3.3 0.00033316 0 0.00033308 0 0.00033318 3.3 0.00033309999999999997 3.3 0.00033319999999999997 0 0.00033312 0 0.00033322 3.3 0.00033314 3.3 0.00033324 0 0.00033316 0 0.00033326 3.3 0.00033318 3.3 0.00033328 0 0.00033319999999999997 0 0.00033329999999999997 3.3 0.00033322 3.3 0.00033332 0 0.00033324 0 0.00033334 3.3 0.00033326 3.3 0.00033336 0 0.00033328 0 0.00033338 3.3 0.00033329999999999997 3.3 0.00033339999999999997 0 0.00033332 0 0.00033342 3.3 0.00033334 3.3 0.00033344 0 0.00033336 0 0.00033346 3.3 0.00033338 3.3 0.00033348 0 0.00033339999999999997 0 0.0003335 3.3 0.00033342 3.3 0.00033352 0 0.00033344 0 0.00033354 3.3 0.00033346 3.3 0.00033356 0 0.00033348 0 0.00033358 3.3 0.0003335 3.3 0.0003336 0 0.00033351999999999996 0 0.00033361999999999997 3.3 0.00033354 3.3 0.00033364 0 0.00033356 0 0.00033366 3.3 0.00033358 3.3 0.00033368 0 0.0003336 0 0.0003337 3.3 0.00033361999999999997 3.3 0.00033371999999999997 0 0.00033364 0 0.00033374 3.3 0.00033366 3.3 0.00033376 0 0.00033368 0 0.00033378 3.3 0.0003337 3.3 0.0003338 0 0.00033371999999999997 0 0.00033381999999999997 3.3 0.00033374 3.3 0.00033384 0 0.00033376 0 0.00033386 3.3 0.00033378 3.3 0.00033388 0 0.0003338 0 0.0003339 3.3 0.00033381999999999997 3.3 0.00033392 0 0.00033384 0 0.00033394 3.3 0.00033386 3.3 0.00033396 0 0.00033388 0 0.00033398 3.3 0.0003339 3.3 0.000334 0 0.00033392 0 0.00033402 3.3 0.00033393999999999996 3.3 0.00033403999999999997 0 0.00033396 0 0.00033406 3.3 0.00033398 3.3 0.00033408 0 0.000334 0 0.0003341 3.3 0.00033402 3.3 0.00033412 0 0.00033403999999999997 0 0.00033413999999999997 3.3 0.00033406 3.3 0.00033416 0 0.00033408 0 0.00033418 3.3 0.0003341 3.3 0.0003342 0 0.00033412 0 0.00033422 3.3 0.00033413999999999997 3.3 0.00033423999999999997 0 0.00033416 0 0.00033426 3.3 0.00033418 3.3 0.00033428 0 0.0003342 0 0.0003343 3.3 0.00033422 3.3 0.00033432 0 0.00033423999999999997 0 0.00033434 3.3 0.00033426 3.3 0.00033436 0 0.00033428 0 0.00033438 3.3 0.0003343 3.3 0.0003344 0 0.00033432 0 0.00033442 3.3 0.00033434 3.3 0.00033444 0 0.00033436 0 0.00033446 3.3 0.00033438 3.3 0.00033448 0 0.0003344 0 0.0003345 3.3 0.00033442 3.3 0.00033452 0 0.00033444 0 0.00033454 3.3 0.00033445999999999997 3.3 0.00033455999999999997 0 0.00033448 0 0.00033458 3.3 0.0003345 3.3 0.0003346 0 0.00033452 0 0.00033462 3.3 0.00033454 3.3 0.00033464 0 0.00033455999999999997 0 0.00033465999999999997 3.3 0.00033458 3.3 0.00033468 0 0.0003346 0 0.0003347 3.3 0.00033462 3.3 0.00033472 0 0.00033464 0 0.00033474 3.3 0.00033465999999999997 3.3 0.00033476 0 0.00033468 0 0.00033478 3.3 0.0003347 3.3 0.0003348 0 0.00033472 0 0.00033482 3.3 0.00033474 3.3 0.00033484 0 0.00033476 0 0.00033486 3.3 0.00033478 3.3 0.00033488 0 0.0003348 0 0.0003349 3.3 0.00033482 3.3 0.00033492 0 0.00033484 0 0.00033494 3.3 0.00033486 3.3 0.00033496 0 0.00033487999999999997 0 0.00033497999999999997 3.3 0.0003349 3.3 0.000335 0 0.00033492 0 0.00033502 3.3 0.00033494 3.3 0.00033504 0 0.00033496 0 0.00033506 3.3 0.00033497999999999997 3.3 0.00033507999999999997 0 0.000335 0 0.0003351 3.3 0.00033502 3.3 0.00033512 0 0.00033504 0 0.00033514 3.3 0.00033506 3.3 0.00033516 0 0.00033507999999999997 0 0.00033517999999999997 3.3 0.0003351 3.3 0.0003352 0 0.00033512 0 0.00033522 3.3 0.00033514 3.3 0.00033524 0 0.00033516 0 0.00033526 3.3 0.00033517999999999997 3.3 0.00033528 0 0.0003352 0 0.0003353 3.3 0.00033522 3.3 0.00033532 0 0.00033524 0 0.00033534 3.3 0.00033526 3.3 0.00033536 0 0.00033528 0 0.00033538 3.3 0.00033529999999999996 3.3 0.00033539999999999997 0 0.00033532 0 0.00033542 3.3 0.00033534 3.3 0.00033544 0 0.00033536 0 0.00033546 3.3 0.00033538 3.3 0.00033548 0 0.00033539999999999997 0 0.00033549999999999997 3.3 0.00033542 3.3 0.00033552 0 0.00033544 0 0.00033554 3.3 0.00033546 3.3 0.00033556 0 0.00033548 0 0.00033558 3.3 0.00033549999999999997 3.3 0.00033559999999999997 0 0.00033552 0 0.00033562 3.3 0.00033554 3.3 0.00033564 0 0.00033556 0 0.00033566 3.3 0.00033558 3.3 0.00033568 0 0.00033559999999999997 0 0.0003357 3.3 0.00033562 3.3 0.00033572 0 0.00033564 0 0.00033574 3.3 0.00033566 3.3 0.00033576 0 0.00033568 0 0.00033578 3.3 0.0003357 3.3 0.0003358 0 0.00033571999999999996 0 0.00033581999999999997 3.3 0.00033574 3.3 0.00033584 0 0.00033576 0 0.00033586 3.3 0.00033578 3.3 0.00033588 0 0.0003358 0 0.0003359 3.3 0.00033581999999999997 3.3 0.00033591999999999997 0 0.00033584 0 0.00033594 3.3 0.00033586 3.3 0.00033596 0 0.00033588 0 0.00033598 3.3 0.0003359 3.3 0.000336 0 0.00033591999999999997 0 0.00033601999999999997 3.3 0.00033594 3.3 0.00033604 0 0.00033596 0 0.00033606 3.3 0.00033598 3.3 0.00033608 0 0.000336 0 0.0003361 3.3 0.00033601999999999997 3.3 0.00033612 0 0.00033604 0 0.00033614 3.3 0.00033606 3.3 0.00033616 0 0.00033608 0 0.00033618 3.3 0.0003361 3.3 0.0003362 0 0.00033612 0 0.00033622 3.3 0.00033614 3.3 0.00033624 0 0.00033616 0 0.00033626 3.3 0.00033618 3.3 0.00033628 0 0.0003362 0 0.0003363 3.3 0.00033622 3.3 0.00033632 0 0.00033623999999999997 0 0.00033633999999999997 3.3 0.00033626 3.3 0.00033636 0 0.00033628 0 0.00033638 3.3 0.0003363 3.3 0.0003364 0 0.00033632 0 0.00033642 3.3 0.00033633999999999997 3.3 0.00033643999999999997 0 0.00033636 0 0.00033646 3.3 0.00033638 3.3 0.00033648 0 0.0003364 0 0.0003365 3.3 0.00033642 3.3 0.00033652 0 0.00033643999999999997 0 0.00033653999999999997 3.3 0.00033646 3.3 0.00033656 0 0.00033648 0 0.00033658 3.3 0.0003365 3.3 0.0003366 0 0.00033652 0 0.00033662 3.3 0.00033653999999999997 3.3 0.00033664 0 0.00033656 0 0.00033666 3.3 0.00033658 3.3 0.00033668 0 0.0003366 0 0.0003367 3.3 0.00033662 3.3 0.00033672 0 0.00033664 0 0.00033674 3.3 0.00033665999999999996 3.3 0.00033675999999999997 0 0.00033668 0 0.00033678 3.3 0.0003367 3.3 0.0003368 0 0.00033672 0 0.00033682 3.3 0.00033674 3.3 0.00033684 0 0.00033675999999999997 0 0.00033685999999999997 3.3 0.00033678 3.3 0.00033688 0 0.0003368 0 0.0003369 3.3 0.00033682 3.3 0.00033692 0 0.00033684 0 0.00033694 3.3 0.00033685999999999997 3.3 0.00033695999999999997 0 0.00033688 0 0.00033698 3.3 0.0003369 3.3 0.000337 0 0.00033692 0 0.00033702 3.3 0.00033694 3.3 0.00033704 0 0.00033695999999999997 0 0.00033706 3.3 0.00033698 3.3 0.00033708 0 0.000337 0 0.0003371 3.3 0.00033702 3.3 0.00033712 0 0.00033704 0 0.00033714 3.3 0.00033706 3.3 0.00033716 0 0.00033707999999999996 0 0.00033717999999999997 3.3 0.0003371 3.3 0.0003372 0 0.00033712 0 0.00033722 3.3 0.00033714 3.3 0.00033724 0 0.00033716 0 0.00033726 3.3 0.00033717999999999997 3.3 0.00033727999999999997 0 0.0003372 0 0.0003373 3.3 0.00033722 3.3 0.00033732 0 0.00033724 0 0.00033734 3.3 0.00033726 3.3 0.00033736 0 0.00033727999999999997 0 0.00033737999999999997 3.3 0.0003373 3.3 0.0003374 0 0.00033732 0 0.00033742 3.3 0.00033734 3.3 0.00033744 0 0.00033736 0 0.00033746 3.3 0.00033737999999999997 3.3 0.00033748 0 0.0003374 0 0.0003375 3.3 0.00033742 3.3 0.00033752 0 0.00033744 0 0.00033754 3.3 0.00033746 3.3 0.00033756 0 0.00033748 0 0.00033758 3.3 0.0003375 3.3 0.0003376 0 0.00033752 0 0.00033762 3.3 0.00033754 3.3 0.00033764 0 0.00033756 0 0.00033766 3.3 0.00033758 3.3 0.00033768 0 0.00033759999999999997 0 0.00033769999999999997 3.3 0.00033762 3.3 0.00033772 0 0.00033764 0 0.00033774 3.3 0.00033766 3.3 0.00033776 0 0.00033768 0 0.00033778 3.3 0.00033769999999999997 3.3 0.00033779999999999997 0 0.00033772 0 0.00033782 3.3 0.00033774 3.3 0.00033784 0 0.00033776 0 0.00033786 3.3 0.00033778 3.3 0.00033788 0 0.00033779999999999997 0 0.0003379 3.3 0.00033782 3.3 0.00033792 0 0.00033784 0 0.00033794 3.3 0.00033786 3.3 0.00033796 0 0.00033788 0 0.00033798 3.3 0.0003379 3.3 0.000338 0 0.00033792 0 0.00033802 3.3 0.00033794 3.3 0.00033804 0 0.00033796 0 0.00033806 3.3 0.00033798 3.3 0.00033808 0 0.000338 0 0.0003381 3.3 0.00033801999999999997 3.3 0.00033811999999999997 0 0.00033804 0 0.00033814 3.3 0.00033806 3.3 0.00033816 0 0.00033808 0 0.00033818 3.3 0.0003381 3.3 0.0003382 0 0.00033811999999999997 0 0.00033821999999999997 3.3 0.00033814 3.3 0.00033824 0 0.00033816 0 0.00033826 3.3 0.00033818 3.3 0.00033828 0 0.0003382 0 0.0003383 3.3 0.00033821999999999997 3.3 0.00033831999999999997 0 0.00033824 0 0.00033834 3.3 0.00033826 3.3 0.00033836 0 0.00033828 0 0.00033838 3.3 0.0003383 3.3 0.0003384 0 0.00033831999999999997 0 0.00033842 3.3 0.00033834 3.3 0.00033844 0 0.00033836 0 0.00033846 3.3 0.00033838 3.3 0.00033848 0 0.0003384 0 0.0003385 3.3 0.00033842 3.3 0.00033852 0 0.00033843999999999996 0 0.00033853999999999997 3.3 0.00033846 3.3 0.00033856 0 0.00033848 0 0.00033858 3.3 0.0003385 3.3 0.0003386 0 0.00033852 0 0.00033862 3.3 0.00033853999999999997 3.3 0.00033863999999999997 0 0.00033856 0 0.00033866 3.3 0.00033858 3.3 0.00033868 0 0.0003386 0 0.0003387 3.3 0.00033862 3.3 0.00033872 0 0.00033863999999999997 0 0.00033873999999999997 3.3 0.00033866 3.3 0.00033876 0 0.00033868 0 0.00033878 3.3 0.0003387 3.3 0.0003388 0 0.00033872 0 0.00033882 3.3 0.00033873999999999997 3.3 0.00033884 0 0.00033876 0 0.00033886 3.3 0.00033878 3.3 0.00033888 0 0.0003388 0 0.0003389 3.3 0.00033882 3.3 0.00033892 0 0.00033884 0 0.00033894 3.3 0.00033885999999999996 3.3 0.00033895999999999997 0 0.00033888 0 0.00033898 3.3 0.0003389 3.3 0.000339 0 0.00033892 0 0.00033902 3.3 0.00033894 3.3 0.00033904 0 0.00033895999999999997 0 0.00033905999999999997 3.3 0.00033898 3.3 0.00033908 0 0.000339 0 0.0003391 3.3 0.00033902 3.3 0.00033912 0 0.00033904 0 0.00033914 3.3 0.00033905999999999997 3.3 0.00033915999999999997 0 0.00033908 0 0.00033918 3.3 0.0003391 3.3 0.0003392 0 0.00033912 0 0.00033922 3.3 0.00033914 3.3 0.00033924 0 0.00033915999999999997 0 0.00033926 3.3 0.00033918 3.3 0.00033928 0 0.0003392 0 0.0003393 3.3 0.00033922 3.3 0.00033932 0 0.00033924 0 0.00033934 3.3 0.00033926 3.3 0.00033936 0 0.00033928 0 0.00033938 3.3 0.0003393 3.3 0.0003394 0 0.00033932 0 0.00033942 3.3 0.00033934 3.3 0.00033944 0 0.00033936 0 0.00033946 3.3 0.00033937999999999997 3.3 0.00033947999999999997 0 0.0003394 0 0.0003395 3.3 0.00033942 3.3 0.00033952 0 0.00033944 0 0.00033954 3.3 0.00033946 3.3 0.00033956 0 0.00033947999999999997 0 0.00033957999999999997 3.3 0.0003395 3.3 0.0003396 0 0.00033952 0 0.00033962 3.3 0.00033954 3.3 0.00033964 0 0.00033956 0 0.00033966 3.3 0.00033957999999999997 3.3 0.00033968 0 0.0003396 0 0.0003397 3.3 0.00033962 3.3 0.00033972 0 0.00033964 0 0.00033974 3.3 0.00033966 3.3 0.00033976 0 0.00033968 0 0.00033978 3.3 0.0003397 3.3 0.0003398 0 0.00033972 0 0.00033982 3.3 0.00033974 3.3 0.00033984 0 0.00033976 0 0.00033986 3.3 0.00033978 3.3 0.00033988 0 0.00033979999999999997 0 0.00033989999999999997 3.3 0.00033982 3.3 0.00033992 0 0.00033984 0 0.00033994 3.3 0.00033986 3.3 0.00033996 0 0.00033988 0 0.00033998 3.3 0.00033989999999999997 3.3 0.00033999999999999997 0 0.00033992 0 0.00034002 3.3 0.00033994 3.3 0.00034004 0 0.00033996 0 0.00034006 3.3 0.00033998 3.3 0.00034008 0 0.00033999999999999997 0 0.00034009999999999997 3.3 0.00034002 3.3 0.00034012 0 0.00034004 0 0.00034014 3.3 0.00034006 3.3 0.00034016 0 0.00034008 0 0.00034018 3.3 0.00034009999999999997 3.3 0.0003402 0 0.00034012 0 0.00034022 3.3 0.00034014 3.3 0.00034024 0 0.00034016 0 0.00034026 3.3 0.00034018 3.3 0.00034028 0 0.0003402 0 0.0003403 3.3 0.00034021999999999996 3.3 0.00034031999999999997 0 0.00034024 0 0.00034034 3.3 0.00034026 3.3 0.00034036 0 0.00034028 0 0.00034038 3.3 0.0003403 3.3 0.0003404 0 0.00034031999999999997 0 0.00034041999999999997 3.3 0.00034034 3.3 0.00034044 0 0.00034036 0 0.00034046 3.3 0.00034038 3.3 0.00034048 0 0.0003404 0 0.0003405 3.3 0.00034041999999999997 3.3 0.00034051999999999997 0 0.00034044 0 0.00034054 3.3 0.00034046 3.3 0.00034056 0 0.00034048 0 0.00034058 3.3 0.0003405 3.3 0.0003406 0 0.00034051999999999997 0 0.00034062 3.3 0.00034054 3.3 0.00034064 0 0.00034056 0 0.00034066 3.3 0.00034058 3.3 0.00034068 0 0.0003406 0 0.0003407 3.3 0.00034062 3.3 0.00034072 0 0.00034063999999999996 0 0.00034073999999999997 3.3 0.00034066 3.3 0.00034076 0 0.00034068 0 0.00034078 3.3 0.0003407 3.3 0.0003408 0 0.00034072 0 0.00034082 3.3 0.00034073999999999997 3.3 0.00034083999999999997 0 0.00034076 0 0.00034086 3.3 0.00034078 3.3 0.00034088 0 0.0003408 0 0.0003409 3.3 0.00034082 3.3 0.00034092 0 0.00034083999999999997 0 0.00034093999999999997 3.3 0.00034086 3.3 0.00034096 0 0.00034088 0 0.00034098 3.3 0.0003409 3.3 0.000341 0 0.00034092 0 0.00034102 3.3 0.00034093999999999997 3.3 0.00034104 0 0.00034096 0 0.00034106 3.3 0.00034098 3.3 0.00034108 0 0.000341 0 0.0003411 3.3 0.00034102 3.3 0.00034112 0 0.00034104 0 0.00034114 3.3 0.00034106 3.3 0.00034116 0 0.00034108 0 0.00034118 3.3 0.0003411 3.3 0.0003412 0 0.00034112 0 0.00034122 3.3 0.00034114 3.3 0.00034124 0 0.00034115999999999997 0 0.00034125999999999997 3.3 0.00034118 3.3 0.00034128 0 0.0003412 0 0.0003413 3.3 0.00034122 3.3 0.00034132 0 0.00034124 0 0.00034134 3.3 0.00034125999999999997 3.3 0.00034135999999999997 0 0.00034128 0 0.00034138 3.3 0.0003413 3.3 0.0003414 0 0.00034132 0 0.00034142 3.3 0.00034134 3.3 0.00034144 0 0.00034135999999999997 0 0.00034146 3.3 0.00034138 3.3 0.00034148 0 0.0003414 0 0.0003415 3.3 0.00034142 3.3 0.00034152 0 0.00034144 0 0.00034154 3.3 0.00034146 3.3 0.00034156 0 0.00034148 0 0.00034158 3.3 0.0003415 3.3 0.0003416 0 0.00034152 0 0.00034162 3.3 0.00034154 3.3 0.00034164 0 0.00034156 0 0.00034166 3.3 0.00034157999999999997 3.3 0.00034167999999999997 0 0.0003416 0 0.0003417 3.3 0.00034162 3.3 0.00034172 0 0.00034164 0 0.00034174 3.3 0.00034166 3.3 0.00034176 0 0.00034167999999999997 0 0.00034177999999999997 3.3 0.0003417 3.3 0.0003418 0 0.00034172 0 0.00034182 3.3 0.00034174 3.3 0.00034184 0 0.00034176 0 0.00034186 3.3 0.00034177999999999997 3.3 0.00034187999999999997 0 0.0003418 0 0.0003419 3.3 0.00034182 3.3 0.00034192 0 0.00034184 0 0.00034194 3.3 0.00034186 3.3 0.00034196 0 0.00034187999999999997 0 0.00034198 3.3 0.0003419 3.3 0.000342 0 0.00034192 0 0.00034202 3.3 0.00034194 3.3 0.00034204 0 0.00034196 0 0.00034206 3.3 0.00034198 3.3 0.00034208 0 0.00034199999999999996 0 0.00034209999999999997 3.3 0.00034202 3.3 0.00034212 0 0.00034204 0 0.00034214 3.3 0.00034206 3.3 0.00034216 0 0.00034208 0 0.00034218 3.3 0.00034209999999999997 3.3 0.00034219999999999997 0 0.00034212 0 0.00034222 3.3 0.00034214 3.3 0.00034224 0 0.00034216 0 0.00034226 3.3 0.00034218 3.3 0.00034228 0 0.00034219999999999997 0 0.00034229999999999997 3.3 0.00034222 3.3 0.00034232 0 0.00034224 0 0.00034234 3.3 0.00034226 3.3 0.00034236 0 0.00034228 0 0.00034238 3.3 0.00034229999999999997 3.3 0.0003424 0 0.00034232 0 0.00034242 3.3 0.00034234 3.3 0.00034244 0 0.00034236 0 0.00034246 3.3 0.00034238 3.3 0.00034248 0 0.0003424 0 0.0003425 3.3 0.00034241999999999996 3.3 0.00034251999999999997 0 0.00034244 0 0.00034254 3.3 0.00034246 3.3 0.00034256 0 0.00034248 0 0.00034258 3.3 0.0003425 3.3 0.0003426 0 0.00034251999999999997 0 0.00034261999999999997 3.3 0.00034254 3.3 0.00034264 0 0.00034256 0 0.00034266 3.3 0.00034258 3.3 0.00034268 0 0.0003426 0 0.0003427 3.3 0.00034261999999999997 3.3 0.00034271999999999997 0 0.00034264 0 0.00034274 3.3 0.00034266 3.3 0.00034276 0 0.00034268 0 0.00034278 3.3 0.0003427 3.3 0.0003428 0 0.00034271999999999997 0 0.00034282 3.3 0.00034274 3.3 0.00034284 0 0.00034276 0 0.00034286 3.3 0.00034278 3.3 0.00034288 0 0.0003428 0 0.0003429 3.3 0.00034282 3.3 0.00034292 0 0.00034284 0 0.00034294 3.3 0.00034286 3.3 0.00034296 0 0.00034288 0 0.00034298 3.3 0.0003429 3.3 0.000343 0 0.00034292 0 0.00034302 3.3 0.00034293999999999997 3.3 0.00034303999999999997 0 0.00034296 0 0.00034306 3.3 0.00034298 3.3 0.00034308 0 0.000343 0 0.0003431 3.3 0.00034302 3.3 0.00034312 0 0.00034303999999999997 0 0.00034313999999999997 3.3 0.00034306 3.3 0.00034316 0 0.00034308 0 0.00034318 3.3 0.0003431 3.3 0.0003432 0 0.00034312 0 0.00034322 3.3 0.00034313999999999997 3.3 0.00034324 0 0.00034316 0 0.00034326 3.3 0.00034318 3.3 0.00034328 0 0.0003432 0 0.0003433 3.3 0.00034322 3.3 0.00034332 0 0.00034324 0 0.00034334 3.3 0.00034326 3.3 0.00034336 0 0.00034328 0 0.00034338 3.3 0.0003433 3.3 0.0003434 0 0.00034332 0 0.00034342 3.3 0.00034334 3.3 0.00034344 0 0.00034335999999999997 0 0.00034345999999999997 3.3 0.00034338 3.3 0.00034348 0 0.0003434 0 0.0003435 3.3 0.00034342 3.3 0.00034352 0 0.00034344 0 0.00034354 3.3 0.00034345999999999997 3.3 0.00034355999999999997 0 0.00034348 0 0.00034358 3.3 0.0003435 3.3 0.0003436 0 0.00034352 0 0.00034362 3.3 0.00034354 3.3 0.00034364 0 0.00034355999999999997 0 0.00034365999999999997 3.3 0.00034358 3.3 0.00034368 0 0.0003436 0 0.0003437 3.3 0.00034362 3.3 0.00034372 0 0.00034364 0 0.00034374 3.3 0.00034365999999999997 3.3 0.00034376 0 0.00034368 0 0.00034378 3.3 0.0003437 3.3 0.0003438 0 0.00034372 0 0.00034382 3.3 0.00034374 3.3 0.00034384 0 0.00034376 0 0.00034386 3.3 0.00034377999999999996 3.3 0.00034387999999999997 0 0.0003438 0 0.0003439 3.3 0.00034382 3.3 0.00034392 0 0.00034384 0 0.00034394 3.3 0.00034386 3.3 0.00034396 0 0.00034387999999999997 0 0.00034397999999999997 3.3 0.0003439 3.3 0.000344 0 0.00034392 0 0.00034402 3.3 0.00034394 3.3 0.00034404 0 0.00034396 0 0.00034406 3.3 0.00034397999999999997 3.3 0.00034407999999999997 0 0.000344 0 0.0003441 3.3 0.00034402 3.3 0.00034412 0 0.00034404 0 0.00034414 3.3 0.00034406 3.3 0.00034416 0 0.00034407999999999997 0 0.00034418 3.3 0.0003441 3.3 0.0003442 0 0.00034412 0 0.00034422 3.3 0.00034414 3.3 0.00034424 0 0.00034416 0 0.00034426 3.3 0.00034418 3.3 0.00034428 0 0.00034419999999999996 0 0.00034429999999999997 3.3 0.00034422 3.3 0.00034432 0 0.00034424 0 0.00034434 3.3 0.00034426 3.3 0.00034436 0 0.00034428 0 0.00034438 3.3 0.00034429999999999997 3.3 0.00034439999999999997 0 0.00034432 0 0.00034442 3.3 0.00034434 3.3 0.00034444 0 0.00034436 0 0.00034446 3.3 0.00034438 3.3 0.00034448 0 0.00034439999999999997 0 0.00034449999999999997 3.3 0.00034442 3.3 0.00034452 0 0.00034444 0 0.00034454 3.3 0.00034446 3.3 0.00034456 0 0.00034448 0 0.00034458 3.3 0.00034449999999999997 3.3 0.0003446 0 0.00034452 0 0.00034462 3.3 0.00034454 3.3 0.00034464 0 0.00034456 0 0.00034466 3.3 0.00034458 3.3 0.00034468 0 0.0003446 0 0.0003447 3.3 0.00034462 3.3 0.00034472 0 0.00034464 0 0.00034474 3.3 0.00034466 3.3 0.00034476 0 0.00034468 0 0.00034478 3.3 0.0003447 3.3 0.0003448 0 0.00034471999999999997 0 0.00034481999999999997 3.3 0.00034474 3.3 0.00034484 0 0.00034476 0 0.00034486 3.3 0.00034478 3.3 0.00034488 0 0.0003448 0 0.0003449 3.3 0.00034481999999999997 3.3 0.00034491999999999997 0 0.00034484 0 0.00034494 3.3 0.00034486 3.3 0.00034496 0 0.00034488 0 0.00034498 3.3 0.0003449 3.3 0.000345 0 0.00034491999999999997 0 0.00034502 3.3 0.00034494 3.3 0.00034504 0 0.00034496 0 0.00034506 3.3 0.00034498 3.3 0.00034508 0 0.000345 0 0.0003451 3.3 0.00034502 3.3 0.00034512 0 0.00034504 0 0.00034514 3.3 0.00034506 3.3 0.00034516 0 0.00034508 0 0.00034518 3.3 0.0003451 3.3 0.0003452 0 0.00034512 0 0.00034522 3.3 0.00034513999999999997 3.3 0.00034523999999999997 0 0.00034516 0 0.00034526 3.3 0.00034518 3.3 0.00034528 0 0.0003452 0 0.0003453 3.3 0.00034522 3.3 0.00034532 0 0.00034523999999999997 0 0.00034533999999999997 3.3 0.00034526 3.3 0.00034536 0 0.00034528 0 0.00034538 3.3 0.0003453 3.3 0.0003454 0 0.00034532 0 0.00034542 3.3 0.00034533999999999997 3.3 0.00034543999999999997 0 0.00034536 0 0.00034546 3.3 0.00034538 3.3 0.00034548 0 0.0003454 0 0.0003455 3.3 0.00034542 3.3 0.00034552 0 0.00034543999999999997 0 0.00034554 3.3 0.00034546 3.3 0.00034556 0 0.00034548 0 0.00034558 3.3 0.0003455 3.3 0.0003456 0 0.00034552 0 0.00034562 3.3 0.00034554 3.3 0.00034564 0 0.00034555999999999996 0 0.00034565999999999997 3.3 0.00034558 3.3 0.00034568 0 0.0003456 0 0.0003457 3.3 0.00034562 3.3 0.00034572 0 0.00034564 0 0.00034574 3.3 0.00034565999999999997 3.3 0.00034575999999999997 0 0.00034568 0 0.00034578 3.3 0.0003457 3.3 0.0003458 0 0.00034572 0 0.00034582 3.3 0.00034574 3.3 0.00034584 0 0.00034575999999999997 0 0.00034585999999999997 3.3 0.00034578 3.3 0.00034588 0 0.0003458 0 0.0003459 3.3 0.00034582 3.3 0.00034592 0 0.00034584 0 0.00034594 3.3 0.00034585999999999997 3.3 0.00034596 0 0.00034588 0 0.00034598 3.3 0.0003459 3.3 0.000346 0 0.00034592 0 0.00034602 3.3 0.00034594 3.3 0.00034604 0 0.00034596 0 0.00034606 3.3 0.00034597999999999996 3.3 0.00034607999999999997 0 0.000346 0 0.0003461 3.3 0.00034602 3.3 0.00034612 0 0.00034604 0 0.00034614 3.3 0.00034606 3.3 0.00034616 0 0.00034607999999999997 0 0.00034617999999999997 3.3 0.0003461 3.3 0.0003462 0 0.00034612 0 0.00034622 3.3 0.00034614 3.3 0.00034624 0 0.00034616 0 0.00034626 3.3 0.00034617999999999997 3.3 0.00034627999999999997 0 0.0003462 0 0.0003463 3.3 0.00034622 3.3 0.00034632 0 0.00034624 0 0.00034634 3.3 0.00034626 3.3 0.00034636 0 0.00034627999999999997 0 0.00034638 3.3 0.0003463 3.3 0.0003464 0 0.00034632 0 0.00034642 3.3 0.00034634 3.3 0.00034644 0 0.00034636 0 0.00034646 3.3 0.00034638 3.3 0.00034648 0 0.0003464 0 0.0003465 3.3 0.00034642 3.3 0.00034652 0 0.00034644 0 0.00034654 3.3 0.00034646 3.3 0.00034656 0 0.00034648 0 0.00034658 3.3 0.00034649999999999997 3.3 0.00034659999999999997 0 0.00034652 0 0.00034662 3.3 0.00034654 3.3 0.00034664 0 0.00034656 0 0.00034666 3.3 0.00034658 3.3 0.00034668 0 0.00034659999999999997 0 0.00034669999999999997 3.3 0.00034662 3.3 0.00034672 0 0.00034664 0 0.00034674 3.3 0.00034666 3.3 0.00034676 0 0.00034668 0 0.00034678 3.3 0.00034669999999999997 3.3 0.00034679999999999997 0 0.00034672 0 0.00034682 3.3 0.00034674 3.3 0.00034684 0 0.00034676 0 0.00034686 3.3 0.00034678 3.3 0.00034688 0 0.00034679999999999997 0 0.0003469 3.3 0.00034682 3.3 0.00034692 0 0.00034684 0 0.00034694 3.3 0.00034686 3.3 0.00034696 0 0.00034688 0 0.00034698 3.3 0.0003469 3.3 0.000347 0 0.00034691999999999996 0 0.00034701999999999997 3.3 0.00034694 3.3 0.00034704 0 0.00034696 0 0.00034706 3.3 0.00034698 3.3 0.00034708 0 0.000347 0 0.0003471 3.3 0.00034701999999999997 3.3 0.00034711999999999997 0 0.00034704 0 0.00034714 3.3 0.00034706 3.3 0.00034716 0 0.00034708 0 0.00034718 3.3 0.0003471 3.3 0.0003472 0 0.00034711999999999997 0 0.00034721999999999997 3.3 0.00034714 3.3 0.00034724 0 0.00034716 0 0.00034726 3.3 0.00034718 3.3 0.00034728 0 0.0003472 0 0.0003473 3.3 0.00034721999999999997 3.3 0.00034732 0 0.00034724 0 0.00034734 3.3 0.00034726 3.3 0.00034736 0 0.00034728 0 0.00034738 3.3 0.0003473 3.3 0.0003474 0 0.00034732 0 0.00034742 3.3 0.00034733999999999996 3.3 0.00034743999999999997 0 0.00034736 0 0.00034746 3.3 0.00034738 3.3 0.00034748 0 0.0003474 0 0.0003475 3.3 0.00034742 3.3 0.00034752 0 0.00034743999999999997 0 0.00034753999999999997 3.3 0.00034746 3.3 0.00034756 0 0.00034748 0 0.00034758 3.3 0.0003475 3.3 0.0003476 0 0.00034752 0 0.00034762 3.3 0.00034753999999999997 3.3 0.00034763999999999997 0 0.00034756 0 0.00034766 3.3 0.00034758 3.3 0.00034768 0 0.0003476 0 0.0003477 3.3 0.00034762 3.3 0.00034772 0 0.00034763999999999997 0 0.00034774 3.3 0.00034766 3.3 0.00034776 0 0.00034768 0 0.00034778 3.3 0.0003477 3.3 0.0003478 0 0.00034772 0 0.00034782 3.3 0.00034774 3.3 0.00034784 0 0.00034775999999999996 0 0.00034785999999999997 3.3 0.00034778 3.3 0.00034788 0 0.0003478 0 0.0003479 3.3 0.00034782 3.3 0.00034792 0 0.00034784 0 0.00034794 3.3 0.00034785999999999997 3.3 0.00034795999999999997 0 0.00034788 0 0.00034798 3.3 0.0003479 3.3 0.000348 0 0.00034792 0 0.00034802 3.3 0.00034794 3.3 0.00034804 0 0.00034795999999999997 0 0.00034805999999999997 3.3 0.00034798 3.3 0.00034808 0 0.000348 0 0.0003481 3.3 0.00034802 3.3 0.00034812 0 0.00034804 0 0.00034814 3.3 0.00034805999999999997 3.3 0.00034816 0 0.00034808 0 0.00034818 3.3 0.0003481 3.3 0.0003482 0 0.00034812 0 0.00034822 3.3 0.00034814 3.3 0.00034824 0 0.00034816 0 0.00034826 3.3 0.00034818 3.3 0.00034828 0 0.0003482 0 0.0003483 3.3 0.00034822 3.3 0.00034832 0 0.00034824 0 0.00034834 3.3 0.00034826 3.3 0.00034836 0 0.00034827999999999997 0 0.00034837999999999997 3.3 0.0003483 3.3 0.0003484 0 0.00034832 0 0.00034842 3.3 0.00034834 3.3 0.00034844 0 0.00034836 0 0.00034846 3.3 0.00034837999999999997 3.3 0.00034847999999999997 0 0.0003484 0 0.0003485 3.3 0.00034842 3.3 0.00034852 0 0.00034844 0 0.00034854 3.3 0.00034846 3.3 0.00034856 0 0.00034847999999999997 0 0.00034857999999999997 3.3 0.0003485 3.3 0.0003486 0 0.00034852 0 0.00034862 3.3 0.00034854 3.3 0.00034864 0 0.00034856 0 0.00034866 3.3 0.00034857999999999997 3.3 0.00034868 0 0.0003486 0 0.0003487 3.3 0.00034862 3.3 0.00034872 0 0.00034864 0 0.00034874 3.3 0.00034866 3.3 0.00034876 0 0.00034868 0 0.00034878 3.3 0.00034869999999999996 3.3 0.00034879999999999997 0 0.00034872 0 0.00034882 3.3 0.00034874 3.3 0.00034884 0 0.00034876 0 0.00034886 3.3 0.00034878 3.3 0.00034888 0 0.00034879999999999997 0 0.00034889999999999997 3.3 0.00034882 3.3 0.00034892 0 0.00034884 0 0.00034894 3.3 0.00034886 3.3 0.00034896 0 0.00034888 0 0.00034898 3.3 0.00034889999999999997 3.3 0.00034899999999999997 0 0.00034892 0 0.00034902 3.3 0.00034894 3.3 0.00034904 0 0.00034896 0 0.00034906 3.3 0.00034898 3.3 0.00034908 0 0.00034899999999999997 0 0.0003491 3.3 0.00034902 3.3 0.00034912 0 0.00034904 0 0.00034914 3.3 0.00034906 3.3 0.00034916 0 0.00034908 0 0.00034918 3.3 0.0003491 3.3 0.0003492 0 0.00034911999999999996 0 0.00034921999999999997 3.3 0.00034914 3.3 0.00034924 0 0.00034916 0 0.00034926 3.3 0.00034918 3.3 0.00034928 0 0.0003492 0 0.0003493 3.3 0.00034921999999999997 3.3 0.00034931999999999997 0 0.00034924 0 0.00034934 3.3 0.00034926 3.3 0.00034936 0 0.00034928 0 0.00034938 3.3 0.0003493 3.3 0.0003494 0 0.00034931999999999997 0 0.00034941999999999997 3.3 0.00034934 3.3 0.00034944 0 0.00034936 0 0.00034946 3.3 0.00034938 3.3 0.00034948 0 0.0003494 0 0.0003495 3.3 0.00034941999999999997 3.3 0.00034952 0 0.00034944 0 0.00034954 3.3 0.00034946 3.3 0.00034956 0 0.00034948 0 0.00034958 3.3 0.0003495 3.3 0.0003496 0 0.00034952 0 0.00034962 3.3 0.00034953999999999996 3.3 0.00034963999999999997 0 0.00034956 0 0.00034966 3.3 0.00034958 3.3 0.00034968 0 0.0003496 0 0.0003497 3.3 0.00034962 3.3 0.00034972 0 0.00034963999999999997 0 0.00034973999999999997 3.3 0.00034966 3.3 0.00034976 0 0.00034968 0 0.00034978 3.3 0.0003497 3.3 0.0003498 0 0.00034972 0 0.00034982 3.3 0.00034973999999999997 3.3 0.00034983999999999997 0 0.00034976 0 0.00034986 3.3 0.00034978 3.3 0.00034988 0 0.0003498 0 0.0003499 3.3 0.00034982 3.3 0.00034992 0 0.00034983999999999997 0 0.00034994 3.3 0.00034986 3.3 0.00034996 0 0.00034988 0 0.00034998 3.3 0.0003499 3.3 0.00035 0 0.00034992 0 0.00035002 3.3 0.00034994 3.3 0.00035004 0 0.00034996 0 0.00035006 3.3 0.00034998 3.3 0.00035008 0 0.00035 0 0.0003501 3.3 0.00035002 3.3 0.00035012 0 0.00035004 0 0.00035014 3.3 0.00035005999999999997 3.3 0.00035015999999999997 0 0.00035008 0 0.00035018 3.3 0.0003501 3.3 0.0003502 0 0.00035012 0 0.00035022 3.3 0.00035014 3.3 0.00035024 0 0.00035015999999999997 0 0.00035025999999999997 3.3 0.00035018 3.3 0.00035028 0 0.0003502 0 0.0003503 3.3 0.00035022 3.3 0.00035032 0 0.00035024 0 0.00035034 3.3 0.00035025999999999997 3.3 0.00035035999999999997 0 0.00035028 0 0.00035038 3.3 0.0003503 3.3 0.0003504 0 0.00035032 0 0.00035042 3.3 0.00035034 3.3 0.00035044 0 0.00035035999999999997 0 0.00035046 3.3 0.00035038 3.3 0.00035048 0 0.0003504 0 0.0003505 3.3 0.00035042 3.3 0.00035052 0 0.00035044 0 0.00035054 3.3 0.00035046 3.3 0.00035056 0 0.00035047999999999996 0 0.00035057999999999997 3.3 0.0003505 3.3 0.0003506 0 0.00035052 0 0.00035062 3.3 0.00035054 3.3 0.00035064 0 0.00035056 0 0.00035066 3.3 0.00035057999999999997 3.3 0.00035067999999999997 0 0.0003506 0 0.0003507 3.3 0.00035062 3.3 0.00035072 0 0.00035064 0 0.00035074 3.3 0.00035066 3.3 0.00035076 0 0.00035067999999999997 0 0.00035077999999999997 3.3 0.0003507 3.3 0.0003508 0 0.00035072 0 0.00035082 3.3 0.00035074 3.3 0.00035084 0 0.00035076 0 0.00035086 3.3 0.00035077999999999997 3.3 0.00035088 0 0.0003508 0 0.0003509 3.3 0.00035082 3.3 0.00035092 0 0.00035084 0 0.00035094 3.3 0.00035086 3.3 0.00035096 0 0.00035088 0 0.00035098 3.3 0.00035089999999999996 3.3 0.00035099999999999997 0 0.00035092 0 0.00035102 3.3 0.00035094 3.3 0.00035104 0 0.00035096 0 0.00035106 3.3 0.00035098 3.3 0.00035108 0 0.00035099999999999997 0 0.00035109999999999997 3.3 0.00035102 3.3 0.00035112 0 0.00035104 0 0.00035114 3.3 0.00035106 3.3 0.00035116 0 0.00035108 0 0.00035118 3.3 0.00035109999999999997 3.3 0.00035119999999999997 0 0.00035112 0 0.00035122 3.3 0.00035114 3.3 0.00035124 0 0.00035116 0 0.00035126 3.3 0.00035118 3.3 0.00035128 0 0.00035119999999999997 0 0.0003513 3.3 0.00035122 3.3 0.00035132 0 0.00035124 0 0.00035134 3.3 0.00035126 3.3 0.00035136 0 0.00035128 0 0.00035138 3.3 0.0003513 3.3 0.0003514 0 0.00035131999999999996 0 0.00035141999999999997 3.3 0.00035134 3.3 0.00035144 0 0.00035136 0 0.00035146 3.3 0.00035138 3.3 0.00035148 0 0.0003514 0 0.0003515 3.3 0.00035141999999999997 3.3 0.00035151999999999997 0 0.00035144 0 0.00035154 3.3 0.00035146 3.3 0.00035156 0 0.00035148 0 0.00035158 3.3 0.0003515 3.3 0.0003516 0 0.00035151999999999997 0 0.00035161999999999997 3.3 0.00035154 3.3 0.00035164 0 0.00035156 0 0.00035166 3.3 0.00035158 3.3 0.00035168 0 0.0003516 0 0.0003517 3.3 0.00035161999999999997 3.3 0.00035172 0 0.00035164 0 0.00035174 3.3 0.00035166 3.3 0.00035176 0 0.00035168 0 0.00035178 3.3 0.0003517 3.3 0.0003518 0 0.00035172 0 0.00035182 3.3 0.00035174 3.3 0.00035184 0 0.00035176 0 0.00035186 3.3 0.00035178 3.3 0.00035188 0 0.0003518 0 0.0003519 3.3 0.00035182 3.3 0.00035192 0 0.00035183999999999997 0 0.00035193999999999997 3.3 0.00035186 3.3 0.00035196 0 0.00035188 0 0.00035198 3.3 0.0003519 3.3 0.000352 0 0.00035192 0 0.00035202 3.3 0.00035193999999999997 3.3 0.00035203999999999997 0 0.00035196 0 0.00035206 3.3 0.00035198 3.3 0.00035208 0 0.000352 0 0.0003521 3.3 0.00035202 3.3 0.00035212 0 0.00035203999999999997 0 0.00035213999999999997 3.3 0.00035206 3.3 0.00035216 0 0.00035208 0 0.00035218 3.3 0.0003521 3.3 0.0003522 0 0.00035212 0 0.00035222 3.3 0.00035213999999999997 3.3 0.00035224 0 0.00035216 0 0.00035226 3.3 0.00035218 3.3 0.00035228 0 0.0003522 0 0.0003523 3.3 0.00035222 3.3 0.00035232 0 0.00035224 0 0.00035234 3.3 0.00035225999999999996 3.3 0.00035235999999999997 0 0.00035228 0 0.00035238 3.3 0.0003523 3.3 0.0003524 0 0.00035232 0 0.00035242 3.3 0.00035234 3.3 0.00035244 0 0.00035235999999999997 0 0.00035245999999999997 3.3 0.00035238 3.3 0.00035248 0 0.0003524 0 0.0003525 3.3 0.00035242 3.3 0.00035252 0 0.00035244 0 0.00035254 3.3 0.00035245999999999997 3.3 0.00035255999999999997 0 0.00035248 0 0.00035258 3.3 0.0003525 3.3 0.0003526 0 0.00035252 0 0.00035262 3.3 0.00035254 3.3 0.00035264 0 0.00035255999999999997 0 0.00035266 3.3 0.00035258 3.3 0.00035268 0 0.0003526 0 0.0003527 3.3 0.00035262 3.3 0.00035272 0 0.00035264 0 0.00035274 3.3 0.00035266 3.3 0.00035276 0 0.00035267999999999996 0 0.00035277999999999997 3.3 0.0003527 3.3 0.0003528 0 0.00035272 0 0.00035282 3.3 0.00035274 3.3 0.00035284 0 0.00035276 0 0.00035286 3.3 0.00035277999999999997 3.3 0.00035287999999999997 0 0.0003528 0 0.0003529 3.3 0.00035282 3.3 0.00035292 0 0.00035284 0 0.00035294 3.3 0.00035286 3.3 0.00035296 0 0.00035287999999999997 0 0.00035297999999999997 3.3 0.0003529 3.3 0.000353 0 0.00035292 0 0.00035302 3.3 0.00035294 3.3 0.00035304 0 0.00035296 0 0.00035306 3.3 0.00035297999999999997 3.3 0.00035308 0 0.000353 0 0.0003531 3.3 0.00035302 3.3 0.00035312 0 0.00035304 0 0.00035314 3.3 0.00035306 3.3 0.00035316 0 0.00035308 0 0.00035318 3.3 0.00035309999999999996 3.3 0.00035319999999999997 0 0.00035312 0 0.00035322 3.3 0.00035314 3.3 0.00035324 0 0.00035316 0 0.00035326 3.3 0.00035318 3.3 0.00035328 0 0.00035319999999999997 0 0.00035329999999999997 3.3 0.00035322 3.3 0.00035332 0 0.00035324 0 0.00035334 3.3 0.00035326 3.3 0.00035336 0 0.00035328 0 0.00035338 3.3 0.00035329999999999997 3.3 0.00035339999999999997 0 0.00035332 0 0.00035342 3.3 0.00035334 3.3 0.00035344 0 0.00035336 0 0.00035346 3.3 0.00035338 3.3 0.00035348 0 0.00035339999999999997 0 0.0003535 3.3 0.00035342 3.3 0.00035352 0 0.00035344 0 0.00035354 3.3 0.00035346 3.3 0.00035356 0 0.00035348 0 0.00035358 3.3 0.0003535 3.3 0.0003536 0 0.00035352 0 0.00035362 3.3 0.00035354 3.3 0.00035364 0 0.00035356 0 0.00035366 3.3 0.00035358 3.3 0.00035368 0 0.0003536 0 0.0003537 3.3 0.00035361999999999997 3.3 0.00035371999999999997 0 0.00035364 0 0.00035374 3.3 0.00035366 3.3 0.00035376 0 0.00035368 0 0.00035378 3.3 0.0003537 3.3 0.0003538 0 0.00035371999999999997 0 0.00035381999999999997 3.3 0.00035374 3.3 0.00035384 0 0.00035376 0 0.00035386 3.3 0.00035378 3.3 0.00035388 0 0.0003538 0 0.0003539 3.3 0.00035381999999999997 3.3 0.00035391999999999997 0 0.00035384 0 0.00035394 3.3 0.00035386 3.3 0.00035396 0 0.00035388 0 0.00035398 3.3 0.0003539 3.3 0.000354 0 0.00035391999999999997 0 0.00035402 3.3 0.00035394 3.3 0.00035404 0 0.00035396 0 0.00035406 3.3 0.00035398 3.3 0.00035408 0 0.000354 0 0.0003541 3.3 0.00035402 3.3 0.00035412 0 0.00035403999999999996 0 0.00035413999999999997 3.3 0.00035406 3.3 0.00035416 0 0.00035408 0 0.00035418 3.3 0.0003541 3.3 0.0003542 0 0.00035412 0 0.00035422 3.3 0.00035413999999999997 3.3 0.00035423999999999997 0 0.00035416 0 0.00035426 3.3 0.00035418 3.3 0.00035428 0 0.0003542 0 0.0003543 3.3 0.00035422 3.3 0.00035432 0 0.00035423999999999997 0 0.00035433999999999997 3.3 0.00035426 3.3 0.00035436 0 0.00035428 0 0.00035438 3.3 0.0003543 3.3 0.0003544 0 0.00035432 0 0.00035442 3.3 0.00035433999999999997 3.3 0.00035444 0 0.00035436 0 0.00035446 3.3 0.00035438 3.3 0.00035448 0 0.0003544 0 0.0003545 3.3 0.00035442 3.3 0.00035452 0 0.00035444 0 0.00035454 3.3 0.00035445999999999996 3.3 0.00035455999999999997 0 0.00035448 0 0.00035458 3.3 0.0003545 3.3 0.0003546 0 0.00035452 0 0.00035462 3.3 0.00035454 3.3 0.00035464 0 0.00035455999999999997 0 0.00035465999999999997 3.3 0.00035458 3.3 0.00035468 0 0.0003546 0 0.0003547 3.3 0.00035462 3.3 0.00035472 0 0.00035464 0 0.00035474 3.3 0.00035465999999999997 3.3 0.00035475999999999997 0 0.00035468 0 0.00035478 3.3 0.0003547 3.3 0.0003548 0 0.00035472 0 0.00035482 3.3 0.00035474 3.3 0.00035484 0 0.00035475999999999997 0 0.00035486 3.3 0.00035478 3.3 0.00035488 0 0.0003548 0 0.0003549 3.3 0.00035482 3.3 0.00035492 0 0.00035484 0 0.00035494 3.3 0.00035486 3.3 0.00035496 0 0.00035488 0 0.00035498 3.3 0.0003549 3.3 0.000355 0 0.00035492 0 0.00035502 3.3 0.00035494 3.3 0.00035504 0 0.00035496 0 0.00035506 3.3 0.00035497999999999997 3.3 0.00035507999999999997 0 0.000355 0 0.0003551 3.3 0.00035502 3.3 0.00035512 0 0.00035504 0 0.00035514 3.3 0.00035506 3.3 0.00035516 0 0.00035507999999999997 0 0.00035517999999999997 3.3 0.0003551 3.3 0.0003552 0 0.00035512 0 0.00035522 3.3 0.00035514 3.3 0.00035524 0 0.00035516 0 0.00035526 3.3 0.00035517999999999997 3.3 0.00035528 0 0.0003552 0 0.0003553 3.3 0.00035522 3.3 0.00035532 0 0.00035524 0 0.00035534 3.3 0.00035526 3.3 0.00035536 0 0.00035528 0 0.00035538 3.3 0.0003553 3.3 0.0003554 0 0.00035532 0 0.00035542 3.3 0.00035534 3.3 0.00035544 0 0.00035536 0 0.00035546 3.3 0.00035538 3.3 0.00035548 0 0.00035539999999999997 0 0.00035549999999999997 3.3 0.00035542 3.3 0.00035552 0 0.00035544 0 0.00035554 3.3 0.00035546 3.3 0.00035556 0 0.00035548 0 0.00035558 3.3 0.00035549999999999997 3.3 0.00035559999999999997 0 0.00035552 0 0.00035562 3.3 0.00035554 3.3 0.00035564 0 0.00035556 0 0.00035566 3.3 0.00035558 3.3 0.00035568 0 0.00035559999999999997 0 0.00035569999999999997 3.3 0.00035562 3.3 0.00035572 0 0.00035564 0 0.00035574 3.3 0.00035566 3.3 0.00035576 0 0.00035568 0 0.00035578 3.3 0.00035569999999999997 3.3 0.0003558 0 0.00035572 0 0.00035582 3.3 0.00035574 3.3 0.00035584 0 0.00035576 0 0.00035586 3.3 0.00035578 3.3 0.00035588 0 0.0003558 0 0.0003559 3.3 0.00035581999999999996 3.3 0.00035591999999999997 0 0.00035584 0 0.00035594 3.3 0.00035586 3.3 0.00035596 0 0.00035588 0 0.00035598 3.3 0.0003559 3.3 0.000356 0 0.00035591999999999997 0 0.00035601999999999997 3.3 0.00035594 3.3 0.00035604 0 0.00035596 0 0.00035606 3.3 0.00035598 3.3 0.00035608 0 0.000356 0 0.0003561 3.3 0.00035601999999999997 3.3 0.00035611999999999997 0 0.00035604 0 0.00035614 3.3 0.00035606 3.3 0.00035616 0 0.00035608 0 0.00035618 3.3 0.0003561 3.3 0.0003562 0 0.00035611999999999997 0 0.00035622 3.3 0.00035614 3.3 0.00035624 0 0.00035616 0 0.00035626 3.3 0.00035618 3.3 0.00035628 0 0.0003562 0 0.0003563 3.3 0.00035622 3.3 0.00035632 0 0.00035623999999999996 0 0.00035633999999999997 3.3 0.00035626 3.3 0.00035636 0 0.00035628 0 0.00035638 3.3 0.0003563 3.3 0.0003564 0 0.00035632 0 0.00035642 3.3 0.00035633999999999997 3.3 0.00035643999999999997 0 0.00035636 0 0.00035646 3.3 0.00035638 3.3 0.00035648 0 0.0003564 0 0.0003565 3.3 0.00035642 3.3 0.00035652 0 0.00035643999999999997 0 0.00035653999999999997 3.3 0.00035646 3.3 0.00035656 0 0.00035648 0 0.00035658 3.3 0.0003565 3.3 0.0003566 0 0.00035652 0 0.00035662 3.3 0.00035653999999999997 3.3 0.00035664 0 0.00035656 0 0.00035666 3.3 0.00035658 3.3 0.00035668 0 0.0003566 0 0.0003567 3.3 0.00035662 3.3 0.00035672 0 0.00035664 0 0.00035674 3.3 0.00035666 3.3 0.00035676 0 0.00035668 0 0.00035678 3.3 0.0003567 3.3 0.0003568 0 0.00035672 0 0.00035682 3.3 0.00035674 3.3 0.00035684 0 0.00035675999999999997 0 0.00035685999999999997 3.3 0.00035678 3.3 0.00035688 0 0.0003568 0 0.0003569 3.3 0.00035682 3.3 0.00035692 0 0.00035684 0 0.00035694 3.3 0.00035685999999999997 3.3 0.00035695999999999997 0 0.00035688 0 0.00035698 3.3 0.0003569 3.3 0.000357 0 0.00035692 0 0.00035702 3.3 0.00035694 3.3 0.00035704 0 0.00035695999999999997 0 0.00035705999999999997 3.3 0.00035698 3.3 0.00035708 0 0.000357 0 0.0003571 3.3 0.00035702 3.3 0.00035712 0 0.00035704 0 0.00035714 3.3 0.00035705999999999997 3.3 0.00035716 0 0.00035708 0 0.00035718 3.3 0.0003571 3.3 0.0003572 0 0.00035712 0 0.00035722 3.3 0.00035714 3.3 0.00035724 0 0.00035716 0 0.00035726 3.3 0.00035717999999999996 3.3 0.00035727999999999997 0 0.0003572 0 0.0003573 3.3 0.00035722 3.3 0.00035732 0 0.00035724 0 0.00035734 3.3 0.00035726 3.3 0.00035736 0 0.00035727999999999997 0 0.00035737999999999997 3.3 0.0003573 3.3 0.0003574 0 0.00035732 0 0.00035742 3.3 0.00035734 3.3 0.00035744 0 0.00035736 0 0.00035746 3.3 0.00035737999999999997 3.3 0.00035747999999999997 0 0.0003574 0 0.0003575 3.3 0.00035742 3.3 0.00035752 0 0.00035744 0 0.00035754 3.3 0.00035746 3.3 0.00035756 0 0.00035747999999999997 0 0.00035758 3.3 0.0003575 3.3 0.0003576 0 0.00035752 0 0.00035762 3.3 0.00035754 3.3 0.00035764 0 0.00035756 0 0.00035766 3.3 0.00035758 3.3 0.00035768 0 0.00035759999999999996 0 0.00035769999999999997 3.3 0.00035762 3.3 0.00035772 0 0.00035764 0 0.00035774 3.3 0.00035766 3.3 0.00035776 0 0.00035768 0 0.00035778 3.3 0.00035769999999999997 3.3 0.00035779999999999997 0 0.00035772 0 0.00035782 3.3 0.00035774 3.3 0.00035784 0 0.00035776 0 0.00035786 3.3 0.00035778 3.3 0.00035788 0 0.00035779999999999997 0 0.00035789999999999997 3.3 0.00035782 3.3 0.00035792 0 0.00035784 0 0.00035794 3.3 0.00035786 3.3 0.00035796 0 0.00035788 0 0.00035798 3.3 0.00035789999999999997 3.3 0.000358 0 0.00035792 0 0.00035802 3.3 0.00035794 3.3 0.00035804 0 0.00035796 0 0.00035806 3.3 0.00035798 3.3 0.00035808 0 0.000358 0 0.0003581 3.3 0.00035801999999999996 3.3 0.00035811999999999997 0 0.00035804 0 0.00035814 3.3 0.00035806 3.3 0.00035816 0 0.00035808 0 0.00035818 3.3 0.0003581 3.3 0.0003582 0 0.00035811999999999997 0 0.00035821999999999997 3.3 0.00035814 3.3 0.00035824 0 0.00035816 0 0.00035826 3.3 0.00035818 3.3 0.00035828 0 0.0003582 0 0.0003583 3.3 0.00035821999999999997 3.3 0.00035831999999999997 0 0.00035824 0 0.00035834 3.3 0.00035826 3.3 0.00035836 0 0.00035828 0 0.00035838 3.3 0.0003583 3.3 0.0003584 0 0.00035831999999999997 0 0.00035842 3.3 0.00035834 3.3 0.00035844 0 0.00035836 0 0.00035846 3.3 0.00035838 3.3 0.00035848 0 0.0003584 0 0.0003585 3.3 0.00035842 3.3 0.00035852 0 0.00035844 0 0.00035854 3.3 0.00035846 3.3 0.00035856 0 0.00035848 0 0.00035858 3.3 0.0003585 3.3 0.0003586 0 0.00035852 0 0.00035862 3.3 0.00035853999999999997 3.3 0.00035863999999999997 0 0.00035856 0 0.00035866 3.3 0.00035858 3.3 0.00035868 0 0.0003586 0 0.0003587 3.3 0.00035862 3.3 0.00035872 0 0.00035863999999999997 0 0.00035873999999999997 3.3 0.00035866 3.3 0.00035876 0 0.00035868 0 0.00035878 3.3 0.0003587 3.3 0.0003588 0 0.00035872 0 0.00035882 3.3 0.00035873999999999997 3.3 0.00035883999999999997 0 0.00035876 0 0.00035886 3.3 0.00035878 3.3 0.00035888 0 0.0003588 0 0.0003589 3.3 0.00035882 3.3 0.00035892 0 0.00035883999999999997 0 0.00035894 3.3 0.00035886 3.3 0.00035896 0 0.00035888 0 0.00035898 3.3 0.0003589 3.3 0.000359 0 0.00035892 0 0.00035902 3.3 0.00035894 3.3 0.00035904 0 0.00035895999999999996 0 0.00035905999999999997 3.3 0.00035898 3.3 0.00035908 0 0.000359 0 0.0003591 3.3 0.00035902 3.3 0.00035912 0 0.00035904 0 0.00035914 3.3 0.00035905999999999997 3.3 0.00035915999999999997 0 0.00035908 0 0.00035918 3.3 0.0003591 3.3 0.0003592 0 0.00035912 0 0.00035922 3.3 0.00035914 3.3 0.00035924 0 0.00035915999999999997 0 0.00035925999999999997 3.3 0.00035918 3.3 0.00035928 0 0.0003592 0 0.0003593 3.3 0.00035922 3.3 0.00035932 0 0.00035924 0 0.00035934 3.3 0.00035925999999999997 3.3 0.00035936 0 0.00035928 0 0.00035938 3.3 0.0003593 3.3 0.0003594 0 0.00035932 0 0.00035942 3.3 0.00035934 3.3 0.00035944 0 0.00035936 0 0.00035946 3.3 0.00035937999999999996 3.3 0.00035947999999999997 0 0.0003594 0 0.0003595 3.3 0.00035942 3.3 0.00035952 0 0.00035944 0 0.00035954 3.3 0.00035946 3.3 0.00035956 0 0.00035947999999999997 0 0.00035957999999999997 3.3 0.0003595 3.3 0.0003596 0 0.00035952 0 0.00035962 3.3 0.00035954 3.3 0.00035964 0 0.00035956 0 0.00035966 3.3 0.00035957999999999997 3.3 0.00035967999999999997 0 0.0003596 0 0.0003597 3.3 0.00035962 3.3 0.00035972 0 0.00035964 0 0.00035974 3.3 0.00035966 3.3 0.00035976 0 0.00035967999999999997 0 0.00035978 3.3 0.0003597 3.3 0.0003598 0 0.00035972 0 0.00035982 3.3 0.00035974 3.3 0.00035984 0 0.00035976 0 0.00035986 3.3 0.00035978 3.3 0.00035988 0 0.00035979999999999996 0 0.00035989999999999997 3.3 0.00035982 3.3 0.00035992 0 0.00035984 0 0.00035994 3.3 0.00035986 3.3 0.00035996 0 0.00035988 0 0.00035998 3.3 0.00035989999999999997 3.3 0.00035999999999999997 0 0.00035992 0 0.00036002 3.3 0.00035994 3.3 0.00036004 0 0.00035996 0 0.00036006 3.3 0.00035998 3.3 0.00036008 0 0.00035999999999999997 0 0.00036009999999999997 3.3 0.00036002 3.3 0.00036012 0 0.00036004 0 0.00036014 3.3 0.00036006 3.3 0.00036016 0 0.00036008 0 0.00036018 3.3 0.00036009999999999997 3.3 0.0003602 0 0.00036012 0 0.00036022 3.3 0.00036014 3.3 0.00036024 0 0.00036016 0 0.00036026 3.3 0.00036018 3.3 0.00036028 0 0.0003602 0 0.0003603 3.3 0.00036022 3.3 0.00036032 0 0.00036024 0 0.00036034 3.3 0.00036026 3.3 0.00036036 0 0.00036028 0 0.00036038 3.3 0.0003603 3.3 0.0003604 0 0.00036031999999999997 0 0.00036041999999999997 3.3 0.00036034 3.3 0.00036044 0 0.00036036 0 0.00036046 3.3 0.00036038 3.3 0.00036048 0 0.0003604 0 0.0003605 3.3 0.00036041999999999997 3.3 0.00036051999999999997 0 0.00036044 0 0.00036054 3.3 0.00036046 3.3 0.00036056 0 0.00036048 0 0.00036058 3.3 0.0003605 3.3 0.0003606 0 0.00036051999999999997 0 0.00036061999999999997 3.3 0.00036054 3.3 0.00036064 0 0.00036056 0 0.00036066 3.3 0.00036058 3.3 0.00036068 0 0.0003606 0 0.0003607 3.3 0.00036061999999999997 3.3 0.00036072 0 0.00036064 0 0.00036074 3.3 0.00036066 3.3 0.00036076 0 0.00036068 0 0.00036078 3.3 0.0003607 3.3 0.0003608 0 0.00036072 0 0.00036082 3.3 0.00036073999999999996 3.3 0.00036083999999999997 0 0.00036076 0 0.00036086 3.3 0.00036078 3.3 0.00036088 0 0.0003608 0 0.0003609 3.3 0.00036082 3.3 0.00036092 0 0.00036083999999999997 0 0.00036093999999999997 3.3 0.00036086 3.3 0.00036096 0 0.00036088 0 0.00036098 3.3 0.0003609 3.3 0.000361 0 0.00036092 0 0.00036102 3.3 0.00036093999999999997 3.3 0.00036103999999999997 0 0.00036096 0 0.00036106 3.3 0.00036098 3.3 0.00036108 0 0.000361 0 0.0003611 3.3 0.00036102 3.3 0.00036112 0 0.00036103999999999997 0 0.00036114 3.3 0.00036106 3.3 0.00036116 0 0.00036108 0 0.00036118 3.3 0.0003611 3.3 0.0003612 0 0.00036112 0 0.00036122 3.3 0.00036114 3.3 0.00036124 0 0.00036115999999999996 0 0.00036125999999999997 3.3 0.00036118 3.3 0.00036128 0 0.0003612 0 0.0003613 3.3 0.00036122 3.3 0.00036132 0 0.00036124 0 0.00036134 3.3 0.00036125999999999997 3.3 0.00036135999999999997 0 0.00036128 0 0.00036138 3.3 0.0003613 3.3 0.0003614 0 0.00036132 0 0.00036142 3.3 0.00036134 3.3 0.00036144 0 0.00036135999999999997 0 0.00036145999999999997 3.3 0.00036138 3.3 0.00036148 0 0.0003614 0 0.0003615 3.3 0.00036142 3.3 0.00036152 0 0.00036144 0 0.00036154 3.3 0.00036145999999999997 3.3 0.00036156 0 0.00036148 0 0.00036158 3.3 0.0003615 3.3 0.0003616 0 0.00036152 0 0.00036162 3.3 0.00036154 3.3 0.00036164 0 0.00036156 0 0.00036166 3.3 0.00036157999999999996 3.3 0.00036167999999999997 0 0.0003616 0 0.0003617 3.3 0.00036162 3.3 0.00036172 0 0.00036164 0 0.00036174 3.3 0.00036166 3.3 0.00036176 0 0.00036167999999999997 0 0.00036177999999999997 3.3 0.0003617 3.3 0.0003618 0 0.00036172 0 0.00036182 3.3 0.00036174 3.3 0.00036184 0 0.00036176 0 0.00036186 3.3 0.00036177999999999997 3.3 0.00036187999999999997 0 0.0003618 0 0.0003619 3.3 0.00036182 3.3 0.00036192 0 0.00036184 0 0.00036194 3.3 0.00036186 3.3 0.00036196 0 0.00036187999999999997 0 0.00036198 3.3 0.0003619 3.3 0.000362 0 0.00036192 0 0.00036202 3.3 0.00036194 3.3 0.00036204 0 0.00036196 0 0.00036206 3.3 0.00036198 3.3 0.00036208 0 0.000362 0 0.0003621 3.3 0.00036202 3.3 0.00036212 0 0.00036204 0 0.00036214 3.3 0.00036206 3.3 0.00036216 0 0.00036208 0 0.00036218 3.3 0.00036209999999999997 3.3 0.00036219999999999997 0 0.00036212 0 0.00036222 3.3 0.00036214 3.3 0.00036224 0 0.00036216 0 0.00036226 3.3 0.00036218 3.3 0.00036228 0 0.00036219999999999997 0 0.00036229999999999997 3.3 0.00036222 3.3 0.00036232 0 0.00036224 0 0.00036234 3.3 0.00036226 3.3 0.00036236 0 0.00036228 0 0.00036238 3.3 0.00036229999999999997 3.3 0.00036239999999999997 0 0.00036232 0 0.00036242 3.3 0.00036234 3.3 0.00036244 0 0.00036236 0 0.00036246 3.3 0.00036238 3.3 0.00036248 0 0.00036239999999999997 0 0.0003625 3.3 0.00036242 3.3 0.00036252 0 0.00036244 0 0.00036254 3.3 0.00036246 3.3 0.00036256 0 0.00036248 0 0.00036258 3.3 0.0003625 3.3 0.0003626 0 0.00036251999999999996 0 0.00036261999999999997 3.3 0.00036254 3.3 0.00036264 0 0.00036256 0 0.00036266 3.3 0.00036258 3.3 0.00036268 0 0.0003626 0 0.0003627 3.3 0.00036261999999999997 3.3 0.00036271999999999997 0 0.00036264 0 0.00036274 3.3 0.00036266 3.3 0.00036276 0 0.00036268 0 0.00036278 3.3 0.0003627 3.3 0.0003628 0 0.00036271999999999997 0 0.00036281999999999997 3.3 0.00036274 3.3 0.00036284 0 0.00036276 0 0.00036286 3.3 0.00036278 3.3 0.00036288 0 0.0003628 0 0.0003629 3.3 0.00036281999999999997 3.3 0.00036292 0 0.00036284 0 0.00036294 3.3 0.00036286 3.3 0.00036296 0 0.00036288 0 0.00036298 3.3 0.0003629 3.3 0.000363 0 0.00036292 0 0.00036302 3.3 0.00036293999999999996 3.3 0.00036303999999999997 0 0.00036296 0 0.00036306 3.3 0.00036298 3.3 0.00036308 0 0.000363 0 0.0003631 3.3 0.00036302 3.3 0.00036312 0 0.00036303999999999997 0 0.00036313999999999997 3.3 0.00036306 3.3 0.00036316 0 0.00036308 0 0.00036318 3.3 0.0003631 3.3 0.0003632 0 0.00036312 0 0.00036322 3.3 0.00036313999999999997 3.3 0.00036323999999999997 0 0.00036316 0 0.00036326 3.3 0.00036318 3.3 0.00036328 0 0.0003632 0 0.0003633 3.3 0.00036322 3.3 0.00036332 0 0.00036323999999999997 0 0.00036334 3.3 0.00036326 3.3 0.00036336 0 0.00036328 0 0.00036338 3.3 0.0003633 3.3 0.0003634 0 0.00036332 0 0.00036342 3.3 0.00036334 3.3 0.00036344 0 0.00036335999999999996 0 0.00036345999999999997 3.3 0.00036338 3.3 0.00036348 0 0.0003634 0 0.0003635 3.3 0.00036342 3.3 0.00036352 0 0.00036344 0 0.00036354 3.3 0.00036345999999999997 3.3 0.00036355999999999997 0 0.00036348 0 0.00036358 3.3 0.0003635 3.3 0.0003636 0 0.00036352 0 0.00036362 3.3 0.00036354 3.3 0.00036364 0 0.00036355999999999997 0 0.00036365999999999997 3.3 0.00036358 3.3 0.00036368 0 0.0003636 0 0.0003637 3.3 0.00036362 3.3 0.00036372 0 0.00036364 0 0.00036374 3.3 0.00036365999999999997 3.3 0.00036376 0 0.00036368 0 0.00036378 3.3 0.0003637 3.3 0.0003638 0 0.00036372 0 0.00036382 3.3 0.00036374 3.3 0.00036384 0 0.00036376 0 0.00036386 3.3 0.00036378 3.3 0.00036388 0 0.0003638 0 0.0003639 3.3 0.00036382 3.3 0.00036392 0 0.00036384 0 0.00036394 3.3 0.00036386 3.3 0.00036396 0 0.00036387999999999997 0 0.00036397999999999997 3.3 0.0003639 3.3 0.000364 0 0.00036392 0 0.00036402 3.3 0.00036394 3.3 0.00036404 0 0.00036396 0 0.00036406 3.3 0.00036397999999999997 3.3 0.00036407999999999997 0 0.000364 0 0.0003641 3.3 0.00036402 3.3 0.00036412 0 0.00036404 0 0.00036414 3.3 0.00036406 3.3 0.00036416 0 0.00036407999999999997 0 0.00036417999999999997 3.3 0.0003641 3.3 0.0003642 0 0.00036412 0 0.00036422 3.3 0.00036414 3.3 0.00036424 0 0.00036416 0 0.00036426 3.3 0.00036417999999999997 3.3 0.00036428 0 0.0003642 0 0.0003643 3.3 0.00036422 3.3 0.00036432 0 0.00036424 0 0.00036434 3.3 0.00036426 3.3 0.00036436 0 0.00036428 0 0.00036438 3.3 0.00036429999999999996 3.3 0.00036439999999999997 0 0.00036432 0 0.00036442 3.3 0.00036434 3.3 0.00036444 0 0.00036436 0 0.00036446 3.3 0.00036438 3.3 0.00036448 0 0.00036439999999999997 0 0.00036449999999999997 3.3 0.00036442 3.3 0.00036452 0 0.00036444 0 0.00036454 3.3 0.00036446 3.3 0.00036456 0 0.00036448 0 0.00036458 3.3 0.00036449999999999997 3.3 0.00036459999999999997 0 0.00036452 0 0.00036462 3.3 0.00036454 3.3 0.00036464 0 0.00036456 0 0.00036466 3.3 0.00036458 3.3 0.00036468 0 0.00036459999999999997 0 0.0003647 3.3 0.00036462 3.3 0.00036472 0 0.00036464 0 0.00036474 3.3 0.00036466 3.3 0.00036476 0 0.00036468 0 0.00036478 3.3 0.0003647 3.3 0.0003648 0 0.00036471999999999996 0 0.00036481999999999997 3.3 0.00036474 3.3 0.00036484 0 0.00036476 0 0.00036486 3.3 0.00036478 3.3 0.00036488 0 0.0003648 0 0.0003649 3.3 0.00036481999999999997 3.3 0.00036491999999999997 0 0.00036484 0 0.00036494 3.3 0.00036486 3.3 0.00036496 0 0.00036488 0 0.00036498 3.3 0.0003649 3.3 0.000365 0 0.00036491999999999997 0 0.00036501999999999997 3.3 0.00036494 3.3 0.00036504 0 0.00036496 0 0.00036506 3.3 0.00036498 3.3 0.00036508 0 0.000365 0 0.0003651 3.3 0.00036501999999999997 3.3 0.00036512 0 0.00036504 0 0.00036514 3.3 0.00036506 3.3 0.00036516 0 0.00036508 0 0.00036518 3.3 0.0003651 3.3 0.0003652 0 0.00036512 0 0.00036522 3.3 0.00036513999999999996 3.3 0.00036523999999999997 0 0.00036516 0 0.00036526 3.3 0.00036518 3.3 0.00036528 0 0.0003652 0 0.0003653 3.3 0.00036522 3.3 0.00036532 0 0.00036523999999999997 0 0.00036533999999999997 3.3 0.00036526 3.3 0.00036536 0 0.00036528 0 0.00036538 3.3 0.0003653 3.3 0.0003654 0 0.00036532 0 0.00036542 3.3 0.00036533999999999997 3.3 0.00036543999999999997 0 0.00036536 0 0.00036546 3.3 0.00036538 3.3 0.00036548 0 0.0003654 0 0.0003655 3.3 0.00036542 3.3 0.00036552 0 0.00036543999999999997 0 0.00036554 3.3 0.00036546 3.3 0.00036556 0 0.00036548 0 0.00036558 3.3 0.0003655 3.3 0.0003656 0 0.00036552 0 0.00036562 3.3 0.00036554 3.3 0.00036564 0 0.00036556 0 0.00036566 3.3 0.00036558 3.3 0.00036568 0 0.0003656 0 0.0003657 3.3 0.00036562 3.3 0.00036572 0 0.00036564 0 0.00036574 3.3 0.00036565999999999997 3.3 0.00036575999999999997 0 0.00036568 0 0.00036578 3.3 0.0003657 3.3 0.0003658 0 0.00036572 0 0.00036582 3.3 0.00036574 3.3 0.00036584 0 0.00036575999999999997 0 0.00036585999999999997 3.3 0.00036578 3.3 0.00036588 0 0.0003658 0 0.0003659 3.3 0.00036582 3.3 0.00036592 0 0.00036584 0 0.00036594 3.3 0.00036585999999999997 3.3 0.00036595999999999997 0 0.00036588 0 0.00036598 3.3 0.0003659 3.3 0.000366 0 0.00036592 0 0.00036602 3.3 0.00036594 3.3 0.00036604 0 0.00036595999999999997 0 0.00036606 3.3 0.00036598 3.3 0.00036608 0 0.000366 0 0.0003661 3.3 0.00036602 3.3 0.00036612 0 0.00036604 0 0.00036614 3.3 0.00036606 3.3 0.00036616 0 0.00036607999999999996 0 0.00036617999999999997 3.3 0.0003661 3.3 0.0003662 0 0.00036612 0 0.00036622 3.3 0.00036614 3.3 0.00036624 0 0.00036616 0 0.00036626 3.3 0.00036617999999999997 3.3 0.00036627999999999997 0 0.0003662 0 0.0003663 3.3 0.00036622 3.3 0.00036632 0 0.00036624 0 0.00036634 3.3 0.00036626 3.3 0.00036636 0 0.00036627999999999997 0 0.00036637999999999997 3.3 0.0003663 3.3 0.0003664 0 0.00036632 0 0.00036642 3.3 0.00036634 3.3 0.00036644 0 0.00036636 0 0.00036646 3.3 0.00036637999999999997 3.3 0.00036648 0 0.0003664 0 0.0003665 3.3 0.00036642 3.3 0.00036652 0 0.00036644 0 0.00036654 3.3 0.00036646 3.3 0.00036656 0 0.00036648 0 0.00036658 3.3 0.00036649999999999996 3.3 0.00036659999999999997 0 0.00036652 0 0.00036662 3.3 0.00036654 3.3 0.00036664 0 0.00036656 0 0.00036666 3.3 0.00036658 3.3 0.00036668 0 0.00036659999999999997 0 0.00036669999999999997 3.3 0.00036662 3.3 0.00036672 0 0.00036664 0 0.00036674 3.3 0.00036666 3.3 0.00036676 0 0.00036668 0 0.00036678 3.3 0.00036669999999999997 3.3 0.00036679999999999997 0 0.00036672 0 0.00036682 3.3 0.00036674 3.3 0.00036684 0 0.00036676 0 0.00036686 3.3 0.00036678 3.3 0.00036688 0 0.00036679999999999997 0 0.0003669 3.3 0.00036682 3.3 0.00036692 0 0.00036684 0 0.00036694 3.3 0.00036686 3.3 0.00036696 0 0.00036688 0 0.00036698 3.3 0.0003669 3.3 0.000367 0 0.00036691999999999996 0 0.00036701999999999997 3.3 0.00036694 3.3 0.00036704 0 0.00036696 0 0.00036706 3.3 0.00036698 3.3 0.00036708 0 0.000367 0 0.0003671 3.3 0.00036701999999999997 3.3 0.00036711999999999997 0 0.00036704 0 0.00036714 3.3 0.00036706 3.3 0.00036716 0 0.00036708 0 0.00036718 3.3 0.0003671 3.3 0.0003672 0 0.00036711999999999997 0 0.00036721999999999997 3.3 0.00036714 3.3 0.00036724 0 0.00036716 0 0.00036726 3.3 0.00036718 3.3 0.00036728 0 0.0003672 0 0.0003673 3.3 0.00036721999999999997 3.3 0.00036732 0 0.00036724 0 0.00036734 3.3 0.00036726 3.3 0.00036736 0 0.00036728 0 0.00036738 3.3 0.0003673 3.3 0.0003674 0 0.00036732 0 0.00036742 3.3 0.00036734 3.3 0.00036744 0 0.00036736 0 0.00036746 3.3 0.00036738 3.3 0.00036748 0 0.0003674 0 0.0003675 3.3 0.00036742 3.3 0.00036752 0 0.00036743999999999996 0 0.00036753999999999997 3.3 0.00036746 3.3 0.00036756 0 0.00036748 0 0.00036758 3.3 0.0003675 3.3 0.0003676 0 0.00036752 0 0.00036762 3.3 0.00036753999999999997 3.3 0.00036763999999999997 0 0.00036756 0 0.00036766 3.3 0.00036758 3.3 0.00036768 0 0.0003676 0 0.0003677 3.3 0.00036762 3.3 0.00036772 0 0.00036763999999999997 0 0.00036773999999999997 3.3 0.00036766 3.3 0.00036776 0 0.00036768 0 0.00036778 3.3 0.0003677 3.3 0.0003678 0 0.00036772 0 0.00036782 3.3 0.00036773999999999997 3.3 0.00036784 0 0.00036776 0 0.00036786 3.3 0.00036778 3.3 0.00036788 0 0.0003678 0 0.0003679 3.3 0.00036782 3.3 0.00036792 0 0.00036784 0 0.00036794 3.3 0.00036785999999999996 3.3 0.00036795999999999997 0 0.00036788 0 0.00036798 3.3 0.0003679 3.3 0.000368 0 0.00036792 0 0.00036802 3.3 0.00036794 3.3 0.00036804 0 0.00036795999999999997 0 0.00036805999999999997 3.3 0.00036798 3.3 0.00036808 0 0.000368 0 0.0003681 3.3 0.00036802 3.3 0.00036812 0 0.00036804 0 0.00036814 3.3 0.00036805999999999997 3.3 0.00036815999999999997 0 0.00036808 0 0.00036818 3.3 0.0003681 3.3 0.0003682 0 0.00036812 0 0.00036822 3.3 0.00036814 3.3 0.00036824 0 0.00036815999999999997 0 0.00036826 3.3 0.00036818 3.3 0.00036828 0 0.0003682 0 0.0003683 3.3 0.00036822 3.3 0.00036832 0 0.00036824 0 0.00036834 3.3 0.00036826 3.3 0.00036836 0 0.00036827999999999996 0 0.00036837999999999997 3.3 0.0003683 3.3 0.0003684 0 0.00036832 0 0.00036842 3.3 0.00036834 3.3 0.00036844 0 0.00036836 0 0.00036846 3.3 0.00036837999999999997 3.3 0.00036847999999999997 0 0.0003684 0 0.0003685 3.3 0.00036842 3.3 0.00036852 0 0.00036844 0 0.00036854 3.3 0.00036846 3.3 0.00036856 0 0.00036847999999999997 0 0.00036857999999999997 3.3 0.0003685 3.3 0.0003686 0 0.00036852 0 0.00036862 3.3 0.00036854 3.3 0.00036864 0 0.00036856 0 0.00036866 3.3 0.00036857999999999997 3.3 0.00036868 0 0.0003686 0 0.0003687 3.3 0.00036862 3.3 0.00036872 0 0.00036864 0 0.00036874 3.3 0.00036866 3.3 0.00036876 0 0.00036868 0 0.00036878 3.3 0.00036869999999999996 3.3 0.00036879999999999997 0 0.00036872 0 0.00036882 3.3 0.00036874 3.3 0.00036884 0 0.00036876 0 0.00036886 3.3 0.00036878 3.3 0.00036888 0 0.00036879999999999997 0 0.00036889999999999997 3.3 0.00036882 3.3 0.00036892 0 0.00036884 0 0.00036894 3.3 0.00036886 3.3 0.00036896 0 0.00036888 0 0.00036898 3.3 0.00036889999999999997 3.3 0.00036899999999999997 0 0.00036892 0 0.00036902 3.3 0.00036894 3.3 0.00036904 0 0.00036896 0 0.00036906 3.3 0.00036898 3.3 0.00036908 0 0.00036899999999999997 0 0.00036909999999999997 3.3 0.00036902 3.3 0.00036912 0 0.00036904 0 0.00036914 3.3 0.00036906 3.3 0.00036916 0 0.00036908 0 0.00036918 3.3 0.00036909999999999997 3.3 0.0003692 0 0.00036912 0 0.00036922 3.3 0.00036914 3.3 0.00036924 0 0.00036916 0 0.00036926 3.3 0.00036918 3.3 0.00036928 0 0.0003692 0 0.0003693 3.3 0.00036921999999999996 3.3 0.00036931999999999997 0 0.00036924 0 0.00036934 3.3 0.00036926 3.3 0.00036936 0 0.00036928 0 0.00036938 3.3 0.0003693 3.3 0.0003694 0 0.00036931999999999997 0 0.00036941999999999997 3.3 0.00036934 3.3 0.00036944 0 0.00036936 0 0.00036946 3.3 0.00036938 3.3 0.00036948 0 0.0003694 0 0.0003695 3.3 0.00036941999999999997 3.3 0.00036951999999999997 0 0.00036944 0 0.00036954 3.3 0.00036946 3.3 0.00036956 0 0.00036948 0 0.00036958 3.3 0.0003695 3.3 0.0003696 0 0.00036951999999999997 0 0.00036962 3.3 0.00036954 3.3 0.00036964 0 0.00036956 0 0.00036966 3.3 0.00036958 3.3 0.00036968 0 0.0003696 0 0.0003697 3.3 0.00036962 3.3 0.00036972 0 0.00036963999999999996 0 0.00036973999999999997 3.3 0.00036966 3.3 0.00036976 0 0.00036968 0 0.00036978 3.3 0.0003697 3.3 0.0003698 0 0.00036972 0 0.00036982 3.3 0.00036973999999999997 3.3 0.00036983999999999997 0 0.00036976 0 0.00036986 3.3 0.00036978 3.3 0.00036988 0 0.0003698 0 0.0003699 3.3 0.00036982 3.3 0.00036992 0 0.00036983999999999997 0 0.00036993999999999997 3.3 0.00036986 3.3 0.00036996 0 0.00036988 0 0.00036998 3.3 0.0003699 3.3 0.00037 0 0.00036992 0 0.00037002 3.3 0.00036993999999999997 3.3 0.00037004 0 0.00036996 0 0.00037006 3.3 0.00036998 3.3 0.00037008 0 0.00037 0 0.0003701 3.3 0.00037002 3.3 0.00037012 0 0.00037004 0 0.00037014 3.3 0.00037005999999999996 3.3 0.00037015999999999997 0 0.00037008 0 0.00037018 3.3 0.0003701 3.3 0.0003702 0 0.00037012 0 0.00037022 3.3 0.00037014 3.3 0.00037024 0 0.00037015999999999997 0 0.00037025999999999997 3.3 0.00037018 3.3 0.00037028 0 0.0003702 0 0.0003703 3.3 0.00037022 3.3 0.00037032 0 0.00037024 0 0.00037034 3.3 0.00037025999999999997 3.3 0.00037035999999999997 0 0.00037028 0 0.00037038 3.3 0.0003703 3.3 0.0003704 0 0.00037032 0 0.00037042 3.3 0.00037034 3.3 0.00037044 0 0.00037035999999999997 0 0.00037046 3.3 0.00037038 3.3 0.00037048 0 0.0003704 0 0.0003705 3.3 0.00037042 3.3 0.00037052 0 0.00037044 0 0.00037054 3.3 0.00037046 3.3 0.00037056 0 0.00037048 0 0.00037058 3.3 0.0003705 3.3 0.0003706 0 0.00037052 0 0.00037062 3.3 0.00037054 3.3 0.00037064 0 0.00037056 0 0.00037066 3.3 0.00037057999999999997 3.3 0.00037067999999999997 0 0.0003706 0 0.0003707 3.3 0.00037062 3.3 0.00037072 0 0.00037064 0 0.00037074 3.3 0.00037066 3.3 0.00037076 0 0.00037067999999999997 0 0.00037077999999999997 3.3 0.0003707 3.3 0.0003708 0 0.00037072 0 0.00037082 3.3 0.00037074 3.3 0.00037084 0 0.00037076 0 0.00037086 3.3 0.00037077999999999997 3.3 0.00037087999999999997 0 0.0003708 0 0.0003709 3.3 0.00037082 3.3 0.00037092 0 0.00037084 0 0.00037094 3.3 0.00037086 3.3 0.00037096 0 0.00037087999999999997 0 0.00037098 3.3 0.0003709 3.3 0.000371 0 0.00037092 0 0.00037102 3.3 0.00037094 3.3 0.00037104 0 0.00037096 0 0.00037106 3.3 0.00037098 3.3 0.00037108 0 0.00037099999999999996 0 0.00037109999999999997 3.3 0.00037102 3.3 0.00037112 0 0.00037104 0 0.00037114 3.3 0.00037106 3.3 0.00037116 0 0.00037108 0 0.00037118 3.3 0.00037109999999999997 3.3 0.00037119999999999997 0 0.00037112 0 0.00037122 3.3 0.00037114 3.3 0.00037124 0 0.00037116 0 0.00037126 3.3 0.00037118 3.3 0.00037128 0 0.00037119999999999997 0 0.00037129999999999997 3.3 0.00037122 3.3 0.00037132 0 0.00037124 0 0.00037134 3.3 0.00037126 3.3 0.00037136 0 0.00037128 0 0.00037138 3.3 0.00037129999999999997 3.3 0.0003714 0 0.00037132 0 0.00037142 3.3 0.00037134 3.3 0.00037144 0 0.00037136 0 0.00037146 3.3 0.00037138 3.3 0.00037148 0 0.0003714 0 0.0003715 3.3 0.00037141999999999996 3.3 0.00037151999999999997 0 0.00037144 0 0.00037154 3.3 0.00037146 3.3 0.00037156 0 0.00037148 0 0.00037158 3.3 0.0003715 3.3 0.0003716 0 0.00037151999999999997 0 0.00037161999999999997 3.3 0.00037154 3.3 0.00037164 0 0.00037156 0 0.00037166 3.3 0.00037158 3.3 0.00037168 0 0.0003716 0 0.0003717 3.3 0.00037161999999999997 3.3 0.00037171999999999997 0 0.00037164 0 0.00037174 3.3 0.00037166 3.3 0.00037176 0 0.00037168 0 0.00037178 3.3 0.0003717 3.3 0.0003718 0 0.00037171999999999997 0 0.00037182 3.3 0.00037174 3.3 0.00037184 0 0.00037176 0 0.00037186 3.3 0.00037178 3.3 0.00037188 0 0.0003718 0 0.0003719 3.3 0.00037182 3.3 0.00037192 0 0.00037183999999999996 0 0.00037193999999999997 3.3 0.00037186 3.3 0.00037196 0 0.00037188 0 0.00037198 3.3 0.0003719 3.3 0.000372 0 0.00037192 0 0.00037202 3.3 0.00037193999999999997 3.3 0.00037203999999999997 0 0.00037196 0 0.00037206 3.3 0.00037198 3.3 0.00037208 0 0.000372 0 0.0003721 3.3 0.00037202 3.3 0.00037212 0 0.00037203999999999997 0 0.00037213999999999997 3.3 0.00037206 3.3 0.00037216 0 0.00037208 0 0.00037218 3.3 0.0003721 3.3 0.0003722 0 0.00037212 0 0.00037222 3.3 0.00037213999999999997 3.3 0.00037224 0 0.00037216 0 0.00037226 3.3 0.00037218 3.3 0.00037228 0 0.0003722 0 0.0003723 3.3 0.00037222 3.3 0.00037232 0 0.00037224 0 0.00037234 3.3 0.00037226 3.3 0.00037236 0 0.00037228 0 0.00037238 3.3 0.0003723 3.3 0.0003724 0 0.00037232 0 0.00037242 3.3 0.00037234 3.3 0.00037244 0 0.00037235999999999997 0 0.00037245999999999997 3.3 0.00037238 3.3 0.00037248 0 0.0003724 0 0.0003725 3.3 0.00037242 3.3 0.00037252 0 0.00037244 0 0.00037254 3.3 0.00037245999999999997 3.3 0.00037255999999999997 0 0.00037248 0 0.00037258 3.3 0.0003725 3.3 0.0003726 0 0.00037252 0 0.00037262 3.3 0.00037254 3.3 0.00037264 0 0.00037255999999999997 0 0.00037265999999999997 3.3 0.00037258 3.3 0.00037268 0 0.0003726 0 0.0003727 3.3 0.00037262 3.3 0.00037272 0 0.00037264 0 0.00037274 3.3 0.00037265999999999997 3.3 0.00037276 0 0.00037268 0 0.00037278 3.3 0.0003727 3.3 0.0003728 0 0.00037272 0 0.00037282 3.3 0.00037274 3.3 0.00037284 0 0.00037276 0 0.00037286 3.3 0.00037277999999999996 3.3 0.00037287999999999997 0 0.0003728 0 0.0003729 3.3 0.00037282 3.3 0.00037292 0 0.00037284 0 0.00037294 3.3 0.00037286 3.3 0.00037296 0 0.00037287999999999997 0 0.00037297999999999997 3.3 0.0003729 3.3 0.000373 0 0.00037292 0 0.00037302 3.3 0.00037294 3.3 0.00037304 0 0.00037296 0 0.00037306 3.3 0.00037297999999999997 3.3 0.00037307999999999997 0 0.000373 0 0.0003731 3.3 0.00037302 3.3 0.00037312 0 0.00037304 0 0.00037314 3.3 0.00037306 3.3 0.00037316 0 0.00037307999999999997 0 0.00037318 3.3 0.0003731 3.3 0.0003732 0 0.00037312 0 0.00037322 3.3 0.00037314 3.3 0.00037324 0 0.00037316 0 0.00037326 3.3 0.00037318 3.3 0.00037328 0 0.00037319999999999996 0 0.00037329999999999997 3.3 0.00037322 3.3 0.00037332 0 0.00037324 0 0.00037334 3.3 0.00037326 3.3 0.00037336 0 0.00037328 0 0.00037338 3.3 0.00037329999999999997 3.3 0.00037339999999999997 0 0.00037332 0 0.00037342 3.3 0.00037334 3.3 0.00037344 0 0.00037336 0 0.00037346 3.3 0.00037338 3.3 0.00037348 0 0.00037339999999999997 0 0.00037349999999999997 3.3 0.00037342 3.3 0.00037352 0 0.00037344 0 0.00037354 3.3 0.00037346 3.3 0.00037356 0 0.00037348 0 0.00037358 3.3 0.00037349999999999997 3.3 0.0003736 0 0.00037352 0 0.00037362 3.3 0.00037354 3.3 0.00037364 0 0.00037356 0 0.00037366 3.3 0.00037358 3.3 0.00037368 0 0.0003736 0 0.0003737 3.3 0.00037361999999999996 3.3 0.00037371999999999997 0 0.00037364 0 0.00037374 3.3 0.00037366 3.3 0.00037376 0 0.00037368 0 0.00037378 3.3 0.0003737 3.3 0.0003738 0 0.00037371999999999997 0 0.00037381999999999997 3.3 0.00037374 3.3 0.00037384 0 0.00037376 0 0.00037386 3.3 0.00037378 3.3 0.00037388 0 0.0003738 0 0.0003739 3.3 0.00037381999999999997 3.3 0.00037391999999999997 0 0.00037384 0 0.00037394 3.3 0.00037386 3.3 0.00037396 0 0.00037388 0 0.00037398 3.3 0.0003739 3.3 0.000374 0 0.00037391999999999997 0 0.00037402 3.3 0.00037394 3.3 0.00037404 0 0.00037396 0 0.00037406 3.3 0.00037398 3.3 0.00037408 0 0.000374 0 0.0003741 3.3 0.00037402 3.3 0.00037412 0 0.00037404 0 0.00037414 3.3 0.00037406 3.3 0.00037416 0 0.00037408 0 0.00037418 3.3 0.0003741 3.3 0.0003742 0 0.00037412 0 0.00037422 3.3 0.00037413999999999997 3.3 0.00037423999999999997 0 0.00037416 0 0.00037426 3.3 0.00037418 3.3 0.00037428 0 0.0003742 0 0.0003743 3.3 0.00037422 3.3 0.00037432 0 0.00037423999999999997 0 0.00037433999999999997 3.3 0.00037426 3.3 0.00037436 0 0.00037428 0 0.00037438 3.3 0.0003743 3.3 0.0003744 0 0.00037432 0 0.00037442 3.3 0.00037433999999999997 3.3 0.00037443999999999997 0 0.00037436 0 0.00037446 3.3 0.00037438 3.3 0.00037448 0 0.0003744 0 0.0003745 3.3 0.00037442 3.3 0.00037452 0 0.00037443999999999997 0 0.00037454 3.3 0.00037446 3.3 0.00037456 0 0.00037448 0 0.00037458 3.3 0.0003745 3.3 0.0003746 0 0.00037452 0 0.00037462 3.3 0.00037454 3.3 0.00037464 0 0.00037455999999999996 0 0.00037465999999999997 3.3 0.00037458 3.3 0.00037468 0 0.0003746 0 0.0003747 3.3 0.00037462 3.3 0.00037472 0 0.00037464 0 0.00037474 3.3 0.00037465999999999997 3.3 0.00037475999999999997 0 0.00037468 0 0.00037478 3.3 0.0003747 3.3 0.0003748 0 0.00037472 0 0.00037482 3.3 0.00037474 3.3 0.00037484 0 0.00037475999999999997 0 0.00037485999999999997 3.3 0.00037478 3.3 0.00037488 0 0.0003748 0 0.0003749 3.3 0.00037482 3.3 0.00037492 0 0.00037484 0 0.00037494 3.3 0.00037485999999999997 3.3 0.00037496 0 0.00037488 0 0.00037498 3.3 0.0003749 3.3 0.000375 0 0.00037492 0 0.00037502 3.3 0.00037494 3.3 0.00037504 0 0.00037496 0 0.00037506 3.3 0.00037497999999999996 3.3 0.00037507999999999997 0 0.000375 0 0.0003751 3.3 0.00037502 3.3 0.00037512 0 0.00037504 0 0.00037514 3.3 0.00037506 3.3 0.00037516 0 0.00037507999999999997 0 0.00037517999999999997 3.3 0.0003751 3.3 0.0003752 0 0.00037512 0 0.00037522 3.3 0.00037514 3.3 0.00037524 0 0.00037516 0 0.00037526 3.3 0.00037517999999999997 3.3 0.00037527999999999997 0 0.0003752 0 0.0003753 3.3 0.00037522 3.3 0.00037532 0 0.00037524 0 0.00037534 3.3 0.00037526 3.3 0.00037536 0 0.00037527999999999997 0 0.00037538 3.3 0.0003753 3.3 0.0003754 0 0.00037532 0 0.00037542 3.3 0.00037534 3.3 0.00037544 0 0.00037536 0 0.00037546 3.3 0.00037538 3.3 0.00037548 0 0.00037539999999999996 0 0.00037549999999999997 3.3 0.00037542 3.3 0.00037552 0 0.00037544 0 0.00037554 3.3 0.00037546 3.3 0.00037556 0 0.00037548 0 0.00037558 3.3 0.00037549999999999997 3.3 0.00037559999999999997 0 0.00037552 0 0.00037562 3.3 0.00037554 3.3 0.00037564 0 0.00037556 0 0.00037566 3.3 0.00037558 3.3 0.00037568 0 0.00037559999999999997 0 0.00037569999999999997 3.3 0.00037562 3.3 0.00037572 0 0.00037564 0 0.00037574 3.3 0.00037566 3.3 0.00037576 0 0.00037568 0 0.00037578 3.3 0.00037569999999999997 3.3 0.0003758 0 0.00037572 0 0.00037582 3.3 0.00037574 3.3 0.00037584 0 0.00037576 0 0.00037586 3.3 0.00037578 3.3 0.00037588 0 0.0003758 0 0.0003759 3.3 0.00037582 3.3 0.00037592 0 0.00037584 0 0.00037594 3.3 0.00037586 3.3 0.00037596 0 0.00037588 0 0.00037598 3.3 0.0003759 3.3 0.000376 0 0.00037591999999999997 0 0.00037601999999999997 3.3 0.00037594 3.3 0.00037604 0 0.00037596 0 0.00037606 3.3 0.00037598 3.3 0.00037608 0 0.000376 0 0.0003761 3.3 0.00037601999999999997 3.3 0.00037611999999999997 0 0.00037604 0 0.00037614 3.3 0.00037606 3.3 0.00037616 0 0.00037608 0 0.00037618 3.3 0.0003761 3.3 0.0003762 0 0.00037611999999999997 0 0.00037621999999999997 3.3 0.00037614 3.3 0.00037624 0 0.00037616 0 0.00037626 3.3 0.00037618 3.3 0.00037628 0 0.0003762 0 0.0003763 3.3 0.00037621999999999997 3.3 0.00037632 0 0.00037624 0 0.00037634 3.3 0.00037626 3.3 0.00037636 0 0.00037628 0 0.00037638 3.3 0.0003763 3.3 0.0003764 0 0.00037632 0 0.00037642 3.3 0.00037633999999999996 3.3 0.00037643999999999997 0 0.00037636 0 0.00037646 3.3 0.00037638 3.3 0.00037648 0 0.0003764 0 0.0003765 3.3 0.00037642 3.3 0.00037652 0 0.00037643999999999997 0 0.00037653999999999997 3.3 0.00037646 3.3 0.00037656 0 0.00037648 0 0.00037658 3.3 0.0003765 3.3 0.0003766 0 0.00037652 0 0.00037662 3.3 0.00037653999999999997 3.3 0.00037663999999999997 0 0.00037656 0 0.00037666 3.3 0.00037658 3.3 0.00037668 0 0.0003766 0 0.0003767 3.3 0.00037662 3.3 0.00037672 0 0.00037663999999999997 0 0.00037674 3.3 0.00037666 3.3 0.00037676 0 0.00037668 0 0.00037678 3.3 0.0003767 3.3 0.0003768 0 0.00037672 0 0.00037682 3.3 0.00037674 3.3 0.00037684 0 0.00037675999999999996 0 0.00037685999999999997 3.3 0.00037678 3.3 0.00037688 0 0.0003768 0 0.0003769 3.3 0.00037682 3.3 0.00037692 0 0.00037684 0 0.00037694 3.3 0.00037685999999999997 3.3 0.00037695999999999997 0 0.00037688 0 0.00037698 3.3 0.0003769 3.3 0.000377 0 0.00037692 0 0.00037702 3.3 0.00037694 3.3 0.00037704 0 0.00037695999999999997 0 0.00037705999999999997 3.3 0.00037698 3.3 0.00037708 0 0.000377 0 0.0003771 3.3 0.00037702 3.3 0.00037712 0 0.00037704 0 0.00037714 3.3 0.00037705999999999997 3.3 0.00037716 0 0.00037708 0 0.00037718 3.3 0.0003771 3.3 0.0003772 0 0.00037712 0 0.00037722 3.3 0.00037714 3.3 0.00037724 0 0.00037716 0 0.00037726 3.3 0.00037717999999999996 3.3 0.00037727999999999997 0 0.0003772 0 0.0003773 3.3 0.00037722 3.3 0.00037732 0 0.00037724 0 0.00037734 3.3 0.00037726 3.3 0.00037736 0 0.00037727999999999997 0 0.00037737999999999997 3.3 0.0003773 3.3 0.0003774 0 0.00037732 0 0.00037742 3.3 0.00037734 3.3 0.00037744 0 0.00037736 0 0.00037746 3.3 0.00037737999999999997 3.3 0.00037747999999999997 0 0.0003774 0 0.0003775 3.3 0.00037742 3.3 0.00037752 0 0.00037744 0 0.00037754 3.3 0.00037746 3.3 0.00037756 0 0.00037747999999999997 0 0.00037758 3.3 0.0003775 3.3 0.0003776 0 0.00037752 0 0.00037762 3.3 0.00037754 3.3 0.00037764 0 0.00037756 0 0.00037766 3.3 0.00037758 3.3 0.00037768 0 0.0003776 0 0.0003777 3.3 0.00037762 3.3 0.00037772 0 0.00037764 0 0.00037774 3.3 0.00037766 3.3 0.00037776 0 0.00037768 0 0.00037778 3.3 0.00037769999999999997 3.3 0.00037779999999999997 0 0.00037772 0 0.00037782 3.3 0.00037774 3.3 0.00037784 0 0.00037776 0 0.00037786 3.3 0.00037778 3.3 0.00037788 0 0.00037779999999999997 0 0.00037789999999999997 3.3 0.00037782 3.3 0.00037792 0 0.00037784 0 0.00037794 3.3 0.00037786 3.3 0.00037796 0 0.00037788 0 0.00037798 3.3 0.00037789999999999997 3.3 0.00037799999999999997 0 0.00037792 0 0.00037802 3.3 0.00037794 3.3 0.00037804 0 0.00037796 0 0.00037806 3.3 0.00037798 3.3 0.00037808 0 0.00037799999999999997 0 0.0003781 3.3 0.00037802 3.3 0.00037812 0 0.00037804 0 0.00037814 3.3 0.00037806 3.3 0.00037816 0 0.00037808 0 0.00037818 3.3 0.0003781 3.3 0.0003782 0 0.00037811999999999996 0 0.00037821999999999997 3.3 0.00037814 3.3 0.00037824 0 0.00037816 0 0.00037826 3.3 0.00037818 3.3 0.00037828 0 0.0003782 0 0.0003783 3.3 0.00037821999999999997 3.3 0.00037831999999999997 0 0.00037824 0 0.00037834 3.3 0.00037826 3.3 0.00037836 0 0.00037828 0 0.00037838 3.3 0.0003783 3.3 0.0003784 0 0.00037831999999999997 0 0.00037841999999999997 3.3 0.00037834 3.3 0.00037844 0 0.00037836 0 0.00037846 3.3 0.00037838 3.3 0.00037848 0 0.0003784 0 0.0003785 3.3 0.00037841999999999997 3.3 0.00037852 0 0.00037844 0 0.00037854 3.3 0.00037846 3.3 0.00037856 0 0.00037848 0 0.00037858 3.3 0.0003785 3.3 0.0003786 0 0.00037852 0 0.00037862 3.3 0.00037853999999999996 3.3 0.00037863999999999997 0 0.00037856 0 0.00037866 3.3 0.00037858 3.3 0.00037868 0 0.0003786 0 0.0003787 3.3 0.00037862 3.3 0.00037872 0 0.00037863999999999997 0 0.00037873999999999997 3.3 0.00037866 3.3 0.00037876 0 0.00037868 0 0.00037878 3.3 0.0003787 3.3 0.0003788 0 0.00037872 0 0.00037882 3.3 0.00037873999999999997 3.3 0.00037883999999999997 0 0.00037876 0 0.00037886 3.3 0.00037878 3.3 0.00037888 0 0.0003788 0 0.0003789 3.3 0.00037882 3.3 0.00037892 0 0.00037883999999999997 0 0.00037894 3.3 0.00037886 3.3 0.00037896 0 0.00037888 0 0.00037898 3.3 0.0003789 3.3 0.000379 0 0.00037892 0 0.00037902 3.3 0.00037894 3.3 0.00037904 0 0.00037895999999999996 0 0.00037905999999999997 3.3 0.00037898 3.3 0.00037908 0 0.000379 0 0.0003791 3.3 0.00037902 3.3 0.00037912 0 0.00037904 0 0.00037914 3.3 0.00037905999999999997 3.3 0.00037915999999999997 0 0.00037908 0 0.00037918 3.3 0.0003791 3.3 0.0003792 0 0.00037912 0 0.00037922 3.3 0.00037914 3.3 0.00037924 0 0.00037915999999999997 0 0.00037925999999999997 3.3 0.00037918 3.3 0.00037928 0 0.0003792 0 0.0003793 3.3 0.00037922 3.3 0.00037932 0 0.00037924 0 0.00037934 3.3 0.00037925999999999997 3.3 0.00037935999999999997 0 0.00037928 0 0.00037938 3.3 0.0003793 3.3 0.0003794 0 0.00037932 0 0.00037942 3.3 0.00037934 3.3 0.00037944 0 0.00037935999999999997 0 0.00037946 3.3 0.00037938 3.3 0.00037948 0 0.0003794 0 0.0003795 3.3 0.00037942 3.3 0.00037952 0 0.00037944 0 0.00037954 3.3 0.00037946 3.3 0.00037956 0 0.00037947999999999996 0 0.00037957999999999997 3.3 0.0003795 3.3 0.0003796 0 0.00037952 0 0.00037962 3.3 0.00037954 3.3 0.00037964 0 0.00037956 0 0.00037966 3.3 0.00037957999999999997 3.3 0.00037967999999999997 0 0.0003796 0 0.0003797 3.3 0.00037962 3.3 0.00037972 0 0.00037964 0 0.00037974 3.3 0.00037966 3.3 0.00037976 0 0.00037967999999999997 0 0.00037977999999999997 3.3 0.0003797 3.3 0.0003798 0 0.00037972 0 0.00037982 3.3 0.00037974 3.3 0.00037984 0 0.00037976 0 0.00037986 3.3 0.00037977999999999997 3.3 0.00037988 0 0.0003798 0 0.0003799 3.3 0.00037982 3.3 0.00037992 0 0.00037984 0 0.00037994 3.3 0.00037986 3.3 0.00037996 0 0.00037988 0 0.00037998 3.3 0.00037989999999999996 3.3 0.00037999999999999997 0 0.00037992 0 0.00038002 3.3 0.00037994 3.3 0.00038004 0 0.00037996 0 0.00038006 3.3 0.00037998 3.3 0.00038008 0 0.00037999999999999997 0 0.00038009999999999997 3.3 0.00038002 3.3 0.00038012 0 0.00038004 0 0.00038014 3.3 0.00038006 3.3 0.00038016 0 0.00038008 0 0.00038018 3.3 0.00038009999999999997 3.3 0.00038019999999999997 0 0.00038012 0 0.00038022 3.3 0.00038014 3.3 0.00038024 0 0.00038016 0 0.00038026 3.3 0.00038018 3.3 0.00038028 0 0.00038019999999999997 0 0.0003803 3.3 0.00038022 3.3 0.00038032 0 0.00038024 0 0.00038034 3.3 0.00038026 3.3 0.00038036 0 0.00038028 0 0.00038038 3.3 0.0003803 3.3 0.0003804 0 0.00038031999999999996 0 0.00038041999999999997 3.3 0.00038034 3.3 0.00038044 0 0.00038036 0 0.00038046 3.3 0.00038038 3.3 0.00038048 0 0.0003804 0 0.0003805 3.3 0.00038041999999999997 3.3 0.00038051999999999997 0 0.00038044 0 0.00038054 3.3 0.00038046 3.3 0.00038056 0 0.00038048 0 0.00038058 3.3 0.0003805 3.3 0.0003806 0 0.00038051999999999997 0 0.00038061999999999997 3.3 0.00038054 3.3 0.00038064 0 0.00038056 0 0.00038066 3.3 0.00038058 3.3 0.00038068 0 0.0003806 0 0.0003807 3.3 0.00038061999999999997 3.3 0.00038072 0 0.00038064 0 0.00038074 3.3 0.00038066 3.3 0.00038076 0 0.00038068 0 0.00038078 3.3 0.0003807 3.3 0.0003808 0 0.00038072 0 0.00038082 3.3 0.00038073999999999996 3.3 0.00038083999999999997 0 0.00038076 0 0.00038086 3.3 0.00038078 3.3 0.00038088 0 0.0003808 0 0.0003809 3.3 0.00038082 3.3 0.00038092 0 0.00038083999999999997 0 0.00038093999999999997 3.3 0.00038086 3.3 0.00038096 0 0.00038088 0 0.00038098 3.3 0.0003809 3.3 0.000381 0 0.00038092 0 0.00038102 3.3 0.00038093999999999997 3.3 0.00038103999999999997 0 0.00038096 0 0.00038106 3.3 0.00038098 3.3 0.00038108 0 0.000381 0 0.0003811 3.3 0.00038102 3.3 0.00038112 0 0.00038103999999999997 0 0.00038113999999999997 3.3 0.00038106 3.3 0.00038116 0 0.00038108 0 0.00038118 3.3 0.0003811 3.3 0.0003812 0 0.00038112 0 0.00038122 3.3 0.00038113999999999997 3.3 0.00038124 0 0.00038116 0 0.00038126 3.3 0.00038118 3.3 0.00038128 0 0.0003812 0 0.0003813 3.3 0.00038122 3.3 0.00038132 0 0.00038124 0 0.00038134 3.3 0.00038125999999999996 3.3 0.00038135999999999997 0 0.00038128 0 0.00038138 3.3 0.0003813 3.3 0.0003814 0 0.00038132 0 0.00038142 3.3 0.00038134 3.3 0.00038144 0 0.00038135999999999997 0 0.00038145999999999997 3.3 0.00038138 3.3 0.00038148 0 0.0003814 0 0.0003815 3.3 0.00038142 3.3 0.00038152 0 0.00038144 0 0.00038154 3.3 0.00038145999999999997 3.3 0.00038155999999999997 0 0.00038148 0 0.00038158 3.3 0.0003815 3.3 0.0003816 0 0.00038152 0 0.00038162 3.3 0.00038154 3.3 0.00038164 0 0.00038155999999999997 0 0.00038166 3.3 0.00038158 3.3 0.00038168 0 0.0003816 0 0.0003817 3.3 0.00038162 3.3 0.00038172 0 0.00038164 0 0.00038174 3.3 0.00038166 3.3 0.00038176 0 0.00038167999999999996 0 0.00038177999999999997 3.3 0.0003817 3.3 0.0003818 0 0.00038172 0 0.00038182 3.3 0.00038174 3.3 0.00038184 0 0.00038176 0 0.00038186 3.3 0.00038177999999999997 3.3 0.00038187999999999997 0 0.0003818 0 0.0003819 3.3 0.00038182 3.3 0.00038192 0 0.00038184 0 0.00038194 3.3 0.00038186 3.3 0.00038196 0 0.00038187999999999997 0 0.00038197999999999997 3.3 0.0003819 3.3 0.000382 0 0.00038192 0 0.00038202 3.3 0.00038194 3.3 0.00038204 0 0.00038196 0 0.00038206 3.3 0.00038197999999999997 3.3 0.00038208 0 0.000382 0 0.0003821 3.3 0.00038202 3.3 0.00038212 0 0.00038204 0 0.00038214 3.3 0.00038206 3.3 0.00038216 0 0.00038208 0 0.00038218 3.3 0.00038209999999999996 3.3 0.00038219999999999997 0 0.00038212 0 0.00038222 3.3 0.00038214 3.3 0.00038224 0 0.00038216 0 0.00038226 3.3 0.00038218 3.3 0.00038228 0 0.00038219999999999997 0 0.00038229999999999997 3.3 0.00038222 3.3 0.00038232 0 0.00038224 0 0.00038234 3.3 0.00038226 3.3 0.00038236 0 0.00038228 0 0.00038238 3.3 0.00038229999999999997 3.3 0.00038239999999999997 0 0.00038232 0 0.00038242 3.3 0.00038234 3.3 0.00038244 0 0.00038236 0 0.00038246 3.3 0.00038238 3.3 0.00038248 0 0.00038239999999999997 0 0.0003825 3.3 0.00038242 3.3 0.00038252 0 0.00038244 0 0.00038254 3.3 0.00038246 3.3 0.00038256 0 0.00038248 0 0.00038258 3.3 0.0003825 3.3 0.0003826 0 0.00038251999999999996 0 0.00038261999999999997 3.3 0.00038254 3.3 0.00038264 0 0.00038256 0 0.00038266 3.3 0.00038258 3.3 0.00038268 0 0.0003826 0 0.0003827 3.3 0.00038261999999999997 3.3 0.00038271999999999997 0 0.00038264 0 0.00038274 3.3 0.00038266 3.3 0.00038276 0 0.00038268 0 0.00038278 3.3 0.0003827 3.3 0.0003828 0 0.00038271999999999997 0 0.00038281999999999997 3.3 0.00038274 3.3 0.00038284 0 0.00038276 0 0.00038286 3.3 0.00038278 3.3 0.00038288 0 0.0003828 0 0.0003829 3.3 0.00038281999999999997 3.3 0.00038291999999999997 0 0.00038284 0 0.00038294 3.3 0.00038286 3.3 0.00038296 0 0.00038288 0 0.00038298 3.3 0.0003829 3.3 0.000383 0 0.00038291999999999997 0 0.00038302 3.3 0.00038294 3.3 0.00038304 0 0.00038296 0 0.00038306 3.3 0.00038298 3.3 0.00038308 0 0.000383 0 0.0003831 3.3 0.00038302 3.3 0.00038312 0 0.00038303999999999996 0 0.00038313999999999997 3.3 0.00038306 3.3 0.00038316 0 0.00038308 0 0.00038318 3.3 0.0003831 3.3 0.0003832 0 0.00038312 0 0.00038322 3.3 0.00038313999999999997 3.3 0.00038323999999999997 0 0.00038316 0 0.00038326 3.3 0.00038318 3.3 0.00038328 0 0.0003832 0 0.0003833 3.3 0.00038322 3.3 0.00038332 0 0.00038323999999999997 0 0.00038333999999999997 3.3 0.00038326 3.3 0.00038336 0 0.00038328 0 0.00038338 3.3 0.0003833 3.3 0.0003834 0 0.00038332 0 0.00038342 3.3 0.00038333999999999997 3.3 0.00038344 0 0.00038336 0 0.00038346 3.3 0.00038338 3.3 0.00038348 0 0.0003834 0 0.0003835 3.3 0.00038342 3.3 0.00038352 0 0.00038344 0 0.00038354 3.3 0.00038345999999999996 3.3 0.00038355999999999997 0 0.00038348 0 0.00038358 3.3 0.0003835 3.3 0.0003836 0 0.00038352 0 0.00038362 3.3 0.00038354 3.3 0.00038364 0 0.00038355999999999997 0 0.00038365999999999997 3.3 0.00038358 3.3 0.00038368 0 0.0003836 0 0.0003837 3.3 0.00038362 3.3 0.00038372 0 0.00038364 0 0.00038374 3.3 0.00038365999999999997 3.3 0.00038375999999999997 0 0.00038368 0 0.00038378 3.3 0.0003837 3.3 0.0003838 0 0.00038372 0 0.00038382 3.3 0.00038374 3.3 0.00038384 0 0.00038375999999999997 0 0.00038386 3.3 0.00038378 3.3 0.00038388 0 0.0003838 0 0.0003839 3.3 0.00038382 3.3 0.00038392 0 0.00038384 0 0.00038394 3.3 0.00038386 3.3 0.00038396 0 0.00038387999999999996 0 0.00038397999999999997 3.3 0.0003839 3.3 0.000384 0 0.00038392 0 0.00038402 3.3 0.00038394 3.3 0.00038404 0 0.00038396 0 0.00038406 3.3 0.00038397999999999997 3.3 0.00038407999999999997 0 0.000384 0 0.0003841 3.3 0.00038402 3.3 0.00038412 0 0.00038404 0 0.00038414 3.3 0.00038406 3.3 0.00038416 0 0.00038407999999999997 0 0.00038417999999999997 3.3 0.0003841 3.3 0.0003842 0 0.00038412 0 0.00038422 3.3 0.00038414 3.3 0.00038424 0 0.00038416 0 0.00038426 3.3 0.00038417999999999997 3.3 0.00038428 0 0.0003842 0 0.0003843 3.3 0.00038422 3.3 0.00038432 0 0.00038424 0 0.00038434 3.3 0.00038426 3.3 0.00038436 0 0.00038428 0 0.00038438 3.3 0.00038429999999999996 3.3 0.00038439999999999997 0 0.00038432 0 0.00038442 3.3 0.00038434 3.3 0.00038444 0 0.00038436 0 0.00038446 3.3 0.00038438 3.3 0.00038448 0 0.00038439999999999997 0 0.00038449999999999997 3.3 0.00038442 3.3 0.00038452 0 0.00038444 0 0.00038454 3.3 0.00038446 3.3 0.00038456 0 0.00038448 0 0.00038458 3.3 0.00038449999999999997 3.3 0.00038459999999999997 0 0.00038452 0 0.00038462 3.3 0.00038454 3.3 0.00038464 0 0.00038456 0 0.00038466 3.3 0.00038458 3.3 0.00038468 0 0.00038459999999999997 0 0.00038469999999999997 3.3 0.00038462 3.3 0.00038472 0 0.00038464 0 0.00038474 3.3 0.00038466 3.3 0.00038476 0 0.00038468 0 0.00038478 3.3 0.00038469999999999997 3.3 0.0003848 0 0.00038472 0 0.00038482 3.3 0.00038474 3.3 0.00038484 0 0.00038476 0 0.00038486 3.3 0.00038478 3.3 0.00038488 0 0.0003848 0 0.0003849 3.3 0.00038481999999999996 3.3 0.00038491999999999997 0 0.00038484 0 0.00038494 3.3 0.00038486 3.3 0.00038496 0 0.00038488 0 0.00038498 3.3 0.0003849 3.3 0.000385 0 0.00038491999999999997 0 0.00038501999999999997 3.3 0.00038494 3.3 0.00038504 0 0.00038496 0 0.00038506 3.3 0.00038498 3.3 0.00038508 0 0.000385 0 0.0003851 3.3 0.00038501999999999997 3.3 0.00038511999999999997 0 0.00038504 0 0.00038514 3.3 0.00038506 3.3 0.00038516 0 0.00038508 0 0.00038518 3.3 0.0003851 3.3 0.0003852 0 0.00038511999999999997 0 0.00038522 3.3 0.00038514 3.3 0.00038524 0 0.00038516 0 0.00038526 3.3 0.00038518 3.3 0.00038528 0 0.0003852 0 0.0003853 3.3 0.00038522 3.3 0.00038532 0 0.00038523999999999996 0 0.00038533999999999997 3.3 0.00038526 3.3 0.00038536 0 0.00038528 0 0.00038538 3.3 0.0003853 3.3 0.0003854 0 0.00038532 0 0.00038542 3.3 0.00038533999999999997 3.3 0.00038543999999999997 0 0.00038536 0 0.00038546 3.3 0.00038538 3.3 0.00038548 0 0.0003854 0 0.0003855 3.3 0.00038542 3.3 0.00038552 0 0.00038543999999999997 0 0.00038553999999999997 3.3 0.00038546 3.3 0.00038556 0 0.00038548 0 0.00038558 3.3 0.0003855 3.3 0.0003856 0 0.00038552 0 0.00038562 3.3 0.00038553999999999997 3.3 0.00038564 0 0.00038556 0 0.00038566 3.3 0.00038558 3.3 0.00038568 0 0.0003856 0 0.0003857 3.3 0.00038562 3.3 0.00038572 0 0.00038564 0 0.00038574 3.3 0.00038565999999999996 3.3 0.00038575999999999997 0 0.00038568 0 0.00038578 3.3 0.0003857 3.3 0.0003858 0 0.00038572 0 0.00038582 3.3 0.00038574 3.3 0.00038584 0 0.00038575999999999997 0 0.00038585999999999997 3.3 0.00038578 3.3 0.00038588 0 0.0003858 0 0.0003859 3.3 0.00038582 3.3 0.00038592 0 0.00038584 0 0.00038594 3.3 0.00038585999999999997 3.3 0.00038595999999999997 0 0.00038588 0 0.00038598 3.3 0.0003859 3.3 0.000386 0 0.00038592 0 0.00038602 3.3 0.00038594 3.3 0.00038604 0 0.00038595999999999997 0 0.00038606 3.3 0.00038598 3.3 0.00038608 0 0.000386 0 0.0003861 3.3 0.00038602 3.3 0.00038612 0 0.00038604 0 0.00038614 3.3 0.00038606 3.3 0.00038616 0 0.00038607999999999996 0 0.00038617999999999997 3.3 0.0003861 3.3 0.0003862 0 0.00038612 0 0.00038622 3.3 0.00038614 3.3 0.00038624 0 0.00038616 0 0.00038626 3.3 0.00038617999999999997 3.3 0.00038627999999999997 0 0.0003862 0 0.0003863 3.3 0.00038622 3.3 0.00038632 0 0.00038624 0 0.00038634 3.3 0.00038626 3.3 0.00038636 0 0.00038627999999999997 0 0.00038637999999999997 3.3 0.0003863 3.3 0.0003864 0 0.00038632 0 0.00038642 3.3 0.00038634 3.3 0.00038644 0 0.00038636 0 0.00038646 3.3 0.00038637999999999997 3.3 0.00038647999999999997 0 0.0003864 0 0.0003865 3.3 0.00038642 3.3 0.00038652 0 0.00038644 0 0.00038654 3.3 0.00038646 3.3 0.00038656 0 0.00038647999999999997 0 0.00038658 3.3 0.0003865 3.3 0.0003866 0 0.00038652 0 0.00038662 3.3 0.00038654 3.3 0.00038664 0 0.00038656 0 0.00038666 3.3 0.00038658 3.3 0.00038668 0 0.00038659999999999996 0 0.00038669999999999997 3.3 0.00038662 3.3 0.00038672 0 0.00038664 0 0.00038674 3.3 0.00038666 3.3 0.00038676 0 0.00038668 0 0.00038678 3.3 0.00038669999999999997 3.3 0.00038679999999999997 0 0.00038672 0 0.00038682 3.3 0.00038674 3.3 0.00038684 0 0.00038676 0 0.00038686 3.3 0.00038678 3.3 0.00038688 0 0.00038679999999999997 0 0.00038689999999999997 3.3 0.00038682 3.3 0.00038692 0 0.00038684 0 0.00038694 3.3 0.00038686 3.3 0.00038696 0 0.00038688 0 0.00038698 3.3 0.00038689999999999997 3.3 0.000387 0 0.00038692 0 0.00038702 3.3 0.00038694 3.3 0.00038704 0 0.00038696 0 0.00038706 3.3 0.00038698 3.3 0.00038708 0 0.000387 0 0.0003871 3.3 0.00038701999999999996 3.3 0.00038711999999999997 0 0.00038704 0 0.00038714 3.3 0.00038706 3.3 0.00038716 0 0.00038708 0 0.00038718 3.3 0.0003871 3.3 0.0003872 0 0.00038711999999999997 0 0.00038721999999999997 3.3 0.00038714 3.3 0.00038724 0 0.00038716 0 0.00038726 3.3 0.00038718 3.3 0.00038728 0 0.0003872 0 0.0003873 3.3 0.00038721999999999997 3.3 0.00038731999999999997 0 0.00038724 0 0.00038734 3.3 0.00038726 3.3 0.00038736 0 0.00038728 0 0.00038738 3.3 0.0003873 3.3 0.0003874 0 0.00038731999999999997 0 0.00038742 3.3 0.00038734 3.3 0.00038744 0 0.00038736 0 0.00038746 3.3 0.00038738 3.3 0.00038748 0 0.0003874 0 0.0003875 3.3 0.00038742 3.3 0.00038752 0 0.00038743999999999996 0 0.00038753999999999997 3.3 0.00038746 3.3 0.00038756 0 0.00038748 0 0.00038758 3.3 0.0003875 3.3 0.0003876 0 0.00038752 0 0.00038762 3.3 0.00038753999999999997 3.3 0.00038763999999999997 0 0.00038756 0 0.00038766 3.3 0.00038758 3.3 0.00038768 0 0.0003876 0 0.0003877 3.3 0.00038762 3.3 0.00038772 0 0.00038763999999999997 0 0.00038773999999999997 3.3 0.00038766 3.3 0.00038776 0 0.00038768 0 0.00038778 3.3 0.0003877 3.3 0.0003878 0 0.00038772 0 0.00038782 3.3 0.00038773999999999997 3.3 0.00038784 0 0.00038776 0 0.00038786 3.3 0.00038778 3.3 0.00038788 0 0.0003878 0 0.0003879 3.3 0.00038782 3.3 0.00038792 0 0.00038784 0 0.00038794 3.3 0.00038786 3.3 0.00038796 0 0.00038788 0 0.00038798 3.3 0.0003879 3.3 0.000388 0 0.00038792 0 0.00038802 3.3 0.00038794 3.3 0.00038804 0 0.00038795999999999997 0 0.00038805999999999997 3.3 0.00038798 3.3 0.00038808 0 0.000388 0 0.0003881 3.3 0.00038802 3.3 0.00038812 0 0.00038804 0 0.00038814 3.3 0.00038805999999999997 3.3 0.00038815999999999997 0 0.00038808 0 0.00038818 3.3 0.0003881 3.3 0.0003882 0 0.00038812 0 0.00038822 3.3 0.00038814 3.3 0.00038824 0 0.00038815999999999997 0 0.00038825999999999997 3.3 0.00038818 3.3 0.00038828 0 0.0003882 0 0.0003883 3.3 0.00038822 3.3 0.00038832 0 0.00038824 0 0.00038834 3.3 0.00038825999999999997 3.3 0.00038836 0 0.00038828 0 0.00038838 3.3 0.0003883 3.3 0.0003884 0 0.00038832 0 0.00038842 3.3 0.00038834 3.3 0.00038844 0 0.00038836 0 0.00038846 3.3 0.00038837999999999996 3.3 0.00038847999999999997 0 0.0003884 0 0.0003885 3.3 0.00038842 3.3 0.00038852 0 0.00038844 0 0.00038854 3.3 0.00038846 3.3 0.00038856 0 0.00038847999999999997 0 0.00038857999999999997 3.3 0.0003885 3.3 0.0003886 0 0.00038852 0 0.00038862 3.3 0.00038854 3.3 0.00038864 0 0.00038856 0 0.00038866 3.3 0.00038857999999999997 3.3 0.00038867999999999997 0 0.0003886 0 0.0003887 3.3 0.00038862 3.3 0.00038872 0 0.00038864 0 0.00038874 3.3 0.00038866 3.3 0.00038876 0 0.00038867999999999997 0 0.00038878 3.3 0.0003887 3.3 0.0003888 0 0.00038872 0 0.00038882 3.3 0.00038874 3.3 0.00038884 0 0.00038876 0 0.00038886 3.3 0.00038878 3.3 0.00038888 0 0.00038879999999999996 0 0.00038889999999999997 3.3 0.00038882 3.3 0.00038892 0 0.00038884 0 0.00038894 3.3 0.00038886 3.3 0.00038896 0 0.00038888 0 0.00038898 3.3 0.00038889999999999997 3.3 0.00038899999999999997 0 0.00038892 0 0.00038902 3.3 0.00038894 3.3 0.00038904 0 0.00038896 0 0.00038906 3.3 0.00038898 3.3 0.00038908 0 0.00038899999999999997 0 0.00038909999999999997 3.3 0.00038902 3.3 0.00038912 0 0.00038904 0 0.00038914 3.3 0.00038906 3.3 0.00038916 0 0.00038908 0 0.00038918 3.3 0.00038909999999999997 3.3 0.0003892 0 0.00038912 0 0.00038922 3.3 0.00038914 3.3 0.00038924 0 0.00038916 0 0.00038926 3.3 0.00038918 3.3 0.00038928 0 0.0003892 0 0.0003893 3.3 0.00038921999999999996 3.3 0.00038931999999999997 0 0.00038924 0 0.00038934 3.3 0.00038926 3.3 0.00038936 0 0.00038928 0 0.00038938 3.3 0.0003893 3.3 0.0003894 0 0.00038931999999999997 0 0.00038941999999999997 3.3 0.00038934 3.3 0.00038944 0 0.00038936 0 0.00038946 3.3 0.00038938 3.3 0.00038948 0 0.0003894 0 0.0003895 3.3 0.00038941999999999997 3.3 0.00038951999999999997 0 0.00038944 0 0.00038954 3.3 0.00038946 3.3 0.00038956 0 0.00038948 0 0.00038958 3.3 0.0003895 3.3 0.0003896 0 0.00038951999999999997 0 0.00038961999999999997 3.3 0.00038954 3.3 0.00038964 0 0.00038956 0 0.00038966 3.3 0.00038958 3.3 0.00038968 0 0.0003896 0 0.0003897 3.3 0.00038961999999999997 3.3 0.00038972 0 0.00038964 0 0.00038974 3.3 0.00038966 3.3 0.00038976 0 0.00038968 0 0.00038978 3.3 0.0003897 3.3 0.0003898 0 0.00038972 0 0.00038982 3.3 0.00038973999999999996 3.3 0.00038983999999999997 0 0.00038976 0 0.00038986 3.3 0.00038978 3.3 0.00038988 0 0.0003898 0 0.0003899 3.3 0.00038982 3.3 0.00038992 0 0.00038983999999999997 0 0.00038993999999999997 3.3 0.00038986 3.3 0.00038996 0 0.00038988 0 0.00038998 3.3 0.0003899 3.3 0.00039 0 0.00038992 0 0.00039002 3.3 0.00038993999999999997 3.3 0.00039003999999999997 0 0.00038996 0 0.00039006 3.3 0.00038998 3.3 0.00039008 0 0.00039 0 0.0003901 3.3 0.00039002 3.3 0.00039012 0 0.00039003999999999997 0 0.00039014 3.3 0.00039006 3.3 0.00039016 0 0.00039008 0 0.00039018 3.3 0.0003901 3.3 0.0003902 0 0.00039012 0 0.00039022 3.3 0.00039014 3.3 0.00039024 0 0.00039015999999999996 0 0.00039025999999999997 3.3 0.00039018 3.3 0.00039028 0 0.0003902 0 0.0003903 3.3 0.00039022 3.3 0.00039032 0 0.00039024 0 0.00039034 3.3 0.00039025999999999997 3.3 0.00039035999999999997 0 0.00039028 0 0.00039038 3.3 0.0003903 3.3 0.0003904 0 0.00039032 0 0.00039042 3.3 0.00039034 3.3 0.00039044 0 0.00039035999999999997 0 0.00039045999999999997 3.3 0.00039038 3.3 0.00039048 0 0.0003904 0 0.0003905 3.3 0.00039042 3.3 0.00039052 0 0.00039044 0 0.00039054 3.3 0.00039045999999999997 3.3 0.00039056 0 0.00039048 0 0.00039058 3.3 0.0003905 3.3 0.0003906 0 0.00039052 0 0.00039062 3.3 0.00039054 3.3 0.00039064 0 0.00039056 0 0.00039066 3.3 0.00039057999999999996 3.3 0.00039067999999999997 0 0.0003906 0 0.0003907 3.3 0.00039062 3.3 0.00039072 0 0.00039064 0 0.00039074 3.3 0.00039066 3.3 0.00039076 0 0.00039067999999999997 0 0.00039077999999999997 3.3 0.0003907 3.3 0.0003908 0 0.00039072 0 0.00039082 3.3 0.00039074 3.3 0.00039084 0 0.00039076 0 0.00039086 3.3 0.00039077999999999997 3.3 0.00039087999999999997 0 0.0003908 0 0.0003909 3.3 0.00039082 3.3 0.00039092 0 0.00039084 0 0.00039094 3.3 0.00039086 3.3 0.00039096 0 0.00039087999999999997 0 0.00039098 3.3 0.0003909 3.3 0.000391 0 0.00039092 0 0.00039102 3.3 0.00039094 3.3 0.00039104 0 0.00039096 0 0.00039106 3.3 0.00039098 3.3 0.00039108 0 0.00039099999999999996 0 0.00039109999999999997 3.3 0.00039102 3.3 0.00039112 0 0.00039104 0 0.00039114 3.3 0.00039106 3.3 0.00039116 0 0.00039108 0 0.00039118 3.3 0.00039109999999999997 3.3 0.00039119999999999997 0 0.00039112 0 0.00039122 3.3 0.00039114 3.3 0.00039124 0 0.00039116 0 0.00039126 3.3 0.00039118 3.3 0.00039128 0 0.00039119999999999997 0 0.00039129999999999997 3.3 0.00039122 3.3 0.00039132 0 0.00039124 0 0.00039134 3.3 0.00039126 3.3 0.00039136 0 0.00039128 0 0.00039138 3.3 0.00039129999999999997 3.3 0.00039139999999999997 0 0.00039132 0 0.00039142 3.3 0.00039134 3.3 0.00039144 0 0.00039136 0 0.00039146 3.3 0.00039138 3.3 0.00039148 0 0.00039139999999999997 0 0.0003915 3.3 0.00039142 3.3 0.00039152 0 0.00039144 0 0.00039154 3.3 0.00039146 3.3 0.00039156 0 0.00039148 0 0.00039158 3.3 0.0003915 3.3 0.0003916 0 0.00039151999999999996 0 0.00039161999999999997 3.3 0.00039154 3.3 0.00039164 0 0.00039156 0 0.00039166 3.3 0.00039158 3.3 0.00039168 0 0.0003916 0 0.0003917 3.3 0.00039161999999999997 3.3 0.00039171999999999997 0 0.00039164 0 0.00039174 3.3 0.00039166 3.3 0.00039176 0 0.00039168 0 0.00039178 3.3 0.0003917 3.3 0.0003918 0 0.00039171999999999997 0 0.00039181999999999997 3.3 0.00039174 3.3 0.00039184 0 0.00039176 0 0.00039186 3.3 0.00039178 3.3 0.00039188 0 0.0003918 0 0.0003919 3.3 0.00039181999999999997 3.3 0.00039192 0 0.00039184 0 0.00039194 3.3 0.00039186 3.3 0.00039196 0 0.00039188 0 0.00039198 3.3 0.0003919 3.3 0.000392 0 0.00039192 0 0.00039202 3.3 0.00039193999999999996 3.3 0.00039203999999999997 0 0.00039196 0 0.00039206 3.3 0.00039198 3.3 0.00039208 0 0.000392 0 0.0003921 3.3 0.00039202 3.3 0.00039212 0 0.00039203999999999997 0 0.00039213999999999997 3.3 0.00039206 3.3 0.00039216 0 0.00039208 0 0.00039218 3.3 0.0003921 3.3 0.0003922 0 0.00039212 0 0.00039222 3.3 0.00039213999999999997 3.3 0.00039223999999999997 0 0.00039216 0 0.00039226 3.3 0.00039218 3.3 0.00039228 0 0.0003922 0 0.0003923 3.3 0.00039222 3.3 0.00039232 0 0.00039223999999999997 0 0.00039234 3.3 0.00039226 3.3 0.00039236 0 0.00039228 0 0.00039238 3.3 0.0003923 3.3 0.0003924 0 0.00039232 0 0.00039242 3.3 0.00039234 3.3 0.00039244 0 0.00039235999999999996 0 0.00039245999999999997 3.3 0.00039238 3.3 0.00039248 0 0.0003924 0 0.0003925 3.3 0.00039242 3.3 0.00039252 0 0.00039244 0 0.00039254 3.3 0.00039245999999999997 3.3 0.00039255999999999997 0 0.00039248 0 0.00039258 3.3 0.0003925 3.3 0.0003926 0 0.00039252 0 0.00039262 3.3 0.00039254 3.3 0.00039264 0 0.00039255999999999997 0 0.00039265999999999997 3.3 0.00039258 3.3 0.00039268 0 0.0003926 0 0.0003927 3.3 0.00039262 3.3 0.00039272 0 0.00039264 0 0.00039274 3.3 0.00039265999999999997 3.3 0.00039276 0 0.00039268 0 0.00039278 3.3 0.0003927 3.3 0.0003928 0 0.00039272 0 0.00039282 3.3 0.00039274 3.3 0.00039284 0 0.00039276 0 0.00039286 3.3 0.00039277999999999996 3.3 0.00039287999999999997 0 0.0003928 0 0.0003929 3.3 0.00039282 3.3 0.00039292 0 0.00039284 0 0.00039294 3.3 0.00039286 3.3 0.00039296 0 0.00039287999999999997 0 0.00039297999999999997 3.3 0.0003929 3.3 0.000393 0 0.00039292 0 0.00039302 3.3 0.00039294 3.3 0.00039304 0 0.00039296 0 0.00039306 3.3 0.00039297999999999997 3.3 0.00039307999999999997 0 0.000393 0 0.0003931 3.3 0.00039302 3.3 0.00039312 0 0.00039304 0 0.00039314 3.3 0.00039306 3.3 0.00039316 0 0.00039307999999999997 0 0.00039317999999999997 3.3 0.0003931 3.3 0.0003932 0 0.00039312 0 0.00039322 3.3 0.00039314 3.3 0.00039324 0 0.00039316 0 0.00039326 3.3 0.00039317999999999997 3.3 0.00039328 0 0.0003932 0 0.0003933 3.3 0.00039322 3.3 0.00039332 0 0.00039324 0 0.00039334 3.3 0.00039326 3.3 0.00039336 0 0.00039328 0 0.00039338 3.3 0.00039329999999999996 3.3 0.00039339999999999997 0 0.00039332 0 0.00039342 3.3 0.00039334 3.3 0.00039344 0 0.00039336 0 0.00039346 3.3 0.00039338 3.3 0.00039348 0 0.00039339999999999997 0 0.00039349999999999997 3.3 0.00039342 3.3 0.00039352 0 0.00039344 0 0.00039354 3.3 0.00039346 3.3 0.00039356 0 0.00039348 0 0.00039358 3.3 0.00039349999999999997 3.3 0.00039359999999999997 0 0.00039352 0 0.00039362 3.3 0.00039354 3.3 0.00039364 0 0.00039356 0 0.00039366 3.3 0.00039358 3.3 0.00039368 0 0.00039359999999999997 0 0.0003937 3.3 0.00039362 3.3 0.00039372 0 0.00039364 0 0.00039374 3.3 0.00039366 3.3 0.00039376 0 0.00039368 0 0.00039378 3.3 0.0003937 3.3 0.0003938 0 0.00039371999999999996 0 0.00039381999999999997 3.3 0.00039374 3.3 0.00039384 0 0.00039376 0 0.00039386 3.3 0.00039378 3.3 0.00039388 0 0.0003938 0 0.0003939 3.3 0.00039381999999999997 3.3 0.00039391999999999997 0 0.00039384 0 0.00039394 3.3 0.00039386 3.3 0.00039396 0 0.00039388 0 0.00039398 3.3 0.0003939 3.3 0.000394 0 0.00039391999999999997 0 0.00039401999999999997 3.3 0.00039394 3.3 0.00039404 0 0.00039396 0 0.00039406 3.3 0.00039398 3.3 0.00039408 0 0.000394 0 0.0003941 3.3 0.00039401999999999997 3.3 0.00039412 0 0.00039404 0 0.00039414 3.3 0.00039406 3.3 0.00039416 0 0.00039408 0 0.00039418 3.3 0.0003941 3.3 0.0003942 0 0.00039412 0 0.00039422 3.3 0.00039413999999999996 3.3 0.00039423999999999997 0 0.00039416 0 0.00039426 3.3 0.00039418 3.3 0.00039428 0 0.0003942 0 0.0003943 3.3 0.00039422 3.3 0.00039432 0 0.00039423999999999997 0 0.00039433999999999997 3.3 0.00039426 3.3 0.00039436 0 0.00039428 0 0.00039438 3.3 0.0003943 3.3 0.0003944 0 0.00039432 0 0.00039442 3.3 0.00039433999999999997 3.3 0.00039443999999999997 0 0.00039436 0 0.00039446 3.3 0.00039438 3.3 0.00039448 0 0.0003944 0 0.0003945 3.3 0.00039442 3.3 0.00039452 0 0.00039443999999999997 0 0.00039454 3.3 0.00039446 3.3 0.00039456 0 0.00039448 0 0.00039458 3.3 0.0003945 3.3 0.0003946 0 0.00039452 0 0.00039462 3.3 0.00039454 3.3 0.00039464 0 0.00039455999999999996 0 0.00039465999999999997 3.3 0.00039458 3.3 0.00039468 0 0.0003946 0 0.0003947 3.3 0.00039462 3.3 0.00039472 0 0.00039464 0 0.00039474 3.3 0.00039465999999999997 3.3 0.00039475999999999997 0 0.00039468 0 0.00039478 3.3 0.0003947 3.3 0.0003948 0 0.00039472 0 0.00039482 3.3 0.00039474 3.3 0.00039484 0 0.00039475999999999997 0 0.00039485999999999997 3.3 0.00039478 3.3 0.00039488 0 0.0003948 0 0.0003949 3.3 0.00039482 3.3 0.00039492 0 0.00039484 0 0.00039494 3.3 0.00039485999999999997 3.3 0.00039495999999999997 0 0.00039488 0 0.00039498 3.3 0.0003949 3.3 0.000395 0 0.00039492 0 0.00039502 3.3 0.00039494 3.3 0.00039504 0 0.00039495999999999997 0 0.00039506 3.3 0.00039498 3.3 0.00039508 0 0.000395 0 0.0003951 3.3 0.00039502 3.3 0.00039512 0 0.00039504 0 0.00039514 3.3 0.00039506 3.3 0.00039516 0 0.00039507999999999996 0 0.00039517999999999997 3.3 0.0003951 3.3 0.0003952 0 0.00039512 0 0.00039522 3.3 0.00039514 3.3 0.00039524 0 0.00039516 0 0.00039526 3.3 0.00039517999999999997 3.3 0.00039527999999999997 0 0.0003952 0 0.0003953 3.3 0.00039522 3.3 0.00039532 0 0.00039524 0 0.00039534 3.3 0.00039526 3.3 0.00039536 0 0.00039527999999999997 0 0.00039537999999999997 3.3 0.0003953 3.3 0.0003954 0 0.00039532 0 0.00039542 3.3 0.00039534 3.3 0.00039544 0 0.00039536 0 0.00039546 3.3 0.00039537999999999997 3.3 0.00039548 0 0.0003954 0 0.0003955 3.3 0.00039542 3.3 0.00039552 0 0.00039544 0 0.00039554 3.3 0.00039546 3.3 0.00039556 0 0.00039548 0 0.00039558 3.3 0.00039549999999999996 3.3 0.00039559999999999997 0 0.00039552 0 0.00039562 3.3 0.00039554 3.3 0.00039564 0 0.00039556 0 0.00039566 3.3 0.00039558 3.3 0.00039568 0 0.00039559999999999997 0 0.00039569999999999997 3.3 0.00039562 3.3 0.00039572 0 0.00039564 0 0.00039574 3.3 0.00039566 3.3 0.00039576 0 0.00039568 0 0.00039578 3.3 0.00039569999999999997 3.3 0.00039579999999999997 0 0.00039572 0 0.00039582 3.3 0.00039574 3.3 0.00039584 0 0.00039576 0 0.00039586 3.3 0.00039578 3.3 0.00039588 0 0.00039579999999999997 0 0.0003959 3.3 0.00039582 3.3 0.00039592 0 0.00039584 0 0.00039594 3.3 0.00039586 3.3 0.00039596 0 0.00039588 0 0.00039598 3.3 0.0003959 3.3 0.000396 0 0.00039591999999999996 0 0.00039601999999999997 3.3 0.00039594 3.3 0.00039604 0 0.00039596 0 0.00039606 3.3 0.00039598 3.3 0.00039608 0 0.000396 0 0.0003961 3.3 0.00039601999999999997 3.3 0.00039611999999999997 0 0.00039604 0 0.00039614 3.3 0.00039606 3.3 0.00039616 0 0.00039608 0 0.00039618 3.3 0.0003961 3.3 0.0003962 0 0.00039611999999999997 0 0.00039621999999999997 3.3 0.00039614 3.3 0.00039624 0 0.00039616 0 0.00039626 3.3 0.00039618 3.3 0.00039628 0 0.0003962 0 0.0003963 3.3 0.00039621999999999997 3.3 0.00039632 0 0.00039624 0 0.00039634 3.3 0.00039626 3.3 0.00039636 0 0.00039628 0 0.00039638 3.3 0.0003963 3.3 0.0003964 0 0.00039632 0 0.00039642 3.3 0.00039633999999999996 3.3 0.00039643999999999997 0 0.00039636 0 0.00039646 3.3 0.00039638 3.3 0.00039648 0 0.0003964 0 0.0003965 3.3 0.00039642 3.3 0.00039652 0 0.00039643999999999997 0 0.00039653999999999997 3.3 0.00039646 3.3 0.00039656 0 0.00039648 0 0.00039658 3.3 0.0003965 3.3 0.0003966 0 0.00039652 0 0.00039662 3.3 0.00039653999999999997 3.3 0.00039663999999999997 0 0.00039656 0 0.00039666 3.3 0.00039658 3.3 0.00039668 0 0.0003966 0 0.0003967 3.3 0.00039662 3.3 0.00039672 0 0.00039663999999999997 0 0.00039673999999999997 3.3 0.00039666 3.3 0.00039676 0 0.00039668 0 0.00039678 3.3 0.0003967 3.3 0.0003968 0 0.00039672 0 0.00039682 3.3 0.00039673999999999997 3.3 0.00039684 0 0.00039676 0 0.00039686 3.3 0.00039678 3.3 0.00039688 0 0.0003968 0 0.0003969 3.3 0.00039682 3.3 0.00039692 0 0.00039684 0 0.00039694 3.3 0.00039685999999999996 3.3 0.00039695999999999997 0 0.00039688 0 0.00039698 3.3 0.0003969 3.3 0.000397 0 0.00039692 0 0.00039702 3.3 0.00039694 3.3 0.00039704 0 0.00039695999999999997 0 0.00039705999999999997 3.3 0.00039698 3.3 0.00039708 0 0.000397 0 0.0003971 3.3 0.00039702 3.3 0.00039712 0 0.00039704 0 0.00039714 3.3 0.00039705999999999997 3.3 0.00039715999999999997 0 0.00039708 0 0.00039718 3.3 0.0003971 3.3 0.0003972 0 0.00039712 0 0.00039722 3.3 0.00039714 3.3 0.00039724 0 0.00039715999999999997 0 0.00039726 3.3 0.00039718 3.3 0.00039728 0 0.0003972 0 0.0003973 3.3 0.00039722 3.3 0.00039732 0 0.00039724 0 0.00039734 3.3 0.00039726 3.3 0.00039736 0 0.00039727999999999996 0 0.00039737999999999997 3.3 0.0003973 3.3 0.0003974 0 0.00039732 0 0.00039742 3.3 0.00039734 3.3 0.00039744 0 0.00039736 0 0.00039746 3.3 0.00039737999999999997 3.3 0.00039747999999999997 0 0.0003974 0 0.0003975 3.3 0.00039742 3.3 0.00039752 0 0.00039744 0 0.00039754 3.3 0.00039746 3.3 0.00039756 0 0.00039747999999999997 0 0.00039757999999999997 3.3 0.0003975 3.3 0.0003976 0 0.00039752 0 0.00039762 3.3 0.00039754 3.3 0.00039764 0 0.00039756 0 0.00039766 3.3 0.00039757999999999997 3.3 0.00039768 0 0.0003976 0 0.0003977 3.3 0.00039762 3.3 0.00039772 0 0.00039764 0 0.00039774 3.3 0.00039766 3.3 0.00039776 0 0.00039768 0 0.00039778 3.3 0.00039769999999999996 3.3 0.00039779999999999997 0 0.00039772 0 0.00039782 3.3 0.00039774 3.3 0.00039784 0 0.00039776 0 0.00039786 3.3 0.00039778 3.3 0.00039788 0 0.00039779999999999997 0 0.00039789999999999997 3.3 0.00039782 3.3 0.00039792 0 0.00039784 0 0.00039794 3.3 0.00039786 3.3 0.00039796 0 0.00039788 0 0.00039798 3.3 0.00039789999999999997 3.3 0.00039799999999999997 0 0.00039792 0 0.00039802 3.3 0.00039794 3.3 0.00039804 0 0.00039796 0 0.00039806 3.3 0.00039798 3.3 0.00039808 0 0.00039799999999999997 0 0.0003981 3.3 0.00039802 3.3 0.00039812 0 0.00039804 0 0.00039814 3.3 0.00039806 3.3 0.00039816 0 0.00039808 0 0.00039818 3.3 0.0003981 3.3 0.0003982 0 0.00039811999999999996 0 0.00039821999999999997 3.3 0.00039814 3.3 0.00039824 0 0.00039816 0 0.00039826 3.3 0.00039818 3.3 0.00039828 0 0.0003982 0 0.0003983 3.3 0.00039821999999999997 3.3 0.00039831999999999997 0 0.00039824 0 0.00039834 3.3 0.00039826 3.3 0.00039836 0 0.00039828 0 0.00039838 3.3 0.0003983 3.3 0.0003984 0 0.00039831999999999997 0 0.00039841999999999997 3.3 0.00039834 3.3 0.00039844 0 0.00039836 0 0.00039846 3.3 0.00039838 3.3 0.00039848 0 0.0003984 0 0.0003985 3.3 0.00039841999999999997 3.3 0.00039851999999999997 0 0.00039844 0 0.00039854 3.3 0.00039846 3.3 0.00039856 0 0.00039848 0 0.00039858 3.3 0.0003985 3.3 0.0003986 0 0.00039851999999999997 0 0.00039862 3.3 0.00039854 3.3 0.00039864 0 0.00039856 0 0.00039866 3.3 0.00039858 3.3 0.00039868 0 0.0003986 0 0.0003987 3.3 0.00039862 3.3 0.00039872 0 0.00039863999999999996 0 0.00039873999999999997 3.3 0.00039866 3.3 0.00039876 0 0.00039868 0 0.00039878 3.3 0.0003987 3.3 0.0003988 0 0.00039872 0 0.00039882 3.3 0.00039873999999999997 3.3 0.00039883999999999997 0 0.00039876 0 0.00039886 3.3 0.00039878 3.3 0.00039888 0 0.0003988 0 0.0003989 3.3 0.00039882 3.3 0.00039892 0 0.00039883999999999997 0 0.00039893999999999997 3.3 0.00039886 3.3 0.00039896 0 0.00039888 0 0.00039898 3.3 0.0003989 3.3 0.000399 0 0.00039892 0 0.00039902 3.3 0.00039893999999999997 3.3 0.00039904 0 0.00039896 0 0.00039906 3.3 0.00039898 3.3 0.00039908 0 0.000399 0 0.0003991 3.3 0.00039902 3.3 0.00039912 0 0.00039904 0 0.00039914 3.3 0.00039905999999999996 3.3 0.00039915999999999997 0 0.00039908 0 0.00039918 3.3 0.0003991 3.3 0.0003992 0 0.00039912 0 0.00039922 3.3 0.00039914 3.3 0.00039924 0 0.00039915999999999997 0 0.00039925999999999997 3.3 0.00039918 3.3 0.00039928 0 0.0003992 0 0.0003993 3.3 0.00039922 3.3 0.00039932 0 0.00039924 0 0.00039934 3.3 0.00039925999999999997 3.3 0.00039935999999999997 0 0.00039928 0 0.00039938 3.3 0.0003993 3.3 0.0003994 0 0.00039932 0 0.00039942 3.3 0.00039934 3.3 0.00039944 0 0.00039935999999999997 0 0.00039946 3.3 0.00039938 3.3 0.00039948 0 0.0003994 0 0.0003995 3.3 0.00039942 3.3 0.00039952 0 0.00039944 0 0.00039954 3.3 0.00039946 3.3 0.00039956 0 0.00039947999999999996 0 0.00039957999999999997 3.3 0.0003995 3.3 0.0003996 0 0.00039952 0 0.00039962 3.3 0.00039954 3.3 0.00039964 0 0.00039956 0 0.00039966 3.3 0.00039957999999999997 3.3 0.00039967999999999997 0 0.0003996 0 0.0003997 3.3 0.00039962 3.3 0.00039972 0 0.00039964 0 0.00039974 3.3 0.00039966 3.3 0.00039976 0 0.00039967999999999997 0 0.00039977999999999997 3.3 0.0003997 3.3 0.0003998 0 0.00039972 0 0.00039982 3.3 0.00039974 3.3 0.00039984 0 0.00039976 0 0.00039986 3.3 0.00039977999999999997 3.3 0.00039987999999999997 0 0.0003998 0 0.0003999 3.3 0.00039982 3.3 0.00039992 0 0.00039984 0 0.00039994 3.3 0.00039986 3.3 0.00039996 0 0.00039987999999999997 0 0.00039998 3.3 0.00039989999999999996 3.3 0.00039999999999999996 0 0.00039992 0 0.00040002 3.3 0.00039994 3.3 0.00040004 0 0.00039996 0 0.00040006 3.3 0.00039998 3.3 0.00040008 0 0.00039999999999999996 0 0.00040009999999999997 3.3 0.00040002 3.3 0.00040012 0 0.00040004 0 0.00040014 3.3 0.00040006 3.3 0.00040016 0 0.00040008 0 0.00040018 3.3 0.00040009999999999997 3.3 0.00040019999999999997 0 0.00040012 0 0.00040022 3.3 0.00040014 3.3 0.00040024 0 0.00040016 0 0.00040026 3.3 0.00040018 3.3 0.00040028 0 0.00040019999999999997 0 0.00040029999999999997 3.3 0.00040022 3.3 0.00040032 0 0.00040024 0 0.00040034 3.3 0.00040026 3.3 0.00040036 0 0.00040028 0 0.00040038 3.3 0.00040029999999999997 3.3 0.0004004 0 0.00040032 0 0.00040042 3.3 0.00040034 3.3 0.00040044 0 0.00040036 0 0.00040046 3.3 0.00040038 3.3 0.00040048 0 0.0004004 0 0.0004005 3.3 0.00040041999999999996 3.3 0.00040051999999999997 0 0.00040044 0 0.00040054 3.3 0.00040046 3.3 0.00040056 0 0.00040048 0 0.00040058 3.3 0.0004005 3.3 0.0004006 0 0.00040051999999999997 0 0.00040061999999999997 3.3 0.00040054 3.3 0.00040064 0 0.00040056 0 0.00040066 3.3 0.00040058 3.3 0.00040068 0 0.0004006 0 0.0004007 3.3 0.00040061999999999997 3.3 0.00040071999999999997 0 0.00040064 0 0.00040074 3.3 0.00040066 3.3 0.00040076 0 0.00040068 0 0.00040078 3.3 0.0004007 3.3 0.0004008 0 0.00040071999999999997 0 0.00040082 3.3 0.00040074 3.3 0.00040084 0 0.00040076 0 0.00040086 3.3 0.00040078 3.3 0.00040088 0 0.0004008 0 0.0004009 3.3 0.00040082 3.3 0.00040092 0 0.00040083999999999996 0 0.00040093999999999997 3.3 0.00040086 3.3 0.00040096 0 0.00040088 0 0.00040098 3.3 0.0004009 3.3 0.000401 0 0.00040092 0 0.00040102 3.3 0.00040093999999999997 3.3 0.00040103999999999997 0 0.00040096 0 0.00040106 3.3 0.00040098 3.3 0.00040108 0 0.000401 0 0.0004011 3.3 0.00040102 3.3 0.00040112 0 0.00040103999999999997 0 0.00040113999999999997 3.3 0.00040106 3.3 0.00040116 0 0.00040108 0 0.00040118 3.3 0.0004011 3.3 0.0004012 0 0.00040112 0 0.00040122 3.3 0.00040113999999999997 3.3 0.00040124 0 0.00040116 0 0.00040126 3.3 0.00040118 3.3 0.00040128 0 0.0004012 0 0.0004013 3.3 0.00040122 3.3 0.00040132 0 0.00040124 0 0.00040134 3.3 0.00040125999999999996 3.3 0.00040135999999999997 0 0.00040128 0 0.00040138 3.3 0.0004013 3.3 0.0004014 0 0.00040132 0 0.00040142 3.3 0.00040134 3.3 0.00040144 0 0.00040135999999999997 0 0.00040145999999999997 3.3 0.00040138 3.3 0.00040148 0 0.0004014 0 0.0004015 3.3 0.00040142 3.3 0.00040152 0 0.00040144 0 0.00040154 3.3 0.00040145999999999997 3.3 0.00040155999999999997 0 0.00040148 0 0.00040158 3.3 0.0004015 3.3 0.0004016 0 0.00040152 0 0.00040162 3.3 0.00040154 3.3 0.00040164 0 0.00040155999999999997 0 0.00040165999999999997 3.3 0.00040158 3.3 0.00040168 0 0.0004016 0 0.0004017 3.3 0.00040162 3.3 0.00040172 0 0.00040164 0 0.00040174 3.3 0.00040165999999999997 3.3 0.00040176 0 0.00040167999999999996 0 0.00040177999999999996 3.3 0.0004017 3.3 0.0004018 0 0.00040172 0 0.00040182 3.3 0.00040174 3.3 0.00040184 0 0.00040176 0 0.00040186 3.3 0.00040177999999999996 3.3 0.00040187999999999997 0 0.0004018 0 0.0004019 3.3 0.00040182 3.3 0.00040192 0 0.00040184 0 0.00040194 3.3 0.00040186 3.3 0.00040196 0 0.00040187999999999997 0 0.00040197999999999997 3.3 0.0004019 3.3 0.000402 0 0.00040192 0 0.00040202 3.3 0.00040194 3.3 0.00040204 0 0.00040196 0 0.00040206 3.3 0.00040197999999999997 3.3 0.00040207999999999997 0 0.000402 0 0.0004021 3.3 0.00040202 3.3 0.00040212 0 0.00040204 0 0.00040214 3.3 0.00040206 3.3 0.00040216 0 0.00040207999999999997 0 0.00040218 3.3 0.0004021 3.3 0.0004022 0 0.00040212 0 0.00040222 3.3 0.00040214 3.3 0.00040224 0 0.00040216 0 0.00040226 3.3 0.00040218 3.3 0.00040228 0 0.00040219999999999996 0 0.00040229999999999997 3.3 0.00040222 3.3 0.00040232 0 0.00040224 0 0.00040234 3.3 0.00040226 3.3 0.00040236 0 0.00040228 0 0.00040238 3.3 0.00040229999999999997 3.3 0.00040239999999999997 0 0.00040232 0 0.00040242 3.3 0.00040234 3.3 0.00040244 0 0.00040236 0 0.00040246 3.3 0.00040238 3.3 0.00040248 0 0.00040239999999999997 0 0.00040249999999999997 3.3 0.00040242 3.3 0.00040252 0 0.00040244 0 0.00040254 3.3 0.00040246 3.3 0.00040256 0 0.00040248 0 0.00040258 3.3 0.00040249999999999997 3.3 0.0004026 0 0.00040252 0 0.00040262 3.3 0.00040254 3.3 0.00040264 0 0.00040256 0 0.00040266 3.3 0.00040258 3.3 0.00040268 0 0.0004026 0 0.0004027 3.3 0.00040261999999999996 3.3 0.00040271999999999997 0 0.00040264 0 0.00040274 3.3 0.00040266 3.3 0.00040276 0 0.00040268 0 0.00040278 3.3 0.0004027 3.3 0.0004028 0 0.00040271999999999997 0 0.00040281999999999997 3.3 0.00040274 3.3 0.00040284 0 0.00040276 0 0.00040286 3.3 0.00040278 3.3 0.00040288 0 0.0004028 0 0.0004029 3.3 0.00040281999999999997 3.3 0.00040291999999999997 0 0.00040284 0 0.00040294 3.3 0.00040286 3.3 0.00040296 0 0.00040288 0 0.00040298 3.3 0.0004029 3.3 0.000403 0 0.00040291999999999997 0 0.00040302 3.3 0.00040294 3.3 0.00040304 0 0.00040296 0 0.00040306 3.3 0.00040298 3.3 0.00040308 0 0.000403 0 0.0004031 3.3 0.00040302 3.3 0.00040312 0 0.00040303999999999996 0 0.00040313999999999997 3.3 0.00040306 3.3 0.00040316 0 0.00040308 0 0.00040318 3.3 0.0004031 3.3 0.0004032 0 0.00040312 0 0.00040322 3.3 0.00040313999999999997 3.3 0.00040323999999999997 0 0.00040316 0 0.00040326 3.3 0.00040318 3.3 0.00040328 0 0.0004032 0 0.0004033 3.3 0.00040322 3.3 0.00040332 0 0.00040323999999999997 0 0.00040333999999999997 3.3 0.00040326 3.3 0.00040336 0 0.00040328 0 0.00040338 3.3 0.0004033 3.3 0.0004034 0 0.00040332 0 0.00040342 3.3 0.00040333999999999997 3.3 0.00040343999999999997 0 0.00040336 0 0.00040346 3.3 0.00040338 3.3 0.00040348 0 0.0004034 0 0.0004035 3.3 0.00040342 3.3 0.00040352 0 0.00040343999999999997 0 0.00040354 3.3 0.00040346 3.3 0.00040356 0 0.00040348 0 0.00040358 3.3 0.0004035 3.3 0.0004036 0 0.00040352 0 0.00040362 3.3 0.00040354 3.3 0.00040364 0 0.00040355999999999996 0 0.00040365999999999997 3.3 0.00040358 3.3 0.00040368 0 0.0004036 0 0.0004037 3.3 0.00040362 3.3 0.00040372 0 0.00040364 0 0.00040374 3.3 0.00040365999999999997 3.3 0.00040375999999999997 0 0.00040368 0 0.00040378 3.3 0.0004037 3.3 0.0004038 0 0.00040372 0 0.00040382 3.3 0.00040374 3.3 0.00040384 0 0.00040375999999999997 0 0.00040385999999999997 3.3 0.00040378 3.3 0.00040388 0 0.0004038 0 0.0004039 3.3 0.00040382 3.3 0.00040392 0 0.00040384 0 0.00040394 3.3 0.00040385999999999997 3.3 0.00040396 0 0.00040388 0 0.00040398 3.3 0.0004039 3.3 0.000404 0 0.00040392 0 0.00040402 3.3 0.00040394 3.3 0.00040404 0 0.00040396 0 0.00040406 3.3 0.00040397999999999996 3.3 0.00040407999999999997 0 0.000404 0 0.0004041 3.3 0.00040402 3.3 0.00040412 0 0.00040404 0 0.00040414 3.3 0.00040406 3.3 0.00040416 0 0.00040407999999999997 0 0.00040417999999999997 3.3 0.0004041 3.3 0.0004042 0 0.00040412 0 0.00040422 3.3 0.00040414 3.3 0.00040424 0 0.00040416 0 0.00040426 3.3 0.00040417999999999997 3.3 0.00040427999999999997 0 0.0004042 0 0.0004043 3.3 0.00040422 3.3 0.00040432 0 0.00040424 0 0.00040434 3.3 0.00040426 3.3 0.00040436 0 0.00040427999999999997 0 0.00040438 3.3 0.0004043 3.3 0.0004044 0 0.00040432 0 0.00040442 3.3 0.00040434 3.3 0.00040444 0 0.00040436 0 0.00040446 3.3 0.00040438 3.3 0.00040448 0 0.00040439999999999996 0 0.00040449999999999997 3.3 0.00040442 3.3 0.00040452 0 0.00040444 0 0.00040454 3.3 0.00040446 3.3 0.00040456 0 0.00040448 0 0.00040458 3.3 0.00040449999999999997 3.3 0.00040459999999999997 0 0.00040452 0 0.00040462 3.3 0.00040454 3.3 0.00040464 0 0.00040456 0 0.00040466 3.3 0.00040458 3.3 0.00040468 0 0.00040459999999999997 0 0.00040469999999999997 3.3 0.00040462 3.3 0.00040472 0 0.00040464 0 0.00040474 3.3 0.00040466 3.3 0.00040476 0 0.00040468 0 0.00040478 3.3 0.00040469999999999997 3.3 0.0004048 0 0.00040472 0 0.00040482 3.3 0.00040474 3.3 0.00040484 0 0.00040476 0 0.00040486 3.3 0.00040478 3.3 0.00040488 0 0.0004048 0 0.0004049 3.3 0.00040481999999999996 3.3 0.00040491999999999997 0 0.00040484 0 0.00040494 3.3 0.00040486 3.3 0.00040496 0 0.00040488 0 0.00040498 3.3 0.0004049 3.3 0.000405 0 0.00040491999999999997 0 0.00040501999999999997 3.3 0.00040494 3.3 0.00040504 0 0.00040496 0 0.00040506 3.3 0.00040498 3.3 0.00040508 0 0.000405 0 0.0004051 3.3 0.00040501999999999997 3.3 0.00040511999999999997 0 0.00040504 0 0.00040514 3.3 0.00040506 3.3 0.00040516 0 0.00040508 0 0.00040518 3.3 0.0004051 3.3 0.0004052 0 0.00040511999999999997 0 0.00040521999999999997 3.3 0.00040514 3.3 0.00040524 0 0.00040516 0 0.00040526 3.3 0.00040518 3.3 0.00040528 0 0.0004052 0 0.0004053 3.3 0.00040521999999999997 3.3 0.00040532 0 0.00040524 0 0.00040534 3.3 0.00040526 3.3 0.00040536 0 0.00040528 0 0.00040538 3.3 0.0004053 3.3 0.0004054 0 0.00040532 0 0.00040542 3.3 0.00040533999999999996 3.3 0.00040543999999999997 0 0.00040536 0 0.00040546 3.3 0.00040538 3.3 0.00040548 0 0.0004054 0 0.0004055 3.3 0.00040542 3.3 0.00040552 0 0.00040543999999999997 0 0.00040553999999999997 3.3 0.00040546 3.3 0.00040556 0 0.00040548 0 0.00040558 3.3 0.0004055 3.3 0.0004056 0 0.00040552 0 0.00040562 3.3 0.00040553999999999997 3.3 0.00040563999999999997 0 0.00040556 0 0.00040566 3.3 0.00040558 3.3 0.00040568 0 0.0004056 0 0.0004057 3.3 0.00040562 3.3 0.00040572 0 0.00040563999999999997 0 0.00040574 3.3 0.00040566 3.3 0.00040576 0 0.00040568 0 0.00040578 3.3 0.0004057 3.3 0.0004058 0 0.00040572 0 0.00040582 3.3 0.00040574 3.3 0.00040584 0 0.00040575999999999996 0 0.00040585999999999997 3.3 0.00040578 3.3 0.00040588 0 0.0004058 0 0.0004059 3.3 0.00040582 3.3 0.00040592 0 0.00040584 0 0.00040594 3.3 0.00040585999999999997 3.3 0.00040595999999999997 0 0.00040588 0 0.00040598 3.3 0.0004059 3.3 0.000406 0 0.00040592 0 0.00040602 3.3 0.00040594 3.3 0.00040604 0 0.00040595999999999997 0 0.00040605999999999997 3.3 0.00040598 3.3 0.00040608 0 0.000406 0 0.0004061 3.3 0.00040602 3.3 0.00040612 0 0.00040604 0 0.00040614 3.3 0.00040605999999999997 3.3 0.00040616 0 0.00040608 0 0.00040618 3.3 0.0004061 3.3 0.0004062 0 0.00040612 0 0.00040622 3.3 0.00040614 3.3 0.00040624 0 0.00040616 0 0.00040626 3.3 0.00040617999999999996 3.3 0.00040627999999999997 0 0.0004062 0 0.0004063 3.3 0.00040622 3.3 0.00040632 0 0.00040624 0 0.00040634 3.3 0.00040626 3.3 0.00040636 0 0.00040627999999999997 0 0.00040637999999999997 3.3 0.0004063 3.3 0.0004064 0 0.00040632 0 0.00040642 3.3 0.00040634 3.3 0.00040644 0 0.00040636 0 0.00040646 3.3 0.00040637999999999997 3.3 0.00040647999999999997 0 0.0004064 0 0.0004065 3.3 0.00040642 3.3 0.00040652 0 0.00040644 0 0.00040654 3.3 0.00040646 3.3 0.00040656 0 0.00040647999999999997 0 0.00040658 3.3 0.0004065 3.3 0.0004066 0 0.00040652 0 0.00040662 3.3 0.00040654 3.3 0.00040664 0 0.00040656 0 0.00040666 3.3 0.00040658 3.3 0.00040668 0 0.00040659999999999996 0 0.00040669999999999997 3.3 0.00040662 3.3 0.00040672 0 0.00040664 0 0.00040674 3.3 0.00040666 3.3 0.00040676 0 0.00040668 0 0.00040678 3.3 0.00040669999999999997 3.3 0.00040679999999999997 0 0.00040672 0 0.00040682 3.3 0.00040674 3.3 0.00040684 0 0.00040676 0 0.00040686 3.3 0.00040678 3.3 0.00040688 0 0.00040679999999999997 0 0.00040689999999999997 3.3 0.00040682 3.3 0.00040692 0 0.00040684 0 0.00040694 3.3 0.00040686 3.3 0.00040696 0 0.00040688 0 0.00040698 3.3 0.00040689999999999997 3.3 0.00040699999999999997 0 0.00040692 0 0.00040702 3.3 0.00040694 3.3 0.00040704 0 0.00040696 0 0.00040706 3.3 0.00040698 3.3 0.00040708 0 0.00040699999999999997 0 0.0004071 3.3 0.00040702 3.3 0.00040712 0 0.00040704 0 0.00040714 3.3 0.00040706 3.3 0.00040716 0 0.00040708 0 0.00040718 3.3 0.0004071 3.3 0.0004072 0 0.00040711999999999996 0 0.00040721999999999997 3.3 0.00040714 3.3 0.00040724 0 0.00040716 0 0.00040726 3.3 0.00040718 3.3 0.00040728 0 0.0004072 0 0.0004073 3.3 0.00040721999999999997 3.3 0.00040731999999999997 0 0.00040724 0 0.00040734 3.3 0.00040726 3.3 0.00040736 0 0.00040728 0 0.00040738 3.3 0.0004073 3.3 0.0004074 0 0.00040731999999999997 0 0.00040741999999999997 3.3 0.00040734 3.3 0.00040744 0 0.00040736 0 0.00040746 3.3 0.00040738 3.3 0.00040748 0 0.0004074 0 0.0004075 3.3 0.00040741999999999997 3.3 0.00040752 0 0.00040744 0 0.00040754 3.3 0.00040746 3.3 0.00040756 0 0.00040748 0 0.00040758 3.3 0.0004075 3.3 0.0004076 0 0.00040752 0 0.00040762 3.3 0.00040753999999999996 3.3 0.00040763999999999997 0 0.00040756 0 0.00040766 3.3 0.00040758 3.3 0.00040768 0 0.0004076 0 0.0004077 3.3 0.00040762 3.3 0.00040772 0 0.00040763999999999997 0 0.00040773999999999997 3.3 0.00040766 3.3 0.00040776 0 0.00040768 0 0.00040778 3.3 0.0004077 3.3 0.0004078 0 0.00040772 0 0.00040782 3.3 0.00040773999999999997 3.3 0.00040783999999999997 0 0.00040776 0 0.00040786 3.3 0.00040778 3.3 0.00040788 0 0.0004078 0 0.0004079 3.3 0.00040782 3.3 0.00040792 0 0.00040783999999999997 0 0.00040794 3.3 0.00040786 3.3 0.00040796 0 0.00040788 0 0.00040798 3.3 0.0004079 3.3 0.000408 0 0.00040792 0 0.00040802 3.3 0.00040794 3.3 0.00040804 0 0.00040795999999999996 0 0.00040805999999999997 3.3 0.00040798 3.3 0.00040808 0 0.000408 0 0.0004081 3.3 0.00040802 3.3 0.00040812 0 0.00040804 0 0.00040814 3.3 0.00040805999999999997 3.3 0.00040815999999999997 0 0.00040808 0 0.00040818 3.3 0.0004081 3.3 0.0004082 0 0.00040812 0 0.00040822 3.3 0.00040814 3.3 0.00040824 0 0.00040815999999999997 0 0.00040825999999999997 3.3 0.00040818 3.3 0.00040828 0 0.0004082 0 0.0004083 3.3 0.00040822 3.3 0.00040832 0 0.00040824 0 0.00040834 3.3 0.00040825999999999997 3.3 0.00040836 0 0.00040828 0 0.00040838 3.3 0.0004083 3.3 0.0004084 0 0.00040832 0 0.00040842 3.3 0.00040834 3.3 0.00040844 0 0.00040836 0 0.00040846 3.3 0.00040837999999999996 3.3 0.00040847999999999997 0 0.0004084 0 0.0004085 3.3 0.00040842 3.3 0.00040852 0 0.00040844 0 0.00040854 3.3 0.00040846 3.3 0.00040856 0 0.00040847999999999997 0 0.00040857999999999997 3.3 0.0004085 3.3 0.0004086 0 0.00040852 0 0.00040862 3.3 0.00040854 3.3 0.00040864 0 0.00040856 0 0.00040866 3.3 0.00040857999999999997 3.3 0.00040867999999999997 0 0.0004086 0 0.0004087 3.3 0.00040862 3.3 0.00040872 0 0.00040864 0 0.00040874 3.3 0.00040866 3.3 0.00040876 0 0.00040867999999999997 0 0.00040877999999999997 3.3 0.0004087 3.3 0.0004088 0 0.00040872 0 0.00040882 3.3 0.00040874 3.3 0.00040884 0 0.00040876 0 0.00040886 3.3 0.00040877999999999997 3.3 0.00040888 0 0.0004088 0 0.0004089 3.3 0.00040882 3.3 0.00040892 0 0.00040884 0 0.00040894 3.3 0.00040886 3.3 0.00040896 0 0.00040888 0 0.00040898 3.3 0.00040889999999999996 3.3 0.00040899999999999997 0 0.00040892 0 0.00040902 3.3 0.00040894 3.3 0.00040904 0 0.00040896 0 0.00040906 3.3 0.00040898 3.3 0.00040908 0 0.00040899999999999997 0 0.00040909999999999997 3.3 0.00040902 3.3 0.00040912 0 0.00040904 0 0.00040914 3.3 0.00040906 3.3 0.00040916 0 0.00040908 0 0.00040918 3.3 0.00040909999999999997 3.3 0.00040919999999999997 0 0.00040912 0 0.00040922 3.3 0.00040914 3.3 0.00040924 0 0.00040916 0 0.00040926 3.3 0.00040918 3.3 0.00040928 0 0.00040919999999999997 0 0.0004093 3.3 0.00040922 3.3 0.00040932 0 0.00040924 0 0.00040934 3.3 0.00040926 3.3 0.00040936 0 0.00040928 0 0.00040938 3.3 0.0004093 3.3 0.0004094 0 0.00040931999999999996 0 0.00040941999999999997 3.3 0.00040934 3.3 0.00040944 0 0.00040936 0 0.00040946 3.3 0.00040938 3.3 0.00040948 0 0.0004094 0 0.0004095 3.3 0.00040941999999999997 3.3 0.00040951999999999997 0 0.00040944 0 0.00040954 3.3 0.00040946 3.3 0.00040956 0 0.00040948 0 0.00040958 3.3 0.0004095 3.3 0.0004096 0 0.00040951999999999997 0 0.00040961999999999997 3.3 0.00040954 3.3 0.00040964 0 0.00040956 0 0.00040966 3.3 0.00040958 3.3 0.00040968 0 0.0004096 0 0.0004097 3.3 0.00040961999999999997 3.3 0.00040972 0 0.00040964 0 0.00040974 3.3 0.00040966 3.3 0.00040976 0 0.00040968 0 0.00040978 3.3 0.0004097 3.3 0.0004098 0 0.00040972 0 0.00040982 3.3 0.00040973999999999996 3.3 0.00040983999999999997 0 0.00040976 0 0.00040986 3.3 0.00040978 3.3 0.00040988 0 0.0004098 0 0.0004099 3.3 0.00040982 3.3 0.00040992 0 0.00040983999999999997 0 0.00040993999999999997 3.3 0.00040986 3.3 0.00040996 0 0.00040988 0 0.00040998 3.3 0.0004099 3.3 0.00041 0 0.00040992 0 0.00041002 3.3 0.00040993999999999997 3.3 0.00041003999999999997 0 0.00040996 0 0.00041006 3.3 0.00040998 3.3 0.00041008 0 0.00041 0 0.0004101 3.3 0.00041002 3.3 0.00041012 0 0.00041003999999999997 0 0.00041014 3.3 0.00041006 3.3 0.00041016 0 0.00041008 0 0.00041018 3.3 0.0004101 3.3 0.0004102 0 0.00041012 0 0.00041022 3.3 0.00041014 3.3 0.00041024 0 0.00041015999999999996 0 0.00041025999999999996 3.3 0.00041018 3.3 0.00041028 0 0.0004102 0 0.0004103 3.3 0.00041022 3.3 0.00041032 0 0.00041024 0 0.00041034 3.3 0.00041025999999999996 3.3 0.00041035999999999997 0 0.00041028 0 0.00041038 3.3 0.0004103 3.3 0.0004104 0 0.00041032 0 0.00041042 3.3 0.00041034 3.3 0.00041044 0 0.00041035999999999997 0 0.00041045999999999997 3.3 0.00041038 3.3 0.00041048 0 0.0004104 0 0.0004105 3.3 0.00041042 3.3 0.00041052 0 0.00041044 0 0.00041054 3.3 0.00041045999999999997 3.3 0.00041055999999999997 0 0.00041048 0 0.00041058 3.3 0.0004105 3.3 0.0004106 0 0.00041052 0 0.00041062 3.3 0.00041054 3.3 0.00041064 0 0.00041055999999999997 0 0.00041066 3.3 0.00041058 3.3 0.00041068 0 0.0004106 0 0.0004107 3.3 0.00041062 3.3 0.00041072 0 0.00041064 0 0.00041074 3.3 0.00041066 3.3 0.00041076 0 0.00041067999999999996 0 0.00041077999999999997 3.3 0.0004107 3.3 0.0004108 0 0.00041072 0 0.00041082 3.3 0.00041074 3.3 0.00041084 0 0.00041076 0 0.00041086 3.3 0.00041077999999999997 3.3 0.00041087999999999997 0 0.0004108 0 0.0004109 3.3 0.00041082 3.3 0.00041092 0 0.00041084 0 0.00041094 3.3 0.00041086 3.3 0.00041096 0 0.00041087999999999997 0 0.00041097999999999997 3.3 0.0004109 3.3 0.000411 0 0.00041092 0 0.00041102 3.3 0.00041094 3.3 0.00041104 0 0.00041096 0 0.00041106 3.3 0.00041097999999999997 3.3 0.00041108 0 0.000411 0 0.0004111 3.3 0.00041102 3.3 0.00041112 0 0.00041104 0 0.00041114 3.3 0.00041106 3.3 0.00041116 0 0.00041108 0 0.00041118 3.3 0.00041109999999999996 3.3 0.00041119999999999997 0 0.00041112 0 0.00041122 3.3 0.00041114 3.3 0.00041124 0 0.00041116 0 0.00041126 3.3 0.00041118 3.3 0.00041128 0 0.00041119999999999997 0 0.00041129999999999997 3.3 0.00041122 3.3 0.00041132 0 0.00041124 0 0.00041134 3.3 0.00041126 3.3 0.00041136 0 0.00041128 0 0.00041138 3.3 0.00041129999999999997 3.3 0.00041139999999999997 0 0.00041132 0 0.00041142 3.3 0.00041134 3.3 0.00041144 0 0.00041136 0 0.00041146 3.3 0.00041138 3.3 0.00041148 0 0.00041139999999999997 0 0.0004115 3.3 0.00041142 3.3 0.00041152 0 0.00041144 0 0.00041154 3.3 0.00041146 3.3 0.00041156 0 0.00041148 0 0.00041158 3.3 0.0004115 3.3 0.0004116 0 0.00041151999999999996 0 0.00041161999999999997 3.3 0.00041154 3.3 0.00041164 0 0.00041156 0 0.00041166 3.3 0.00041158 3.3 0.00041168 0 0.0004116 0 0.0004117 3.3 0.00041161999999999997 3.3 0.00041171999999999997 0 0.00041164 0 0.00041174 3.3 0.00041166 3.3 0.00041176 0 0.00041168 0 0.00041178 3.3 0.0004117 3.3 0.0004118 0 0.00041171999999999997 0 0.00041181999999999997 3.3 0.00041174 3.3 0.00041184 0 0.00041176 0 0.00041186 3.3 0.00041178 3.3 0.00041188 0 0.0004118 0 0.0004119 3.3 0.00041181999999999997 3.3 0.00041191999999999997 0 0.00041184 0 0.00041194 3.3 0.00041186 3.3 0.00041196 0 0.00041188 0 0.00041198 3.3 0.0004119 3.3 0.000412 0 0.00041191999999999997 0 0.00041202 3.3 0.00041193999999999996 3.3 0.00041203999999999996 0 0.00041196 0 0.00041206 3.3 0.00041198 3.3 0.00041208 0 0.000412 0 0.0004121 3.3 0.00041202 3.3 0.00041212 0 0.00041203999999999996 0 0.00041213999999999997 3.3 0.00041206 3.3 0.00041216 0 0.00041208 0 0.00041218 3.3 0.0004121 3.3 0.0004122 0 0.00041212 0 0.00041222 3.3 0.00041213999999999997 3.3 0.00041223999999999997 0 0.00041216 0 0.00041226 3.3 0.00041218 3.3 0.00041228 0 0.0004122 0 0.0004123 3.3 0.00041222 3.3 0.00041232 0 0.00041223999999999997 0 0.00041233999999999997 3.3 0.00041226 3.3 0.00041236 0 0.00041228 0 0.00041238 3.3 0.0004123 3.3 0.0004124 0 0.00041232 0 0.00041242 3.3 0.00041233999999999997 3.3 0.00041244 0 0.00041236 0 0.00041246 3.3 0.00041238 3.3 0.00041248 0 0.0004124 0 0.0004125 3.3 0.00041242 3.3 0.00041252 0 0.00041244 0 0.00041254 3.3 0.00041245999999999996 3.3 0.00041255999999999997 0 0.00041248 0 0.00041258 3.3 0.0004125 3.3 0.0004126 0 0.00041252 0 0.00041262 3.3 0.00041254 3.3 0.00041264 0 0.00041255999999999997 0 0.00041265999999999997 3.3 0.00041258 3.3 0.00041268 0 0.0004126 0 0.0004127 3.3 0.00041262 3.3 0.00041272 0 0.00041264 0 0.00041274 3.3 0.00041265999999999997 3.3 0.00041275999999999997 0 0.00041268 0 0.00041278 3.3 0.0004127 3.3 0.0004128 0 0.00041272 0 0.00041282 3.3 0.00041274 3.3 0.00041284 0 0.00041275999999999997 0 0.00041286 3.3 0.00041278 3.3 0.00041288 0 0.0004128 0 0.0004129 3.3 0.00041282 3.3 0.00041292 0 0.00041284 0 0.00041294 3.3 0.00041286 3.3 0.00041296 0 0.00041287999999999996 0 0.00041297999999999997 3.3 0.0004129 3.3 0.000413 0 0.00041292 0 0.00041302 3.3 0.00041294 3.3 0.00041304 0 0.00041296 0 0.00041306 3.3 0.00041297999999999997 3.3 0.00041307999999999997 0 0.000413 0 0.0004131 3.3 0.00041302 3.3 0.00041312 0 0.00041304 0 0.00041314 3.3 0.00041306 3.3 0.00041316 0 0.00041307999999999997 0 0.00041317999999999997 3.3 0.0004131 3.3 0.0004132 0 0.00041312 0 0.00041322 3.3 0.00041314 3.3 0.00041324 0 0.00041316 0 0.00041326 3.3 0.00041317999999999997 3.3 0.00041328 0 0.0004132 0 0.0004133 3.3 0.00041322 3.3 0.00041332 0 0.00041324 0 0.00041334 3.3 0.00041326 3.3 0.00041336 0 0.00041328 0 0.00041338 3.3 0.00041329999999999996 3.3 0.00041339999999999997 0 0.00041332 0 0.00041342 3.3 0.00041334 3.3 0.00041344 0 0.00041336 0 0.00041346 3.3 0.00041338 3.3 0.00041348 0 0.00041339999999999997 0 0.00041349999999999997 3.3 0.00041342 3.3 0.00041352 0 0.00041344 0 0.00041354 3.3 0.00041346 3.3 0.00041356 0 0.00041348 0 0.00041358 3.3 0.00041349999999999997 3.3 0.00041359999999999997 0 0.00041352 0 0.00041362 3.3 0.00041354 3.3 0.00041364 0 0.00041356 0 0.00041366 3.3 0.00041358 3.3 0.00041368 0 0.00041359999999999997 0 0.00041369999999999997 3.3 0.00041362 3.3 0.00041372 0 0.00041364 0 0.00041374 3.3 0.00041366 3.3 0.00041376 0 0.00041368 0 0.00041378 3.3 0.00041369999999999997 3.3 0.0004138 0 0.00041371999999999996 0 0.00041381999999999996 3.3 0.00041374 3.3 0.00041384 0 0.00041376 0 0.00041386 3.3 0.00041378 3.3 0.00041388 0 0.0004138 0 0.0004139 3.3 0.00041381999999999996 3.3 0.00041391999999999997 0 0.00041384 0 0.00041394 3.3 0.00041386 3.3 0.00041396 0 0.00041388 0 0.00041398 3.3 0.0004139 3.3 0.000414 0 0.00041391999999999997 0 0.00041401999999999997 3.3 0.00041394 3.3 0.00041404 0 0.00041396 0 0.00041406 3.3 0.00041398 3.3 0.00041408 0 0.000414 0 0.0004141 3.3 0.00041401999999999997 3.3 0.00041411999999999997 0 0.00041404 0 0.00041414 3.3 0.00041406 3.3 0.00041416 0 0.00041408 0 0.00041418 3.3 0.0004141 3.3 0.0004142 0 0.00041411999999999997 0 0.00041422 3.3 0.00041414 3.3 0.00041424 0 0.00041416 0 0.00041426 3.3 0.00041418 3.3 0.00041428 0 0.0004142 0 0.0004143 3.3 0.00041422 3.3 0.00041432 0 0.00041423999999999996 0 0.00041433999999999997 3.3 0.00041426 3.3 0.00041436 0 0.00041428 0 0.00041438 3.3 0.0004143 3.3 0.0004144 0 0.00041432 0 0.00041442 3.3 0.00041433999999999997 3.3 0.00041443999999999997 0 0.00041436 0 0.00041446 3.3 0.00041438 3.3 0.00041448 0 0.0004144 0 0.0004145 3.3 0.00041442 3.3 0.00041452 0 0.00041443999999999997 0 0.00041453999999999997 3.3 0.00041446 3.3 0.00041456 0 0.00041448 0 0.00041458 3.3 0.0004145 3.3 0.0004146 0 0.00041452 0 0.00041462 3.3 0.00041453999999999997 3.3 0.00041464 0 0.00041456 0 0.00041466 3.3 0.00041458 3.3 0.00041468 0 0.0004146 0 0.0004147 3.3 0.00041462 3.3 0.00041472 0 0.00041464 0 0.00041474 3.3 0.00041465999999999996 3.3 0.00041475999999999997 0 0.00041468 0 0.00041478 3.3 0.0004147 3.3 0.0004148 0 0.00041472 0 0.00041482 3.3 0.00041474 3.3 0.00041484 0 0.00041475999999999997 0 0.00041485999999999997 3.3 0.00041478 3.3 0.00041488 0 0.0004148 0 0.0004149 3.3 0.00041482 3.3 0.00041492 0 0.00041484 0 0.00041494 3.3 0.00041485999999999997 3.3 0.00041495999999999997 0 0.00041488 0 0.00041498 3.3 0.0004149 3.3 0.000415 0 0.00041492 0 0.00041502 3.3 0.00041494 3.3 0.00041504 0 0.00041495999999999997 0 0.00041506 3.3 0.00041498 3.3 0.00041508 0 0.000415 0 0.0004151 3.3 0.00041502 3.3 0.00041512 0 0.00041504 0 0.00041514 3.3 0.00041506 3.3 0.00041516 0 0.00041507999999999996 0 0.00041517999999999997 3.3 0.0004151 3.3 0.0004152 0 0.00041512 0 0.00041522 3.3 0.00041514 3.3 0.00041524 0 0.00041516 0 0.00041526 3.3 0.00041517999999999997 3.3 0.00041527999999999997 0 0.0004152 0 0.0004153 3.3 0.00041522 3.3 0.00041532 0 0.00041524 0 0.00041534 3.3 0.00041526 3.3 0.00041536 0 0.00041527999999999997 0 0.00041537999999999997 3.3 0.0004153 3.3 0.0004154 0 0.00041532 0 0.00041542 3.3 0.00041534 3.3 0.00041544 0 0.00041536 0 0.00041546 3.3 0.00041537999999999997 3.3 0.00041547999999999997 0 0.0004154 0 0.0004155 3.3 0.00041542 3.3 0.00041552 0 0.00041544 0 0.00041554 3.3 0.00041546 3.3 0.00041556 0 0.00041547999999999997 0 0.00041558 3.3 0.00041549999999999996 3.3 0.00041559999999999996 0 0.00041552 0 0.00041562 3.3 0.00041554 3.3 0.00041564 0 0.00041556 0 0.00041566 3.3 0.00041558 3.3 0.00041568 0 0.00041559999999999996 0 0.00041569999999999997 3.3 0.00041562 3.3 0.00041572 0 0.00041564 0 0.00041574 3.3 0.00041566 3.3 0.00041576 0 0.00041568 0 0.00041578 3.3 0.00041569999999999997 3.3 0.00041579999999999997 0 0.00041572 0 0.00041582 3.3 0.00041574 3.3 0.00041584 0 0.00041576 0 0.00041586 3.3 0.00041578 3.3 0.00041588 0 0.00041579999999999997 0 0.00041589999999999997 3.3 0.00041582 3.3 0.00041592 0 0.00041584 0 0.00041594 3.3 0.00041586 3.3 0.00041596 0 0.00041588 0 0.00041598 3.3 0.00041589999999999997 3.3 0.000416 0 0.00041592 0 0.00041602 3.3 0.00041594 3.3 0.00041604 0 0.00041596 0 0.00041606 3.3 0.00041598 3.3 0.00041608 0 0.000416 0 0.0004161 3.3 0.00041601999999999996 3.3 0.00041611999999999997 0 0.00041604 0 0.00041614 3.3 0.00041606 3.3 0.00041616 0 0.00041608 0 0.00041618 3.3 0.0004161 3.3 0.0004162 0 0.00041611999999999997 0 0.00041621999999999997 3.3 0.00041614 3.3 0.00041624 0 0.00041616 0 0.00041626 3.3 0.00041618 3.3 0.00041628 0 0.0004162 0 0.0004163 3.3 0.00041621999999999997 3.3 0.00041631999999999997 0 0.00041624 0 0.00041634 3.3 0.00041626 3.3 0.00041636 0 0.00041628 0 0.00041638 3.3 0.0004163 3.3 0.0004164 0 0.00041631999999999997 0 0.00041642 3.3 0.00041634 3.3 0.00041644 0 0.00041636 0 0.00041646 3.3 0.00041638 3.3 0.00041648 0 0.0004164 0 0.0004165 3.3 0.00041642 3.3 0.00041652 0 0.00041643999999999996 0 0.00041653999999999997 3.3 0.00041646 3.3 0.00041656 0 0.00041648 0 0.00041658 3.3 0.0004165 3.3 0.0004166 0 0.00041652 0 0.00041662 3.3 0.00041653999999999997 3.3 0.00041663999999999997 0 0.00041656 0 0.00041666 3.3 0.00041658 3.3 0.00041668 0 0.0004166 0 0.0004167 3.3 0.00041662 3.3 0.00041672 0 0.00041663999999999997 0 0.00041673999999999997 3.3 0.00041666 3.3 0.00041676 0 0.00041668 0 0.00041678 3.3 0.0004167 3.3 0.0004168 0 0.00041672 0 0.00041682 3.3 0.00041673999999999997 3.3 0.00041684 0 0.00041676 0 0.00041686 3.3 0.00041678 3.3 0.00041688 0 0.0004168 0 0.0004169 3.3 0.00041682 3.3 0.00041692 0 0.00041684 0 0.00041694 3.3 0.00041685999999999996 3.3 0.00041695999999999997 0 0.00041688 0 0.00041698 3.3 0.0004169 3.3 0.000417 0 0.00041692 0 0.00041702 3.3 0.00041694 3.3 0.00041704 0 0.00041695999999999997 0 0.00041705999999999997 3.3 0.00041698 3.3 0.00041708 0 0.000417 0 0.0004171 3.3 0.00041702 3.3 0.00041712 0 0.00041704 0 0.00041714 3.3 0.00041705999999999997 3.3 0.00041715999999999997 0 0.00041708 0 0.00041718 3.3 0.0004171 3.3 0.0004172 0 0.00041712 0 0.00041722 3.3 0.00041714 3.3 0.00041724 0 0.00041715999999999997 0 0.00041725999999999997 3.3 0.00041718 3.3 0.00041728 0 0.0004172 0 0.0004173 3.3 0.00041722 3.3 0.00041732 0 0.00041724 0 0.00041734 3.3 0.00041725999999999997 3.3 0.00041736 0 0.00041727999999999996 0 0.00041737999999999996 3.3 0.0004173 3.3 0.0004174 0 0.00041732 0 0.00041742 3.3 0.00041734 3.3 0.00041744 0 0.00041736 0 0.00041746 3.3 0.00041737999999999996 3.3 0.00041747999999999997 0 0.0004174 0 0.0004175 3.3 0.00041742 3.3 0.00041752 0 0.00041744 0 0.00041754 3.3 0.00041746 3.3 0.00041756 0 0.00041747999999999997 0 0.00041757999999999997 3.3 0.0004175 3.3 0.0004176 0 0.00041752 0 0.00041762 3.3 0.00041754 3.3 0.00041764 0 0.00041756 0 0.00041766 3.3 0.00041757999999999997 3.3 0.00041767999999999997 0 0.0004176 0 0.0004177 3.3 0.00041762 3.3 0.00041772 0 0.00041764 0 0.00041774 3.3 0.00041766 3.3 0.00041776 0 0.00041767999999999997 0 0.00041778 3.3 0.0004177 3.3 0.0004178 0 0.00041772 0 0.00041782 3.3 0.00041774 3.3 0.00041784 0 0.00041776 0 0.00041786 3.3 0.00041778 3.3 0.00041788 0 0.00041779999999999996 0 0.00041789999999999997 3.3 0.00041782 3.3 0.00041792 0 0.00041784 0 0.00041794 3.3 0.00041786 3.3 0.00041796 0 0.00041788 0 0.00041798 3.3 0.00041789999999999997 3.3 0.00041799999999999997 0 0.00041792 0 0.00041802 3.3 0.00041794 3.3 0.00041804 0 0.00041796 0 0.00041806 3.3 0.00041798 3.3 0.00041808 0 0.00041799999999999997 0 0.00041809999999999997 3.3 0.00041802 3.3 0.00041812 0 0.00041804 0 0.00041814 3.3 0.00041806 3.3 0.00041816 0 0.00041808 0 0.00041818 3.3 0.00041809999999999997 3.3 0.0004182 0 0.00041812 0 0.00041822 3.3 0.00041814 3.3 0.00041824 0 0.00041816 0 0.00041826 3.3 0.00041818 3.3 0.00041828 0 0.0004182 0 0.0004183 3.3 0.00041821999999999996 3.3 0.00041831999999999997 0 0.00041824 0 0.00041834 3.3 0.00041826 3.3 0.00041836 0 0.00041828 0 0.00041838 3.3 0.0004183 3.3 0.0004184 0 0.00041831999999999997 0 0.00041841999999999997 3.3 0.00041834 3.3 0.00041844 0 0.00041836 0 0.00041846 3.3 0.00041838 3.3 0.00041848 0 0.0004184 0 0.0004185 3.3 0.00041841999999999997 3.3 0.00041851999999999997 0 0.00041844 0 0.00041854 3.3 0.00041846 3.3 0.00041856 0 0.00041848 0 0.00041858 3.3 0.0004185 3.3 0.0004186 0 0.00041851999999999997 0 0.00041862 3.3 0.00041854 3.3 0.00041864 0 0.00041856 0 0.00041866 3.3 0.00041858 3.3 0.00041868 0 0.0004186 0 0.0004187 3.3 0.00041862 3.3 0.00041872 0 0.00041863999999999996 0 0.00041873999999999997 3.3 0.00041866 3.3 0.00041876 0 0.00041868 0 0.00041878 3.3 0.0004187 3.3 0.0004188 0 0.00041872 0 0.00041882 3.3 0.00041873999999999997 3.3 0.00041883999999999997 0 0.00041876 0 0.00041886 3.3 0.00041878 3.3 0.00041888 0 0.0004188 0 0.0004189 3.3 0.00041882 3.3 0.00041892 0 0.00041883999999999997 0 0.00041893999999999997 3.3 0.00041886 3.3 0.00041896 0 0.00041888 0 0.00041898 3.3 0.0004189 3.3 0.000419 0 0.00041892 0 0.00041902 3.3 0.00041893999999999997 3.3 0.00041903999999999997 0 0.00041896 0 0.00041906 3.3 0.00041898 3.3 0.00041908 0 0.000419 0 0.0004191 3.3 0.00041902 3.3 0.00041912 0 0.00041903999999999997 0 0.00041914 3.3 0.00041905999999999996 3.3 0.00041915999999999996 0 0.00041908 0 0.00041918 3.3 0.0004191 3.3 0.0004192 0 0.00041912 0 0.00041922 3.3 0.00041914 3.3 0.00041924 0 0.00041915999999999996 0 0.00041925999999999997 3.3 0.00041918 3.3 0.00041928 0 0.0004192 0 0.0004193 3.3 0.00041922 3.3 0.00041932 0 0.00041924 0 0.00041934 3.3 0.00041925999999999997 3.3 0.00041935999999999997 0 0.00041928 0 0.00041938 3.3 0.0004193 3.3 0.0004194 0 0.00041932 0 0.00041942 3.3 0.00041934 3.3 0.00041944 0 0.00041935999999999997 0 0.00041945999999999997 3.3 0.00041938 3.3 0.00041948 0 0.0004194 0 0.0004195 3.3 0.00041942 3.3 0.00041952 0 0.00041944 0 0.00041954 3.3 0.00041945999999999997 3.3 0.00041956 0 0.00041948 0 0.00041958 3.3 0.0004195 3.3 0.0004196 0 0.00041952 0 0.00041962 3.3 0.00041954 3.3 0.00041964 0 0.00041956 0 0.00041966 3.3 0.00041957999999999996 3.3 0.00041967999999999997 0 0.0004196 0 0.0004197 3.3 0.00041962 3.3 0.00041972 0 0.00041964 0 0.00041974 3.3 0.00041966 3.3 0.00041976 0 0.00041967999999999997 0 0.00041977999999999997 3.3 0.0004197 3.3 0.0004198 0 0.00041972 0 0.00041982 3.3 0.00041974 3.3 0.00041984 0 0.00041976 0 0.00041986 3.3 0.00041977999999999997 3.3 0.00041987999999999997 0 0.0004198 0 0.0004199 3.3 0.00041982 3.3 0.00041992 0 0.00041984 0 0.00041994 3.3 0.00041986 3.3 0.00041996 0 0.00041987999999999997 0 0.00041998 3.3 0.0004199 3.3 0.00042 0 0.00041992 0 0.00042002 3.3 0.00041994 3.3 0.00042004 0 0.00041996 0 0.00042006 3.3 0.00041998 3.3 0.00042008 0 0.00041999999999999996 0 0.00042009999999999997 3.3 0.00042002 3.3 0.00042012 0 0.00042004 0 0.00042014 3.3 0.00042006 3.3 0.00042016 0 0.00042008 0 0.00042018 3.3 0.00042009999999999997 3.3 0.00042019999999999997 0 0.00042012 0 0.00042022 3.3 0.00042014 3.3 0.00042024 0 0.00042016 0 0.00042026 3.3 0.00042018 3.3 0.00042028 0 0.00042019999999999997 0 0.00042029999999999997 3.3 0.00042022 3.3 0.00042032 0 0.00042024 0 0.00042034 3.3 0.00042026 3.3 0.00042036 0 0.00042028 0 0.00042038 3.3 0.00042029999999999997 3.3 0.0004204 0 0.00042032 0 0.00042042 3.3 0.00042034 3.3 0.00042044 0 0.00042036 0 0.00042046 3.3 0.00042038 3.3 0.00042048 0 0.0004204 0 0.0004205 3.3 0.00042041999999999996 3.3 0.00042051999999999997 0 0.00042044 0 0.00042054 3.3 0.00042046 3.3 0.00042056 0 0.00042048 0 0.00042058 3.3 0.0004205 3.3 0.0004206 0 0.00042051999999999997 0 0.00042061999999999997 3.3 0.00042054 3.3 0.00042064 0 0.00042056 0 0.00042066 3.3 0.00042058 3.3 0.00042068 0 0.0004206 0 0.0004207 3.3 0.00042061999999999997 3.3 0.00042071999999999997 0 0.00042064 0 0.00042074 3.3 0.00042066 3.3 0.00042076 0 0.00042068 0 0.00042078 3.3 0.0004207 3.3 0.0004208 0 0.00042071999999999997 0 0.00042081999999999997 3.3 0.00042074 3.3 0.00042084 0 0.00042076 0 0.00042086 3.3 0.00042078 3.3 0.00042088 0 0.0004208 0 0.0004209 3.3 0.00042081999999999997 3.3 0.00042092 0 0.00042084 0 0.00042094 3.3 0.00042086 3.3 0.00042096 0 0.00042088 0 0.00042098 3.3 0.0004209 3.3 0.000421 0 0.00042092 0 0.00042102 3.3 0.00042093999999999996 3.3 0.00042103999999999997 0 0.00042096 0 0.00042106 3.3 0.00042098 3.3 0.00042108 0 0.000421 0 0.0004211 3.3 0.00042102 3.3 0.00042112 0 0.00042103999999999997 0 0.00042113999999999997 3.3 0.00042106 3.3 0.00042116 0 0.00042108 0 0.00042118 3.3 0.0004211 3.3 0.0004212 0 0.00042112 0 0.00042122 3.3 0.00042113999999999997 3.3 0.00042123999999999997 0 0.00042116 0 0.00042126 3.3 0.00042118 3.3 0.00042128 0 0.0004212 0 0.0004213 3.3 0.00042122 3.3 0.00042132 0 0.00042123999999999997 0 0.00042134 3.3 0.00042126 3.3 0.00042136 0 0.00042128 0 0.00042138 3.3 0.0004213 3.3 0.0004214 0 0.00042132 0 0.00042142 3.3 0.00042134 3.3 0.00042144 0 0.00042135999999999996 0 0.00042145999999999997 3.3 0.00042138 3.3 0.00042148 0 0.0004214 0 0.0004215 3.3 0.00042142 3.3 0.00042152 0 0.00042144 0 0.00042154 3.3 0.00042145999999999997 3.3 0.00042155999999999997 0 0.00042148 0 0.00042158 3.3 0.0004215 3.3 0.0004216 0 0.00042152 0 0.00042162 3.3 0.00042154 3.3 0.00042164 0 0.00042155999999999997 0 0.00042165999999999997 3.3 0.00042158 3.3 0.00042168 0 0.0004216 0 0.0004217 3.3 0.00042162 3.3 0.00042172 0 0.00042164 0 0.00042174 3.3 0.00042165999999999997 3.3 0.00042176 0 0.00042168 0 0.00042178 3.3 0.0004217 3.3 0.0004218 0 0.00042172 0 0.00042182 3.3 0.00042174 3.3 0.00042184 0 0.00042176 0 0.00042186 3.3 0.00042177999999999996 3.3 0.00042187999999999997 0 0.0004218 0 0.0004219 3.3 0.00042182 3.3 0.00042192 0 0.00042184 0 0.00042194 3.3 0.00042186 3.3 0.00042196 0 0.00042187999999999997 0 0.00042197999999999997 3.3 0.0004219 3.3 0.000422 0 0.00042192 0 0.00042202 3.3 0.00042194 3.3 0.00042204 0 0.00042196 0 0.00042206 3.3 0.00042197999999999997 3.3 0.00042207999999999997 0 0.000422 0 0.0004221 3.3 0.00042202 3.3 0.00042212 0 0.00042204 0 0.00042214 3.3 0.00042206 3.3 0.00042216 0 0.00042207999999999997 0 0.00042217999999999997 3.3 0.0004221 3.3 0.0004222 0 0.00042212 0 0.00042222 3.3 0.00042214 3.3 0.00042224 0 0.00042216 0 0.00042226 3.3 0.00042217999999999997 3.3 0.00042228 0 0.00042219999999999996 0 0.00042229999999999996 3.3 0.00042222 3.3 0.00042232 0 0.00042224 0 0.00042234 3.3 0.00042226 3.3 0.00042236 0 0.00042228 0 0.00042238 3.3 0.00042229999999999996 3.3 0.00042239999999999997 0 0.00042232 0 0.00042242 3.3 0.00042234 3.3 0.00042244 0 0.00042236 0 0.00042246 3.3 0.00042238 3.3 0.00042248 0 0.00042239999999999997 0 0.00042249999999999997 3.3 0.00042242 3.3 0.00042252 0 0.00042244 0 0.00042254 3.3 0.00042246 3.3 0.00042256 0 0.00042248 0 0.00042258 3.3 0.00042249999999999997 3.3 0.00042259999999999997 0 0.00042252 0 0.00042262 3.3 0.00042254 3.3 0.00042264 0 0.00042256 0 0.00042266 3.3 0.00042258 3.3 0.00042268 0 0.00042259999999999997 0 0.0004227 3.3 0.00042262 3.3 0.00042272 0 0.00042264 0 0.00042274 3.3 0.00042266 3.3 0.00042276 0 0.00042268 0 0.00042278 3.3 0.0004227 3.3 0.0004228 0 0.00042271999999999996 0 0.00042281999999999997 3.3 0.00042274 3.3 0.00042284 0 0.00042276 0 0.00042286 3.3 0.00042278 3.3 0.00042288 0 0.0004228 0 0.0004229 3.3 0.00042281999999999997 3.3 0.00042291999999999997 0 0.00042284 0 0.00042294 3.3 0.00042286 3.3 0.00042296 0 0.00042288 0 0.00042298 3.3 0.0004229 3.3 0.000423 0 0.00042291999999999997 0 0.00042301999999999997 3.3 0.00042294 3.3 0.00042304 0 0.00042296 0 0.00042306 3.3 0.00042298 3.3 0.00042308 0 0.000423 0 0.0004231 3.3 0.00042301999999999997 3.3 0.00042312 0 0.00042304 0 0.00042314 3.3 0.00042306 3.3 0.00042316 0 0.00042308 0 0.00042318 3.3 0.0004231 3.3 0.0004232 0 0.00042312 0 0.00042322 3.3 0.00042313999999999996 3.3 0.00042323999999999997 0 0.00042316 0 0.00042326 3.3 0.00042318 3.3 0.00042328 0 0.0004232 0 0.0004233 3.3 0.00042322 3.3 0.00042332 0 0.00042323999999999997 0 0.00042333999999999997 3.3 0.00042326 3.3 0.00042336 0 0.00042328 0 0.00042338 3.3 0.0004233 3.3 0.0004234 0 0.00042332 0 0.00042342 3.3 0.00042333999999999997 3.3 0.00042343999999999997 0 0.00042336 0 0.00042346 3.3 0.00042338 3.3 0.00042348 0 0.0004234 0 0.0004235 3.3 0.00042342 3.3 0.00042352 0 0.00042343999999999997 0 0.00042354 3.3 0.00042346 3.3 0.00042356 0 0.00042348 0 0.00042358 3.3 0.0004235 3.3 0.0004236 0 0.00042352 0 0.00042362 3.3 0.00042354 3.3 0.00042364 0 0.00042355999999999996 0 0.00042365999999999997 3.3 0.00042358 3.3 0.00042368 0 0.0004236 0 0.0004237 3.3 0.00042362 3.3 0.00042372 0 0.00042364 0 0.00042374 3.3 0.00042365999999999997 3.3 0.00042375999999999997 0 0.00042368 0 0.00042378 3.3 0.0004237 3.3 0.0004238 0 0.00042372 0 0.00042382 3.3 0.00042374 3.3 0.00042384 0 0.00042375999999999997 0 0.00042385999999999997 3.3 0.00042378 3.3 0.00042388 0 0.0004238 0 0.0004239 3.3 0.00042382 3.3 0.00042392 0 0.00042384 0 0.00042394 3.3 0.00042385999999999997 3.3 0.00042395999999999997 0 0.00042388 0 0.00042398 3.3 0.0004239 3.3 0.000424 0 0.00042392 0 0.00042402 3.3 0.00042394 3.3 0.00042404 0 0.00042395999999999997 0 0.00042406 3.3 0.00042397999999999996 3.3 0.00042407999999999996 0 0.000424 0 0.0004241 3.3 0.00042402 3.3 0.00042412 0 0.00042404 0 0.00042414 3.3 0.00042406 3.3 0.00042416 0 0.00042407999999999996 0 0.00042417999999999997 3.3 0.0004241 3.3 0.0004242 0 0.00042412 0 0.00042422 3.3 0.00042414 3.3 0.00042424 0 0.00042416 0 0.00042426 3.3 0.00042417999999999997 3.3 0.00042427999999999997 0 0.0004242 0 0.0004243 3.3 0.00042422 3.3 0.00042432 0 0.00042424 0 0.00042434 3.3 0.00042426 3.3 0.00042436 0 0.00042427999999999997 0 0.00042437999999999997 3.3 0.0004243 3.3 0.0004244 0 0.00042432 0 0.00042442 3.3 0.00042434 3.3 0.00042444 0 0.00042436 0 0.00042446 3.3 0.00042437999999999997 3.3 0.00042448 0 0.0004244 0 0.0004245 3.3 0.00042442 3.3 0.00042452 0 0.00042444 0 0.00042454 3.3 0.00042446 3.3 0.00042456 0 0.00042448 0 0.00042458 3.3 0.00042449999999999996 3.3 0.00042459999999999997 0 0.00042452 0 0.00042462 3.3 0.00042454 3.3 0.00042464 0 0.00042456 0 0.00042466 3.3 0.00042458 3.3 0.00042468 0 0.00042459999999999997 0 0.00042469999999999997 3.3 0.00042462 3.3 0.00042472 0 0.00042464 0 0.00042474 3.3 0.00042466 3.3 0.00042476 0 0.00042468 0 0.00042478 3.3 0.00042469999999999997 3.3 0.00042479999999999997 0 0.00042472 0 0.00042482 3.3 0.00042474 3.3 0.00042484 0 0.00042476 0 0.00042486 3.3 0.00042478 3.3 0.00042488 0 0.00042479999999999997 0 0.0004249 3.3 0.00042482 3.3 0.00042492 0 0.00042484 0 0.00042494 3.3 0.00042486 3.3 0.00042496 0 0.00042488 0 0.00042498 3.3 0.0004249 3.3 0.000425 0 0.00042491999999999996 0 0.00042501999999999997 3.3 0.00042494 3.3 0.00042504 0 0.00042496 0 0.00042506 3.3 0.00042498 3.3 0.00042508 0 0.000425 0 0.0004251 3.3 0.00042501999999999997 3.3 0.00042511999999999997 0 0.00042504 0 0.00042514 3.3 0.00042506 3.3 0.00042516 0 0.00042508 0 0.00042518 3.3 0.0004251 3.3 0.0004252 0 0.00042511999999999997 0 0.00042521999999999997 3.3 0.00042514 3.3 0.00042524 0 0.00042516 0 0.00042526 3.3 0.00042518 3.3 0.00042528 0 0.0004252 0 0.0004253 3.3 0.00042521999999999997 3.3 0.00042532 0 0.00042524 0 0.00042534 3.3 0.00042526 3.3 0.00042536 0 0.00042528 0 0.00042538 3.3 0.0004253 3.3 0.0004254 0 0.00042532 0 0.00042542 3.3 0.00042533999999999996 3.3 0.00042543999999999997 0 0.00042536 0 0.00042546 3.3 0.00042538 3.3 0.00042548 0 0.0004254 0 0.0004255 3.3 0.00042542 3.3 0.00042552 0 0.00042543999999999997 0 0.00042553999999999997 3.3 0.00042546 3.3 0.00042556 0 0.00042548 0 0.00042558 3.3 0.0004255 3.3 0.0004256 0 0.00042552 0 0.00042562 3.3 0.00042553999999999997 3.3 0.00042563999999999997 0 0.00042556 0 0.00042566 3.3 0.00042558 3.3 0.00042568 0 0.0004256 0 0.0004257 3.3 0.00042562 3.3 0.00042572 0 0.00042563999999999997 0 0.00042573999999999997 3.3 0.00042566 3.3 0.00042576 0 0.00042568 0 0.00042578 3.3 0.0004257 3.3 0.0004258 0 0.00042572 0 0.00042582 3.3 0.00042573999999999997 3.3 0.00042584 0 0.00042575999999999996 0 0.00042585999999999996 3.3 0.00042578 3.3 0.00042588 0 0.0004258 0 0.0004259 3.3 0.00042582 3.3 0.00042592 0 0.00042584 0 0.00042594 3.3 0.00042585999999999996 3.3 0.00042595999999999997 0 0.00042588 0 0.00042598 3.3 0.0004259 3.3 0.000426 0 0.00042592 0 0.00042602 3.3 0.00042594 3.3 0.00042604 0 0.00042595999999999997 0 0.00042605999999999997 3.3 0.00042598 3.3 0.00042608 0 0.000426 0 0.0004261 3.3 0.00042602 3.3 0.00042612 0 0.00042604 0 0.00042614 3.3 0.00042605999999999997 3.3 0.00042615999999999997 0 0.00042608 0 0.00042618 3.3 0.0004261 3.3 0.0004262 0 0.00042612 0 0.00042622 3.3 0.00042614 3.3 0.00042624 0 0.00042615999999999997 0 0.00042626 3.3 0.00042618 3.3 0.00042628 0 0.0004262 0 0.0004263 3.3 0.00042622 3.3 0.00042632 0 0.00042624 0 0.00042634 3.3 0.00042626 3.3 0.00042636 0 0.00042627999999999996 0 0.00042637999999999997 3.3 0.0004263 3.3 0.0004264 0 0.00042632 0 0.00042642 3.3 0.00042634 3.3 0.00042644 0 0.00042636 0 0.00042646 3.3 0.00042637999999999997 3.3 0.00042647999999999997 0 0.0004264 0 0.0004265 3.3 0.00042642 3.3 0.00042652 0 0.00042644 0 0.00042654 3.3 0.00042646 3.3 0.00042656 0 0.00042647999999999997 0 0.00042657999999999997 3.3 0.0004265 3.3 0.0004266 0 0.00042652 0 0.00042662 3.3 0.00042654 3.3 0.00042664 0 0.00042656 0 0.00042666 3.3 0.00042657999999999997 3.3 0.00042668 0 0.0004266 0 0.0004267 3.3 0.00042662 3.3 0.00042672 0 0.00042664 0 0.00042674 3.3 0.00042666 3.3 0.00042676 0 0.00042668 0 0.00042678 3.3 0.00042669999999999996 3.3 0.00042679999999999997 0 0.00042672 0 0.00042682 3.3 0.00042674 3.3 0.00042684 0 0.00042676 0 0.00042686 3.3 0.00042678 3.3 0.00042688 0 0.00042679999999999997 0 0.00042689999999999997 3.3 0.00042682 3.3 0.00042692 0 0.00042684 0 0.00042694 3.3 0.00042686 3.3 0.00042696 0 0.00042688 0 0.00042698 3.3 0.00042689999999999997 3.3 0.00042699999999999997 0 0.00042692 0 0.00042702 3.3 0.00042694 3.3 0.00042704 0 0.00042696 0 0.00042706 3.3 0.00042698 3.3 0.00042708 0 0.00042699999999999997 0 0.0004271 3.3 0.00042702 3.3 0.00042712 0 0.00042704 0 0.00042714 3.3 0.00042706 3.3 0.00042716 0 0.00042708 0 0.00042718 3.3 0.0004271 3.3 0.0004272 0 0.00042711999999999996 0 0.00042721999999999997 3.3 0.00042714 3.3 0.00042724 0 0.00042716 0 0.00042726 3.3 0.00042718 3.3 0.00042728 0 0.0004272 0 0.0004273 3.3 0.00042721999999999997 3.3 0.00042731999999999997 0 0.00042724 0 0.00042734 3.3 0.00042726 3.3 0.00042736 0 0.00042728 0 0.00042738 3.3 0.0004273 3.3 0.0004274 0 0.00042731999999999997 0 0.00042741999999999997 3.3 0.00042734 3.3 0.00042744 0 0.00042736 0 0.00042746 3.3 0.00042738 3.3 0.00042748 0 0.0004274 0 0.0004275 3.3 0.00042741999999999997 3.3 0.00042751999999999997 0 0.00042744 0 0.00042754 3.3 0.00042746 3.3 0.00042756 0 0.00042748 0 0.00042758 3.3 0.0004275 3.3 0.0004276 0 0.00042751999999999997 0 0.00042762 3.3 0.00042753999999999996 3.3 0.00042763999999999996 0 0.00042756 0 0.00042766 3.3 0.00042758 3.3 0.00042768 0 0.0004276 0 0.0004277 3.3 0.00042762 3.3 0.00042772 0 0.00042763999999999996 0 0.00042773999999999997 3.3 0.00042766 3.3 0.00042776 0 0.00042768 0 0.00042778 3.3 0.0004277 3.3 0.0004278 0 0.00042772 0 0.00042782 3.3 0.00042773999999999997 3.3 0.00042783999999999997 0 0.00042776 0 0.00042786 3.3 0.00042778 3.3 0.00042788 0 0.0004278 0 0.0004279 3.3 0.00042782 3.3 0.00042792 0 0.00042783999999999997 0 0.00042793999999999997 3.3 0.00042786 3.3 0.00042796 0 0.00042788 0 0.00042798 3.3 0.0004279 3.3 0.000428 0 0.00042792 0 0.00042802 3.3 0.00042793999999999997 3.3 0.00042804 0 0.00042796 0 0.00042806 3.3 0.00042798 3.3 0.00042808 0 0.000428 0 0.0004281 3.3 0.00042802 3.3 0.00042812 0 0.00042804 0 0.00042814 3.3 0.00042805999999999996 3.3 0.00042815999999999997 0 0.00042808 0 0.00042818 3.3 0.0004281 3.3 0.0004282 0 0.00042812 0 0.00042822 3.3 0.00042814 3.3 0.00042824 0 0.00042815999999999997 0 0.00042825999999999997 3.3 0.00042818 3.3 0.00042828 0 0.0004282 0 0.0004283 3.3 0.00042822 3.3 0.00042832 0 0.00042824 0 0.00042834 3.3 0.00042825999999999997 3.3 0.00042835999999999997 0 0.00042828 0 0.00042838 3.3 0.0004283 3.3 0.0004284 0 0.00042832 0 0.00042842 3.3 0.00042834 3.3 0.00042844 0 0.00042835999999999997 0 0.00042846 3.3 0.00042838 3.3 0.00042848 0 0.0004284 0 0.0004285 3.3 0.00042842 3.3 0.00042852 0 0.00042844 0 0.00042854 3.3 0.00042846 3.3 0.00042856 0 0.00042847999999999996 0 0.00042857999999999997 3.3 0.0004285 3.3 0.0004286 0 0.00042852 0 0.00042862 3.3 0.00042854 3.3 0.00042864 0 0.00042856 0 0.00042866 3.3 0.00042857999999999997 3.3 0.00042867999999999997 0 0.0004286 0 0.0004287 3.3 0.00042862 3.3 0.00042872 0 0.00042864 0 0.00042874 3.3 0.00042866 3.3 0.00042876 0 0.00042867999999999997 0 0.00042877999999999997 3.3 0.0004287 3.3 0.0004288 0 0.00042872 0 0.00042882 3.3 0.00042874 3.3 0.00042884 0 0.00042876 0 0.00042886 3.3 0.00042877999999999997 3.3 0.00042888 0 0.0004288 0 0.0004289 3.3 0.00042882 3.3 0.00042892 0 0.00042884 0 0.00042894 3.3 0.00042886 3.3 0.00042896 0 0.00042888 0 0.00042898 3.3 0.00042889999999999996 3.3 0.00042899999999999997 0 0.00042892 0 0.00042902 3.3 0.00042894 3.3 0.00042904 0 0.00042896 0 0.00042906 3.3 0.00042898 3.3 0.00042908 0 0.00042899999999999997 0 0.00042909999999999997 3.3 0.00042902 3.3 0.00042912 0 0.00042904 0 0.00042914 3.3 0.00042906 3.3 0.00042916 0 0.00042908 0 0.00042918 3.3 0.00042909999999999997 3.3 0.00042919999999999997 0 0.00042912 0 0.00042922 3.3 0.00042914 3.3 0.00042924 0 0.00042916 0 0.00042926 3.3 0.00042918 3.3 0.00042928 0 0.00042919999999999997 0 0.00042929999999999997 3.3 0.00042922 3.3 0.00042932 0 0.00042924 0 0.00042934 3.3 0.00042926 3.3 0.00042936 0 0.00042928 0 0.00042938 3.3 0.00042929999999999997 3.3 0.0004294 0 0.00042931999999999996 0 0.00042941999999999996 3.3 0.00042934 3.3 0.00042944 0 0.00042936 0 0.00042946 3.3 0.00042938 3.3 0.00042948 0 0.0004294 0 0.0004295 3.3 0.00042941999999999996 3.3 0.00042951999999999997 0 0.00042944 0 0.00042954 3.3 0.00042946 3.3 0.00042956 0 0.00042948 0 0.00042958 3.3 0.0004295 3.3 0.0004296 0 0.00042951999999999997 0 0.00042961999999999997 3.3 0.00042954 3.3 0.00042964 0 0.00042956 0 0.00042966 3.3 0.00042958 3.3 0.00042968 0 0.0004296 0 0.0004297 3.3 0.00042961999999999997 3.3 0.00042971999999999997 0 0.00042964 0 0.00042974 3.3 0.00042966 3.3 0.00042976 0 0.00042968 0 0.00042978 3.3 0.0004297 3.3 0.0004298 0 0.00042971999999999997 0 0.00042982 3.3 0.00042974 3.3 0.00042984 0 0.00042976 0 0.00042986 3.3 0.00042978 3.3 0.00042988 0 0.0004298 0 0.0004299 3.3 0.00042982 3.3 0.00042992 0 0.00042983999999999996 0 0.00042993999999999997 3.3 0.00042986 3.3 0.00042996 0 0.00042988 0 0.00042998 3.3 0.0004299 3.3 0.00043 0 0.00042992 0 0.00043002 3.3 0.00042993999999999997 3.3 0.00043003999999999997 0 0.00042996 0 0.00043006 3.3 0.00042998 3.3 0.00043008 0 0.00043 0 0.0004301 3.3 0.00043002 3.3 0.00043012 0 0.00043003999999999997 0 0.00043013999999999997 3.3 0.00043006 3.3 0.00043016 0 0.00043008 0 0.00043018 3.3 0.0004301 3.3 0.0004302 0 0.00043012 0 0.00043022 3.3 0.00043013999999999997 3.3 0.00043024 0 0.00043016 0 0.00043026 3.3 0.00043018 3.3 0.00043028 0 0.0004302 0 0.0004303 3.3 0.00043022 3.3 0.00043032 0 0.00043024 0 0.00043034 3.3 0.00043025999999999996 3.3 0.00043035999999999997 0 0.00043028 0 0.00043038 3.3 0.0004303 3.3 0.0004304 0 0.00043032 0 0.00043042 3.3 0.00043034 3.3 0.00043044 0 0.00043035999999999997 0 0.00043045999999999997 3.3 0.00043038 3.3 0.00043048 0 0.0004304 0 0.0004305 3.3 0.00043042 3.3 0.00043052 0 0.00043044 0 0.00043054 3.3 0.00043045999999999997 3.3 0.00043055999999999997 0 0.00043048 0 0.00043058 3.3 0.0004305 3.3 0.0004306 0 0.00043052 0 0.00043062 3.3 0.00043054 3.3 0.00043064 0 0.00043055999999999997 0 0.00043066 3.3 0.00043058 3.3 0.00043068 0 0.0004306 0 0.0004307 3.3 0.00043062 3.3 0.00043072 0 0.00043064 0 0.00043074 3.3 0.00043066 3.3 0.00043076 0 0.00043067999999999996 0 0.00043077999999999997 3.3 0.0004307 3.3 0.0004308 0 0.00043072 0 0.00043082 3.3 0.00043074 3.3 0.00043084 0 0.00043076 0 0.00043086 3.3 0.00043077999999999997 3.3 0.00043087999999999997 0 0.0004308 0 0.0004309 3.3 0.00043082 3.3 0.00043092 0 0.00043084 0 0.00043094 3.3 0.00043086 3.3 0.00043096 0 0.00043087999999999997 0 0.00043097999999999997 3.3 0.0004309 3.3 0.000431 0 0.00043092 0 0.00043102 3.3 0.00043094 3.3 0.00043104 0 0.00043096 0 0.00043106 3.3 0.00043097999999999997 3.3 0.00043107999999999997 0 0.000431 0 0.0004311 3.3 0.00043102 3.3 0.00043112 0 0.00043104 0 0.00043114 3.3 0.00043106 3.3 0.00043116 0 0.00043107999999999997 0 0.00043118 3.3 0.00043109999999999996 3.3 0.00043119999999999996 0 0.00043112 0 0.00043122 3.3 0.00043114 3.3 0.00043124 0 0.00043116 0 0.00043126 3.3 0.00043118 3.3 0.00043128 0 0.00043119999999999996 0 0.00043129999999999997 3.3 0.00043122 3.3 0.00043132 0 0.00043124 0 0.00043134 3.3 0.00043126 3.3 0.00043136 0 0.00043128 0 0.00043138 3.3 0.00043129999999999997 3.3 0.00043139999999999997 0 0.00043132 0 0.00043142 3.3 0.00043134 3.3 0.00043144 0 0.00043136 0 0.00043146 3.3 0.00043138 3.3 0.00043148 0 0.00043139999999999997 0 0.00043149999999999997 3.3 0.00043142 3.3 0.00043152 0 0.00043144 0 0.00043154 3.3 0.00043146 3.3 0.00043156 0 0.00043148 0 0.00043158 3.3 0.00043149999999999997 3.3 0.0004316 0 0.00043152 0 0.00043162 3.3 0.00043154 3.3 0.00043164 0 0.00043156 0 0.00043166 3.3 0.00043158 3.3 0.00043168 0 0.0004316 0 0.0004317 3.3 0.00043161999999999996 3.3 0.00043171999999999997 0 0.00043164 0 0.00043174 3.3 0.00043166 3.3 0.00043176 0 0.00043168 0 0.00043178 3.3 0.0004317 3.3 0.0004318 0 0.00043171999999999997 0 0.00043181999999999997 3.3 0.00043174 3.3 0.00043184 0 0.00043176 0 0.00043186 3.3 0.00043178 3.3 0.00043188 0 0.0004318 0 0.0004319 3.3 0.00043181999999999997 3.3 0.00043191999999999997 0 0.00043184 0 0.00043194 3.3 0.00043186 3.3 0.00043196 0 0.00043188 0 0.00043198 3.3 0.0004319 3.3 0.000432 0 0.00043191999999999997 0 0.00043202 3.3 0.00043194 3.3 0.00043204 0 0.00043196 0 0.00043206 3.3 0.00043198 3.3 0.00043208 0 0.000432 0 0.0004321 3.3 0.00043202 3.3 0.00043212 0 0.00043203999999999996 0 0.00043213999999999997 3.3 0.00043206 3.3 0.00043216 0 0.00043208 0 0.00043218 3.3 0.0004321 3.3 0.0004322 0 0.00043212 0 0.00043222 3.3 0.00043213999999999997 3.3 0.00043223999999999997 0 0.00043216 0 0.00043226 3.3 0.00043218 3.3 0.00043228 0 0.0004322 0 0.0004323 3.3 0.00043222 3.3 0.00043232 0 0.00043223999999999997 0 0.00043233999999999997 3.3 0.00043226 3.3 0.00043236 0 0.00043228 0 0.00043238 3.3 0.0004323 3.3 0.0004324 0 0.00043232 0 0.00043242 3.3 0.00043233999999999997 3.3 0.00043243999999999997 0 0.00043236 0 0.00043246 3.3 0.00043238 3.3 0.00043248 0 0.0004324 0 0.0004325 3.3 0.00043242 3.3 0.00043252 0 0.00043243999999999997 0 0.00043254 3.3 0.00043245999999999996 3.3 0.00043255999999999996 0 0.00043248 0 0.00043258 3.3 0.0004325 3.3 0.0004326 0 0.00043252 0 0.00043262 3.3 0.00043254 3.3 0.00043264 0 0.00043255999999999996 0 0.00043265999999999997 3.3 0.00043258 3.3 0.00043268 0 0.0004326 0 0.0004327 3.3 0.00043262 3.3 0.00043272 0 0.00043264 0 0.00043274 3.3 0.00043265999999999997 3.3 0.00043275999999999997 0 0.00043268 0 0.00043278 3.3 0.0004327 3.3 0.0004328 0 0.00043272 0 0.00043282 3.3 0.00043274 3.3 0.00043284 0 0.00043275999999999997 0 0.00043285999999999997 3.3 0.00043278 3.3 0.00043288 0 0.0004328 0 0.0004329 3.3 0.00043282 3.3 0.00043292 0 0.00043284 0 0.00043294 3.3 0.00043285999999999997 3.3 0.00043296 0 0.00043287999999999996 0 0.00043297999999999996 3.3 0.0004329 3.3 0.000433 0 0.00043292 0 0.00043302 3.3 0.00043294 3.3 0.00043304 0 0.00043296 0 0.00043306 3.3 0.00043297999999999996 3.3 0.00043307999999999997 0 0.000433 0 0.0004331 3.3 0.00043302 3.3 0.00043312 0 0.00043304 0 0.00043314 3.3 0.00043306 3.3 0.00043316 0 0.00043307999999999997 0 0.00043317999999999997 3.3 0.0004331 3.3 0.0004332 0 0.00043312 0 0.00043322 3.3 0.00043314 3.3 0.00043324 0 0.00043316 0 0.00043326 3.3 0.00043317999999999997 3.3 0.00043327999999999997 0 0.0004332 0 0.0004333 3.3 0.00043322 3.3 0.00043332 0 0.00043324 0 0.00043334 3.3 0.00043326 3.3 0.00043336 0 0.00043327999999999997 0 0.00043338 3.3 0.0004333 3.3 0.0004334 0 0.00043332 0 0.00043342 3.3 0.00043334 3.3 0.00043344 0 0.00043336 0 0.00043346 3.3 0.00043338 3.3 0.00043348 0 0.00043339999999999996 0 0.00043349999999999997 3.3 0.00043342 3.3 0.00043352 0 0.00043344 0 0.00043354 3.3 0.00043346 3.3 0.00043356 0 0.00043348 0 0.00043358 3.3 0.00043349999999999997 3.3 0.00043359999999999997 0 0.00043352 0 0.00043362 3.3 0.00043354 3.3 0.00043364 0 0.00043356 0 0.00043366 3.3 0.00043358 3.3 0.00043368 0 0.00043359999999999997 0 0.00043369999999999997 3.3 0.00043362 3.3 0.00043372 0 0.00043364 0 0.00043374 3.3 0.00043366 3.3 0.00043376 0 0.00043368 0 0.00043378 3.3 0.00043369999999999997 3.3 0.0004338 0 0.00043372 0 0.00043382 3.3 0.00043374 3.3 0.00043384 0 0.00043376 0 0.00043386 3.3 0.00043378 3.3 0.00043388 0 0.0004338 0 0.0004339 3.3 0.00043381999999999996 3.3 0.00043391999999999997 0 0.00043384 0 0.00043394 3.3 0.00043386 3.3 0.00043396 0 0.00043388 0 0.00043398 3.3 0.0004339 3.3 0.000434 0 0.00043391999999999997 0 0.00043401999999999997 3.3 0.00043394 3.3 0.00043404 0 0.00043396 0 0.00043406 3.3 0.00043398 3.3 0.00043408 0 0.000434 0 0.0004341 3.3 0.00043401999999999997 3.3 0.00043411999999999997 0 0.00043404 0 0.00043414 3.3 0.00043406 3.3 0.00043416 0 0.00043408 0 0.00043418 3.3 0.0004341 3.3 0.0004342 0 0.00043411999999999997 0 0.00043421999999999997 3.3 0.00043414 3.3 0.00043424 0 0.00043416 0 0.00043426 3.3 0.00043418 3.3 0.00043428 0 0.0004342 0 0.0004343 3.3 0.00043421999999999997 3.3 0.00043432 0 0.00043423999999999996 0 0.00043433999999999996 3.3 0.00043426 3.3 0.00043436 0 0.00043428 0 0.00043438 3.3 0.0004343 3.3 0.0004344 0 0.00043432 0 0.00043442 3.3 0.00043433999999999996 3.3 0.00043443999999999997 0 0.00043436 0 0.00043446 3.3 0.00043438 3.3 0.00043448 0 0.0004344 0 0.0004345 3.3 0.00043442 3.3 0.00043452 0 0.00043443999999999997 0 0.00043453999999999997 3.3 0.00043446 3.3 0.00043456 0 0.00043448 0 0.00043458 3.3 0.0004345 3.3 0.0004346 0 0.00043452 0 0.00043462 3.3 0.00043453999999999997 3.3 0.00043463999999999997 0 0.00043456 0 0.00043466 3.3 0.00043458 3.3 0.00043468 0 0.0004346 0 0.0004347 3.3 0.00043462 3.3 0.00043472 0 0.00043463999999999997 0 0.00043474 3.3 0.00043465999999999996 3.3 0.00043475999999999996 0 0.00043468 0 0.00043478 3.3 0.0004347 3.3 0.0004348 0 0.00043472 0 0.00043482 3.3 0.00043474 3.3 0.00043484 0 0.00043475999999999996 0 0.00043485999999999997 3.3 0.00043478 3.3 0.00043488 0 0.0004348 0 0.0004349 3.3 0.00043482 3.3 0.00043492 0 0.00043484 0 0.00043494 3.3 0.00043485999999999997 3.3 0.00043495999999999997 0 0.00043488 0 0.00043498 3.3 0.0004349 3.3 0.000435 0 0.00043492 0 0.00043502 3.3 0.00043494 3.3 0.00043504 0 0.00043495999999999997 0 0.00043505999999999997 3.3 0.00043498 3.3 0.00043508 0 0.000435 0 0.0004351 3.3 0.00043502 3.3 0.00043512 0 0.00043504 0 0.00043514 3.3 0.00043505999999999997 3.3 0.00043516 0 0.00043508 0 0.00043518 3.3 0.0004351 3.3 0.0004352 0 0.00043512 0 0.00043522 3.3 0.00043514 3.3 0.00043524 0 0.00043516 0 0.00043526 3.3 0.00043517999999999996 3.3 0.00043527999999999997 0 0.0004352 0 0.0004353 3.3 0.00043522 3.3 0.00043532 0 0.00043524 0 0.00043534 3.3 0.00043526 3.3 0.00043536 0 0.00043527999999999997 0 0.00043537999999999997 3.3 0.0004353 3.3 0.0004354 0 0.00043532 0 0.00043542 3.3 0.00043534 3.3 0.00043544 0 0.00043536 0 0.00043546 3.3 0.00043537999999999997 3.3 0.00043547999999999997 0 0.0004354 0 0.0004355 3.3 0.00043542 3.3 0.00043552 0 0.00043544 0 0.00043554 3.3 0.00043546 3.3 0.00043556 0 0.00043547999999999997 0 0.00043558 3.3 0.0004355 3.3 0.0004356 0 0.00043552 0 0.00043562 3.3 0.00043554 3.3 0.00043564 0 0.00043556 0 0.00043566 3.3 0.00043558 3.3 0.00043568 0 0.00043559999999999996 0 0.00043569999999999997 3.3 0.00043562 3.3 0.00043572 0 0.00043564 0 0.00043574 3.3 0.00043566 3.3 0.00043576 0 0.00043568 0 0.00043578 3.3 0.00043569999999999997 3.3 0.00043579999999999997 0 0.00043572 0 0.00043582 3.3 0.00043574 3.3 0.00043584 0 0.00043576 0 0.00043586 3.3 0.00043578 3.3 0.00043588 0 0.00043579999999999997 0 0.00043589999999999997 3.3 0.00043582 3.3 0.00043592 0 0.00043584 0 0.00043594 3.3 0.00043586 3.3 0.00043596 0 0.00043588 0 0.00043598 3.3 0.00043589999999999997 3.3 0.00043599999999999997 0 0.00043592 0 0.00043602 3.3 0.00043594 3.3 0.00043604 0 0.00043596 0 0.00043606 3.3 0.00043598 3.3 0.00043608 0 0.00043599999999999997 0 0.0004361 3.3 0.00043601999999999996 3.3 0.00043611999999999996 0 0.00043604 0 0.00043614 3.3 0.00043606 3.3 0.00043616 0 0.00043608 0 0.00043618 3.3 0.0004361 3.3 0.0004362 0 0.00043611999999999996 0 0.00043621999999999997 3.3 0.00043614 3.3 0.00043624 0 0.00043616 0 0.00043626 3.3 0.00043618 3.3 0.00043628 0 0.0004362 0 0.0004363 3.3 0.00043621999999999997 3.3 0.00043631999999999997 0 0.00043624 0 0.00043634 3.3 0.00043626 3.3 0.00043636 0 0.00043628 0 0.00043638 3.3 0.0004363 3.3 0.0004364 0 0.00043631999999999997 0 0.00043641999999999997 3.3 0.00043634 3.3 0.00043644 0 0.00043636 0 0.00043646 3.3 0.00043638 3.3 0.00043648 0 0.0004364 0 0.0004365 3.3 0.00043641999999999997 3.3 0.00043652 0 0.00043644 0 0.00043654 3.3 0.00043646 3.3 0.00043656 0 0.00043648 0 0.00043658 3.3 0.0004365 3.3 0.0004366 0 0.00043652 0 0.00043662 3.3 0.00043653999999999996 3.3 0.00043663999999999997 0 0.00043656 0 0.00043666 3.3 0.00043658 3.3 0.00043668 0 0.0004366 0 0.0004367 3.3 0.00043662 3.3 0.00043672 0 0.00043663999999999997 0 0.00043673999999999997 3.3 0.00043666 3.3 0.00043676 0 0.00043668 0 0.00043678 3.3 0.0004367 3.3 0.0004368 0 0.00043672 0 0.00043682 3.3 0.00043673999999999997 3.3 0.00043683999999999997 0 0.00043676 0 0.00043686 3.3 0.00043678 3.3 0.00043688 0 0.0004368 0 0.0004369 3.3 0.00043682 3.3 0.00043692 0 0.00043683999999999997 0 0.00043694 3.3 0.00043686 3.3 0.00043696 0 0.00043688 0 0.00043698 3.3 0.0004369 3.3 0.000437 0 0.00043692 0 0.00043702 3.3 0.00043694 3.3 0.00043704 0 0.00043695999999999996 0 0.00043705999999999997 3.3 0.00043698 3.3 0.00043708 0 0.000437 0 0.0004371 3.3 0.00043702 3.3 0.00043712 0 0.00043704 0 0.00043714 3.3 0.00043705999999999997 3.3 0.00043715999999999997 0 0.00043708 0 0.00043718 3.3 0.0004371 3.3 0.0004372 0 0.00043712 0 0.00043722 3.3 0.00043714 3.3 0.00043724 0 0.00043715999999999997 0 0.00043725999999999997 3.3 0.00043718 3.3 0.00043728 0 0.0004372 0 0.0004373 3.3 0.00043722 3.3 0.00043732 0 0.00043724 0 0.00043734 3.3 0.00043725999999999997 3.3 0.00043736 0 0.00043728 0 0.00043738 3.3 0.0004373 3.3 0.0004374 0 0.00043732 0 0.00043742 3.3 0.00043734 3.3 0.00043744 0 0.00043736 0 0.00043746 3.3 0.00043737999999999996 3.3 0.00043747999999999997 0 0.0004374 0 0.0004375 3.3 0.00043742 3.3 0.00043752 0 0.00043744 0 0.00043754 3.3 0.00043746 3.3 0.00043756 0 0.00043747999999999997 0 0.00043757999999999997 3.3 0.0004375 3.3 0.0004376 0 0.00043752 0 0.00043762 3.3 0.00043754 3.3 0.00043764 0 0.00043756 0 0.00043766 3.3 0.00043757999999999997 3.3 0.00043767999999999997 0 0.0004376 0 0.0004377 3.3 0.00043762 3.3 0.00043772 0 0.00043764 0 0.00043774 3.3 0.00043766 3.3 0.00043776 0 0.00043767999999999997 0 0.00043777999999999997 3.3 0.0004377 3.3 0.0004378 0 0.00043772 0 0.00043782 3.3 0.00043774 3.3 0.00043784 0 0.00043776 0 0.00043786 3.3 0.00043777999999999997 3.3 0.00043788 0 0.00043779999999999996 0 0.00043789999999999996 3.3 0.00043782 3.3 0.00043792 0 0.00043784 0 0.00043794 3.3 0.00043786 3.3 0.00043796 0 0.00043788 0 0.00043798 3.3 0.00043789999999999996 3.3 0.00043799999999999997 0 0.00043792 0 0.00043802 3.3 0.00043794 3.3 0.00043804 0 0.00043796 0 0.00043806 3.3 0.00043798 3.3 0.00043808 0 0.00043799999999999997 0 0.00043809999999999997 3.3 0.00043802 3.3 0.00043812 0 0.00043804 0 0.00043814 3.3 0.00043806 3.3 0.00043816 0 0.00043808 0 0.00043818 3.3 0.00043809999999999997 3.3 0.00043819999999999997 0 0.00043812 0 0.00043822 3.3 0.00043814 3.3 0.00043824 0 0.00043816 0 0.00043826 3.3 0.00043818 3.3 0.00043828 0 0.00043819999999999997 0 0.0004383 3.3 0.00043822 3.3 0.00043832 0 0.00043824 0 0.00043834 3.3 0.00043826 3.3 0.00043836 0 0.00043828 0 0.00043838 3.3 0.0004383 3.3 0.0004384 0 0.00043831999999999996 0 0.00043841999999999997 3.3 0.00043834 3.3 0.00043844 0 0.00043836 0 0.00043846 3.3 0.00043838 3.3 0.00043848 0 0.0004384 0 0.0004385 3.3 0.00043841999999999997 3.3 0.00043851999999999997 0 0.00043844 0 0.00043854 3.3 0.00043846 3.3 0.00043856 0 0.00043848 0 0.00043858 3.3 0.0004385 3.3 0.0004386 0 0.00043851999999999997 0 0.00043861999999999997 3.3 0.00043854 3.3 0.00043864 0 0.00043856 0 0.00043866 3.3 0.00043858 3.3 0.00043868 0 0.0004386 0 0.0004387 3.3 0.00043861999999999997 3.3 0.00043872 0 0.00043864 0 0.00043874 3.3 0.00043866 3.3 0.00043876 0 0.00043868 0 0.00043878 3.3 0.0004387 3.3 0.0004388 0 0.00043872 0 0.00043882 3.3 0.00043873999999999996 3.3 0.00043883999999999997 0 0.00043876 0 0.00043886 3.3 0.00043878 3.3 0.00043888 0 0.0004388 0 0.0004389 3.3 0.00043882 3.3 0.00043892 0 0.00043883999999999997 0 0.00043893999999999997 3.3 0.00043886 3.3 0.00043896 0 0.00043888 0 0.00043898 3.3 0.0004389 3.3 0.000439 0 0.00043892 0 0.00043902 3.3 0.00043893999999999997 3.3 0.00043903999999999997 0 0.00043896 0 0.00043906 3.3 0.00043898 3.3 0.00043908 0 0.000439 0 0.0004391 3.3 0.00043902 3.3 0.00043912 0 0.00043903999999999997 0 0.00043914 3.3 0.00043906 3.3 0.00043916 0 0.00043908 0 0.00043918 3.3 0.0004391 3.3 0.0004392 0 0.00043912 0 0.00043922 3.3 0.00043914 3.3 0.00043924 0 0.00043915999999999996 0 0.00043925999999999997 3.3 0.00043918 3.3 0.00043928 0 0.0004392 0 0.0004393 3.3 0.00043922 3.3 0.00043932 0 0.00043924 0 0.00043934 3.3 0.00043925999999999997 3.3 0.00043935999999999997 0 0.00043928 0 0.00043938 3.3 0.0004393 3.3 0.0004394 0 0.00043932 0 0.00043942 3.3 0.00043934 3.3 0.00043944 0 0.00043935999999999997 0 0.00043945999999999997 3.3 0.00043938 3.3 0.00043948 0 0.0004394 0 0.0004395 3.3 0.00043942 3.3 0.00043952 0 0.00043944 0 0.00043954 3.3 0.00043945999999999997 3.3 0.00043955999999999997 0 0.00043948 0 0.00043958 3.3 0.0004395 3.3 0.0004396 0 0.00043952 0 0.00043962 3.3 0.00043954 3.3 0.00043964 0 0.00043955999999999997 0 0.00043966 3.3 0.00043957999999999996 3.3 0.00043967999999999996 0 0.0004396 0 0.0004397 3.3 0.00043962 3.3 0.00043972 0 0.00043964 0 0.00043974 3.3 0.00043966 3.3 0.00043976 0 0.00043967999999999996 0 0.00043977999999999997 3.3 0.0004397 3.3 0.0004398 0 0.00043972 0 0.00043982 3.3 0.00043974 3.3 0.00043984 0 0.00043976 0 0.00043986 3.3 0.00043977999999999997 3.3 0.00043987999999999997 0 0.0004398 0 0.0004399 3.3 0.00043982 3.3 0.00043992 0 0.00043984 0 0.00043994 3.3 0.00043986 3.3 0.00043996 0 0.00043987999999999997 0 0.00043997999999999997 3.3 0.0004399 3.3 0.00044 0 0.00043992 0 0.00044002 3.3 0.00043994 3.3 0.00044004 0 0.00043996 0 0.00044006 3.3 0.00043997999999999997 3.3 0.00044008 0 0.00044 0 0.0004401 3.3 0.00044002 3.3 0.00044012 0 0.00044004 0 0.00044014 3.3 0.00044006 3.3 0.00044016 0 0.00044008 0 0.00044018 3.3 0.00044009999999999996 3.3 0.00044019999999999997 0 0.00044012 0 0.00044022 3.3 0.00044014 3.3 0.00044024 0 0.00044016 0 0.00044026 3.3 0.00044018 3.3 0.00044028 0 0.00044019999999999997 0 0.00044029999999999997 3.3 0.00044022 3.3 0.00044032 0 0.00044024 0 0.00044034 3.3 0.00044026 3.3 0.00044036 0 0.00044028 0 0.00044038 3.3 0.00044029999999999997 3.3 0.00044039999999999997 0 0.00044032 0 0.00044042 3.3 0.00044034 3.3 0.00044044 0 0.00044036 0 0.00044046 3.3 0.00044038 3.3 0.00044048 0 0.00044039999999999997 0 0.0004405 3.3 0.00044042 3.3 0.00044052 0 0.00044044 0 0.00044054 3.3 0.00044046 3.3 0.00044056 0 0.00044048 0 0.00044058 3.3 0.0004405 3.3 0.0004406 0 0.00044051999999999996 0 0.00044061999999999997 3.3 0.00044054 3.3 0.00044064 0 0.00044056 0 0.00044066 3.3 0.00044058 3.3 0.00044068 0 0.0004406 0 0.0004407 3.3 0.00044061999999999997 3.3 0.00044071999999999997 0 0.00044064 0 0.00044074 3.3 0.00044066 3.3 0.00044076 0 0.00044068 0 0.00044078 3.3 0.0004407 3.3 0.0004408 0 0.00044071999999999997 0 0.00044081999999999997 3.3 0.00044074 3.3 0.00044084 0 0.00044076 0 0.00044086 3.3 0.00044078 3.3 0.00044088 0 0.0004408 0 0.0004409 3.3 0.00044081999999999997 3.3 0.00044092 0 0.00044084 0 0.00044094 3.3 0.00044086 3.3 0.00044096 0 0.00044088 0 0.00044098 3.3 0.0004409 3.3 0.000441 0 0.00044092 0 0.00044102 3.3 0.00044093999999999996 3.3 0.00044103999999999997 0 0.00044096 0 0.00044106 3.3 0.00044098 3.3 0.00044108 0 0.000441 0 0.0004411 3.3 0.00044102 3.3 0.00044112 0 0.00044103999999999997 0 0.00044113999999999997 3.3 0.00044106 3.3 0.00044116 0 0.00044108 0 0.00044118 3.3 0.0004411 3.3 0.0004412 0 0.00044112 0 0.00044122 3.3 0.00044113999999999997 3.3 0.00044123999999999997 0 0.00044116 0 0.00044126 3.3 0.00044118 3.3 0.00044128 0 0.0004412 0 0.0004413 3.3 0.00044122 3.3 0.00044132 0 0.00044123999999999997 0 0.00044133999999999997 3.3 0.00044126 3.3 0.00044136 0 0.00044128 0 0.00044138 3.3 0.0004413 3.3 0.0004414 0 0.00044132 0 0.00044142 3.3 0.00044133999999999997 3.3 0.00044144 0 0.00044135999999999996 0 0.00044145999999999996 3.3 0.00044138 3.3 0.00044148 0 0.0004414 0 0.0004415 3.3 0.00044142 3.3 0.00044152 0 0.00044144 0 0.00044154 3.3 0.00044145999999999996 3.3 0.00044155999999999997 0 0.00044148 0 0.00044158 3.3 0.0004415 3.3 0.0004416 0 0.00044152 0 0.00044162 3.3 0.00044154 3.3 0.00044164 0 0.00044155999999999997 0 0.00044165999999999997 3.3 0.00044158 3.3 0.00044168 0 0.0004416 0 0.0004417 3.3 0.00044162 3.3 0.00044172 0 0.00044164 0 0.00044174 3.3 0.00044165999999999997 3.3 0.00044175999999999997 0 0.00044168 0 0.00044178 3.3 0.0004417 3.3 0.0004418 0 0.00044172 0 0.00044182 3.3 0.00044174 3.3 0.00044184 0 0.00044175999999999997 0 0.00044186 3.3 0.00044178 3.3 0.00044188 0 0.0004418 0 0.0004419 3.3 0.00044182 3.3 0.00044192 0 0.00044184 0 0.00044194 3.3 0.00044186 3.3 0.00044196 0 0.00044187999999999996 0 0.00044197999999999997 3.3 0.0004419 3.3 0.000442 0 0.00044192 0 0.00044202 3.3 0.00044194 3.3 0.00044204 0 0.00044196 0 0.00044206 3.3 0.00044197999999999997 3.3 0.00044207999999999997 0 0.000442 0 0.0004421 3.3 0.00044202 3.3 0.00044212 0 0.00044204 0 0.00044214 3.3 0.00044206 3.3 0.00044216 0 0.00044207999999999997 0 0.00044217999999999997 3.3 0.0004421 3.3 0.0004422 0 0.00044212 0 0.00044222 3.3 0.00044214 3.3 0.00044224 0 0.00044216 0 0.00044226 3.3 0.00044217999999999997 3.3 0.00044228 0 0.0004422 0 0.0004423 3.3 0.00044222 3.3 0.00044232 0 0.00044224 0 0.00044234 3.3 0.00044226 3.3 0.00044236 0 0.00044228 0 0.00044238 3.3 0.00044229999999999996 3.3 0.00044239999999999997 0 0.00044232 0 0.00044242 3.3 0.00044234 3.3 0.00044244 0 0.00044236 0 0.00044246 3.3 0.00044238 3.3 0.00044248 0 0.00044239999999999997 0 0.00044249999999999997 3.3 0.00044242 3.3 0.00044252 0 0.00044244 0 0.00044254 3.3 0.00044246 3.3 0.00044256 0 0.00044248 0 0.00044258 3.3 0.00044249999999999997 3.3 0.00044259999999999997 0 0.00044252 0 0.00044262 3.3 0.00044254 3.3 0.00044264 0 0.00044256 0 0.00044266 3.3 0.00044258 3.3 0.00044268 0 0.00044259999999999997 0 0.00044269999999999997 3.3 0.00044262 3.3 0.00044272 0 0.00044264 0 0.00044274 3.3 0.00044266 3.3 0.00044276 0 0.00044268 0 0.00044278 3.3 0.00044269999999999997 3.3 0.0004428 0 0.00044271999999999996 0 0.00044281999999999996 3.3 0.00044274 3.3 0.00044284 0 0.00044276 0 0.00044286 3.3 0.00044278 3.3 0.00044288 0 0.0004428 0 0.0004429 3.3 0.00044281999999999996 3.3 0.00044291999999999997 0 0.00044284 0 0.00044294 3.3 0.00044286 3.3 0.00044296 0 0.00044288 0 0.00044298 3.3 0.0004429 3.3 0.000443 0 0.00044291999999999997 0 0.00044301999999999997 3.3 0.00044294 3.3 0.00044304 0 0.00044296 0 0.00044306 3.3 0.00044298 3.3 0.00044308 0 0.000443 0 0.0004431 3.3 0.00044301999999999997 3.3 0.00044311999999999997 0 0.00044304 0 0.00044314 3.3 0.00044306 3.3 0.00044316 0 0.00044308 0 0.00044318 3.3 0.0004431 3.3 0.0004432 0 0.00044311999999999997 0 0.00044322 3.3 0.00044313999999999996 3.3 0.00044323999999999996 0 0.00044316 0 0.00044326 3.3 0.00044318 3.3 0.00044328 0 0.0004432 0 0.0004433 3.3 0.00044322 3.3 0.00044332 0 0.00044323999999999996 0 0.00044333999999999997 3.3 0.00044326 3.3 0.00044336 0 0.00044328 0 0.00044338 3.3 0.0004433 3.3 0.0004434 0 0.00044332 0 0.00044342 3.3 0.00044333999999999997 3.3 0.00044343999999999997 0 0.00044336 0 0.00044346 3.3 0.00044338 3.3 0.00044348 0 0.0004434 0 0.0004435 3.3 0.00044342 3.3 0.00044352 0 0.00044343999999999997 0 0.00044353999999999997 3.3 0.00044346 3.3 0.00044356 0 0.00044348 0 0.00044358 3.3 0.0004435 3.3 0.0004436 0 0.00044352 0 0.00044362 3.3 0.00044353999999999997 3.3 0.00044364 0 0.00044356 0 0.00044366 3.3 0.00044358 3.3 0.00044368 0 0.0004436 0 0.0004437 3.3 0.00044362 3.3 0.00044372 0 0.00044364 0 0.00044374 3.3 0.00044365999999999996 3.3 0.00044375999999999997 0 0.00044368 0 0.00044378 3.3 0.0004437 3.3 0.0004438 0 0.00044372 0 0.00044382 3.3 0.00044374 3.3 0.00044384 0 0.00044375999999999997 0 0.00044385999999999997 3.3 0.00044378 3.3 0.00044388 0 0.0004438 0 0.0004439 3.3 0.00044382 3.3 0.00044392 0 0.00044384 0 0.00044394 3.3 0.00044385999999999997 3.3 0.00044395999999999997 0 0.00044388 0 0.00044398 3.3 0.0004439 3.3 0.000444 0 0.00044392 0 0.00044402 3.3 0.00044394 3.3 0.00044404 0 0.00044395999999999997 0 0.00044406 3.3 0.00044398 3.3 0.00044408 0 0.000444 0 0.0004441 3.3 0.00044402 3.3 0.00044412 0 0.00044404 0 0.00044414 3.3 0.00044406 3.3 0.00044416 0 0.00044407999999999996 0 0.00044417999999999997 3.3 0.0004441 3.3 0.0004442 0 0.00044412 0 0.00044422 3.3 0.00044414 3.3 0.00044424 0 0.00044416 0 0.00044426 3.3 0.00044417999999999997 3.3 0.00044427999999999997 0 0.0004442 0 0.0004443 3.3 0.00044422 3.3 0.00044432 0 0.00044424 0 0.00044434 3.3 0.00044426 3.3 0.00044436 0 0.00044427999999999997 0 0.00044437999999999997 3.3 0.0004443 3.3 0.0004444 0 0.00044432 0 0.00044442 3.3 0.00044434 3.3 0.00044444 0 0.00044436 0 0.00044446 3.3 0.00044437999999999997 3.3 0.00044447999999999997 0 0.0004444 0 0.0004445 3.3 0.00044442 3.3 0.00044452 0 0.00044444 0 0.00044454 3.3 0.00044446 3.3 0.00044456 0 0.00044447999999999997 0 0.00044458 3.3 0.00044449999999999996 3.3 0.00044459999999999996 0 0.00044452 0 0.00044462 3.3 0.00044454 3.3 0.00044464 0 0.00044456 0 0.00044466 3.3 0.00044458 3.3 0.00044468 0 0.00044459999999999996 0 0.00044469999999999997 3.3 0.00044462 3.3 0.00044472 0 0.00044464 0 0.00044474 3.3 0.00044466 3.3 0.00044476 0 0.00044468 0 0.00044478 3.3 0.00044469999999999997 3.3 0.00044479999999999997 0 0.00044472 0 0.00044482 3.3 0.00044474 3.3 0.00044484 0 0.00044476 0 0.00044486 3.3 0.00044478 3.3 0.00044488 0 0.00044479999999999997 0 0.00044489999999999997 3.3 0.00044482 3.3 0.00044492 0 0.00044484 0 0.00044494 3.3 0.00044486 3.3 0.00044496 0 0.00044488 0 0.00044498 3.3 0.00044489999999999997 3.3 0.000445 0 0.00044491999999999996 0 0.00044501999999999996 3.3 0.00044494 3.3 0.00044504 0 0.00044496 0 0.00044506 3.3 0.00044498 3.3 0.00044508 0 0.000445 0 0.0004451 3.3 0.00044501999999999996 3.3 0.00044511999999999997 0 0.00044504 0 0.00044514 3.3 0.00044506 3.3 0.00044516 0 0.00044508 0 0.00044518 3.3 0.0004451 3.3 0.0004452 0 0.00044511999999999997 0 0.00044521999999999997 3.3 0.00044514 3.3 0.00044524 0 0.00044516 0 0.00044526 3.3 0.00044518 3.3 0.00044528 0 0.0004452 0 0.0004453 3.3 0.00044521999999999997 3.3 0.00044531999999999997 0 0.00044524 0 0.00044534 3.3 0.00044526 3.3 0.00044536 0 0.00044528 0 0.00044538 3.3 0.0004453 3.3 0.0004454 0 0.00044531999999999997 0 0.00044542 3.3 0.00044534 3.3 0.00044544 0 0.00044536 0 0.00044546 3.3 0.00044538 3.3 0.00044548 0 0.0004454 0 0.0004455 3.3 0.00044542 3.3 0.00044552 0 0.00044543999999999996 0 0.00044553999999999997 3.3 0.00044546 3.3 0.00044556 0 0.00044548 0 0.00044558 3.3 0.0004455 3.3 0.0004456 0 0.00044552 0 0.00044562 3.3 0.00044553999999999997 3.3 0.00044563999999999997 0 0.00044556 0 0.00044566 3.3 0.00044558 3.3 0.00044568 0 0.0004456 0 0.0004457 3.3 0.00044562 3.3 0.00044572 0 0.00044563999999999997 0 0.00044573999999999997 3.3 0.00044566 3.3 0.00044576 0 0.00044568 0 0.00044578 3.3 0.0004457 3.3 0.0004458 0 0.00044572 0 0.00044582 3.3 0.00044573999999999997 3.3 0.00044584 0 0.00044576 0 0.00044586 3.3 0.00044578 3.3 0.00044588 0 0.0004458 0 0.0004459 3.3 0.00044582 3.3 0.00044592 0 0.00044584 0 0.00044594 3.3 0.00044585999999999996 3.3 0.00044595999999999997 0 0.00044588 0 0.00044598 3.3 0.0004459 3.3 0.000446 0 0.00044592 0 0.00044602 3.3 0.00044594 3.3 0.00044604 0 0.00044595999999999997 0 0.00044605999999999997 3.3 0.00044598 3.3 0.00044608 0 0.000446 0 0.0004461 3.3 0.00044602 3.3 0.00044612 0 0.00044604 0 0.00044614 3.3 0.00044605999999999997 3.3 0.00044615999999999997 0 0.00044608 0 0.00044618 3.3 0.0004461 3.3 0.0004462 0 0.00044612 0 0.00044622 3.3 0.00044614 3.3 0.00044624 0 0.00044615999999999997 0 0.00044625999999999997 3.3 0.00044618 3.3 0.00044628 0 0.0004462 0 0.0004463 3.3 0.00044622 3.3 0.00044632 0 0.00044624 0 0.00044634 3.3 0.00044625999999999997 3.3 0.00044636 0 0.00044627999999999996 0 0.00044637999999999996 3.3 0.0004463 3.3 0.0004464 0 0.00044632 0 0.00044642 3.3 0.00044634 3.3 0.00044644 0 0.00044636 0 0.00044646 3.3 0.00044637999999999996 3.3 0.00044647999999999997 0 0.0004464 0 0.0004465 3.3 0.00044642 3.3 0.00044652 0 0.00044644 0 0.00044654 3.3 0.00044646 3.3 0.00044656 0 0.00044647999999999997 0 0.00044657999999999997 3.3 0.0004465 3.3 0.0004466 0 0.00044652 0 0.00044662 3.3 0.00044654 3.3 0.00044664 0 0.00044656 0 0.00044666 3.3 0.00044657999999999997 3.3 0.00044667999999999997 0 0.0004466 0 0.0004467 3.3 0.00044662 3.3 0.00044672 0 0.00044664 0 0.00044674 3.3 0.00044666 3.3 0.00044676 0 0.00044667999999999997 0 0.00044678 3.3 0.00044669999999999996 3.3 0.00044679999999999996 0 0.00044672 0 0.00044682 3.3 0.00044674 3.3 0.00044684 0 0.00044676 0 0.00044686 3.3 0.00044678 3.3 0.00044688 0 0.00044679999999999996 0 0.00044689999999999997 3.3 0.00044682 3.3 0.00044692 0 0.00044684 0 0.00044694 3.3 0.00044686 3.3 0.00044696 0 0.00044688 0 0.00044698 3.3 0.00044689999999999997 3.3 0.00044699999999999997 0 0.00044692 0 0.00044702 3.3 0.00044694 3.3 0.00044704 0 0.00044696 0 0.00044706 3.3 0.00044698 3.3 0.00044708 0 0.00044699999999999997 0 0.00044709999999999997 3.3 0.00044702 3.3 0.00044712 0 0.00044704 0 0.00044714 3.3 0.00044706 3.3 0.00044716 0 0.00044708 0 0.00044718 3.3 0.00044709999999999997 3.3 0.0004472 0 0.00044712 0 0.00044722 3.3 0.00044714 3.3 0.00044724 0 0.00044716 0 0.00044726 3.3 0.00044718 3.3 0.00044728 0 0.0004472 0 0.0004473 3.3 0.00044721999999999996 3.3 0.00044731999999999997 0 0.00044724 0 0.00044734 3.3 0.00044726 3.3 0.00044736 0 0.00044728 0 0.00044738 3.3 0.0004473 3.3 0.0004474 0 0.00044731999999999997 0 0.00044741999999999997 3.3 0.00044734 3.3 0.00044744 0 0.00044736 0 0.00044746 3.3 0.00044738 3.3 0.00044748 0 0.0004474 0 0.0004475 3.3 0.00044741999999999997 3.3 0.00044751999999999997 0 0.00044744 0 0.00044754 3.3 0.00044746 3.3 0.00044756 0 0.00044748 0 0.00044758 3.3 0.0004475 3.3 0.0004476 0 0.00044751999999999997 0 0.00044762 3.3 0.00044754 3.3 0.00044764 0 0.00044756 0 0.00044766 3.3 0.00044758 3.3 0.00044768 0 0.0004476 0 0.0004477 3.3 0.00044762 3.3 0.00044772 0 0.00044763999999999996 0 0.00044773999999999997 3.3 0.00044766 3.3 0.00044776 0 0.00044768 0 0.00044778 3.3 0.0004477 3.3 0.0004478 0 0.00044772 0 0.00044782 3.3 0.00044773999999999997 3.3 0.00044783999999999997 0 0.00044776 0 0.00044786 3.3 0.00044778 3.3 0.00044788 0 0.0004478 0 0.0004479 3.3 0.00044782 3.3 0.00044792 0 0.00044783999999999997 0 0.00044793999999999997 3.3 0.00044786 3.3 0.00044796 0 0.00044788 0 0.00044798 3.3 0.0004479 3.3 0.000448 0 0.00044792 0 0.00044802 3.3 0.00044793999999999997 3.3 0.00044803999999999997 0 0.00044796 0 0.00044806 3.3 0.00044798 3.3 0.00044808 0 0.000448 0 0.0004481 3.3 0.00044802 3.3 0.00044812 0 0.00044803999999999997 0 0.00044814 3.3 0.00044805999999999996 3.3 0.00044815999999999996 0 0.00044808 0 0.00044818 3.3 0.0004481 3.3 0.0004482 0 0.00044812 0 0.00044822 3.3 0.00044814 3.3 0.00044824 0 0.00044815999999999996 0 0.00044825999999999997 3.3 0.00044818 3.3 0.00044828 0 0.0004482 0 0.0004483 3.3 0.00044822 3.3 0.00044832 0 0.00044824 0 0.00044834 3.3 0.00044825999999999997 3.3 0.00044835999999999997 0 0.00044828 0 0.00044838 3.3 0.0004483 3.3 0.0004484 0 0.00044832 0 0.00044842 3.3 0.00044834 3.3 0.00044844 0 0.00044835999999999997 0 0.00044845999999999997 3.3 0.00044838 3.3 0.00044848 0 0.0004484 0 0.0004485 3.3 0.00044842 3.3 0.00044852 0 0.00044844 0 0.00044854 3.3 0.00044845999999999997 3.3 0.00044856 0 0.00044847999999999996 0 0.00044857999999999996 3.3 0.0004485 3.3 0.0004486 0 0.00044852 0 0.00044862 3.3 0.00044854 3.3 0.00044864 0 0.00044856 0 0.00044866 3.3 0.00044857999999999996 3.3 0.00044867999999999997 0 0.0004486 0 0.0004487 3.3 0.00044862 3.3 0.00044872 0 0.00044864 0 0.00044874 3.3 0.00044866 3.3 0.00044876 0 0.00044867999999999997 0 0.00044877999999999997 3.3 0.0004487 3.3 0.0004488 0 0.00044872 0 0.00044882 3.3 0.00044874 3.3 0.00044884 0 0.00044876 0 0.00044886 3.3 0.00044877999999999997 3.3 0.00044887999999999997 0 0.0004488 0 0.0004489 3.3 0.00044882 3.3 0.00044892 0 0.00044884 0 0.00044894 3.3 0.00044886 3.3 0.00044896 0 0.00044887999999999997 0 0.00044898 3.3 0.0004489 3.3 0.000449 0 0.00044892 0 0.00044902 3.3 0.00044894 3.3 0.00044904 0 0.00044896 0 0.00044906 3.3 0.00044898 3.3 0.00044908 0 0.00044899999999999996 0 0.00044909999999999997 3.3 0.00044902 3.3 0.00044912 0 0.00044904 0 0.00044914 3.3 0.00044906 3.3 0.00044916 0 0.00044908 0 0.00044918 3.3 0.00044909999999999997 3.3 0.00044919999999999997 0 0.00044912 0 0.00044922 3.3 0.00044914 3.3 0.00044924 0 0.00044916 0 0.00044926 3.3 0.00044918 3.3 0.00044928 0 0.00044919999999999997 0 0.00044929999999999997 3.3 0.00044922 3.3 0.00044932 0 0.00044924 0 0.00044934 3.3 0.00044926 3.3 0.00044936 0 0.00044928 0 0.00044938 3.3 0.00044929999999999997 3.3 0.0004494 0 0.00044932 0 0.00044942 3.3 0.00044934 3.3 0.00044944 0 0.00044936 0 0.00044946 3.3 0.00044938 3.3 0.00044948 0 0.0004494 0 0.0004495 3.3 0.00044941999999999996 3.3 0.00044951999999999997 0 0.00044944 0 0.00044954 3.3 0.00044946 3.3 0.00044956 0 0.00044948 0 0.00044958 3.3 0.0004495 3.3 0.0004496 0 0.00044951999999999997 0 0.00044961999999999997 3.3 0.00044954 3.3 0.00044964 0 0.00044956 0 0.00044966 3.3 0.00044958 3.3 0.00044968 0 0.0004496 0 0.0004497 3.3 0.00044961999999999997 3.3 0.00044971999999999997 0 0.00044964 0 0.00044974 3.3 0.00044966 3.3 0.00044976 0 0.00044968 0 0.00044978 3.3 0.0004497 3.3 0.0004498 0 0.00044971999999999997 0 0.00044981999999999997 3.3 0.00044974 3.3 0.00044984 0 0.00044976 0 0.00044986 3.3 0.00044978 3.3 0.00044988 0 0.0004498 0 0.0004499 3.3 0.00044981999999999997 3.3 0.00044992 0 0.00044983999999999996 0 0.00044993999999999996 3.3 0.00044986 3.3 0.00044996 0 0.00044988 0 0.00044998 3.3 0.0004499 3.3 0.00045 0 0.00044992 0 0.00045002 3.3 0.00044993999999999996 3.3 0.00045003999999999997 0 0.00044996 0 0.00045006 3.3 0.00044998 3.3 0.00045008 0 0.00045 0 0.0004501 3.3 0.00045002 3.3 0.00045012 0 0.00045003999999999997 0 0.00045013999999999997 3.3 0.00045006 3.3 0.00045016 0 0.00045008 0 0.00045018 3.3 0.0004501 3.3 0.0004502 0 0.00045012 0 0.00045022 3.3 0.00045013999999999997 3.3 0.00045023999999999997 0 0.00045016 0 0.00045026 3.3 0.00045018 3.3 0.00045028 0 0.0004502 0 0.0004503 3.3 0.00045022 3.3 0.00045032 0 0.00045023999999999997 0 0.00045034 3.3 0.00045025999999999996 3.3 0.00045035999999999996 0 0.00045028 0 0.00045038 3.3 0.0004503 3.3 0.0004504 0 0.00045032 0 0.00045042 3.3 0.00045034 3.3 0.00045044 0 0.00045035999999999996 0 0.00045045999999999997 3.3 0.00045038 3.3 0.00045048 0 0.0004504 0 0.0004505 3.3 0.00045042 3.3 0.00045052 0 0.00045044 0 0.00045054 3.3 0.00045045999999999997 3.3 0.00045055999999999997 0 0.00045048 0 0.00045058 3.3 0.0004505 3.3 0.0004506 0 0.00045052 0 0.00045062 3.3 0.00045054 3.3 0.00045064 0 0.00045055999999999997 0 0.00045065999999999997 3.3 0.00045058 3.3 0.00045068 0 0.0004506 0 0.0004507 3.3 0.00045062 3.3 0.00045072 0 0.00045064 0 0.00045074 3.3 0.00045065999999999997 3.3 0.00045076 0 0.00045068 0 0.00045078 3.3 0.0004507 3.3 0.0004508 0 0.00045072 0 0.00045082 3.3 0.00045074 3.3 0.00045084 0 0.00045076 0 0.00045086 3.3 0.00045077999999999996 3.3 0.00045087999999999997 0 0.0004508 0 0.0004509 3.3 0.00045082 3.3 0.00045092 0 0.00045084 0 0.00045094 3.3 0.00045086 3.3 0.00045096 0 0.00045087999999999997 0 0.00045097999999999997 3.3 0.0004509 3.3 0.000451 0 0.00045092 0 0.00045102 3.3 0.00045094 3.3 0.00045104 0 0.00045096 0 0.00045106 3.3 0.00045097999999999997 3.3 0.00045107999999999997 0 0.000451 0 0.0004511 3.3 0.00045102 3.3 0.00045112 0 0.00045104 0 0.00045114 3.3 0.00045106 3.3 0.00045116 0 0.00045107999999999997 0 0.00045118 3.3 0.0004511 3.3 0.0004512 0 0.00045112 0 0.00045122 3.3 0.00045114 3.3 0.00045124 0 0.00045116 0 0.00045126 3.3 0.00045118 3.3 0.00045128 0 0.00045119999999999996 0 0.00045129999999999997 3.3 0.00045122 3.3 0.00045132 0 0.00045124 0 0.00045134 3.3 0.00045126 3.3 0.00045136 0 0.00045128 0 0.00045138 3.3 0.00045129999999999997 3.3 0.00045139999999999997 0 0.00045132 0 0.00045142 3.3 0.00045134 3.3 0.00045144 0 0.00045136 0 0.00045146 3.3 0.00045138 3.3 0.00045148 0 0.00045139999999999997 0 0.00045149999999999997 3.3 0.00045142 3.3 0.00045152 0 0.00045144 0 0.00045154 3.3 0.00045146 3.3 0.00045156 0 0.00045148 0 0.00045158 3.3 0.00045149999999999997 3.3 0.00045159999999999997 0 0.00045152 0 0.00045162 3.3 0.00045154 3.3 0.00045164 0 0.00045156 0 0.00045166 3.3 0.00045158 3.3 0.00045168 0 0.00045159999999999997 0 0.0004517 3.3 0.00045161999999999996 3.3 0.00045171999999999996 0 0.00045164 0 0.00045174 3.3 0.00045166 3.3 0.00045176 0 0.00045168 0 0.00045178 3.3 0.0004517 3.3 0.0004518 0 0.00045171999999999996 0 0.00045181999999999997 3.3 0.00045174 3.3 0.00045184 0 0.00045176 0 0.00045186 3.3 0.00045178 3.3 0.00045188 0 0.0004518 0 0.0004519 3.3 0.00045181999999999997 3.3 0.00045191999999999997 0 0.00045184 0 0.00045194 3.3 0.00045186 3.3 0.00045196 0 0.00045188 0 0.00045198 3.3 0.0004519 3.3 0.000452 0 0.00045191999999999997 0 0.00045201999999999997 3.3 0.00045194 3.3 0.00045204 0 0.00045196 0 0.00045206 3.3 0.00045198 3.3 0.00045208 0 0.000452 0 0.0004521 3.3 0.00045201999999999997 3.3 0.00045212 0 0.00045203999999999996 0 0.00045213999999999996 3.3 0.00045206 3.3 0.00045216 0 0.00045208 0 0.00045218 3.3 0.0004521 3.3 0.0004522 0 0.00045212 0 0.00045222 3.3 0.00045213999999999996 3.3 0.00045223999999999997 0 0.00045216 0 0.00045226 3.3 0.00045218 3.3 0.00045228 0 0.0004522 0 0.0004523 3.3 0.00045222 3.3 0.00045232 0 0.00045223999999999997 0 0.00045233999999999997 3.3 0.00045226 3.3 0.00045236 0 0.00045228 0 0.00045238 3.3 0.0004523 3.3 0.0004524 0 0.00045232 0 0.00045242 3.3 0.00045233999999999997 3.3 0.00045243999999999997 0 0.00045236 0 0.00045246 3.3 0.00045238 3.3 0.00045248 0 0.0004524 0 0.0004525 3.3 0.00045242 3.3 0.00045252 0 0.00045243999999999997 0 0.00045254 3.3 0.00045246 3.3 0.00045256 0 0.00045248 0 0.00045258 3.3 0.0004525 3.3 0.0004526 0 0.00045252 0 0.00045262 3.3 0.00045254 3.3 0.00045264 0 0.00045255999999999996 0 0.00045265999999999997 3.3 0.00045258 3.3 0.00045268 0 0.0004526 0 0.0004527 3.3 0.00045262 3.3 0.00045272 0 0.00045264 0 0.00045274 3.3 0.00045265999999999997 3.3 0.00045275999999999997 0 0.00045268 0 0.00045278 3.3 0.0004527 3.3 0.0004528 0 0.00045272 0 0.00045282 3.3 0.00045274 3.3 0.00045284 0 0.00045275999999999997 0 0.00045285999999999997 3.3 0.00045278 3.3 0.00045288 0 0.0004528 0 0.0004529 3.3 0.00045282 3.3 0.00045292 0 0.00045284 0 0.00045294 3.3 0.00045285999999999997 3.3 0.00045296 0 0.00045288 0 0.00045298 3.3 0.0004529 3.3 0.000453 0 0.00045292 0 0.00045302 3.3 0.00045294 3.3 0.00045304 0 0.00045296 0 0.00045306 3.3 0.00045297999999999996 3.3 0.00045307999999999996 0 0.000453 0 0.0004531 3.3 0.00045302 3.3 0.00045312 0 0.00045304 0 0.00045314 3.3 0.00045306 3.3 0.00045316 0 0.00045307999999999996 0 0.00045317999999999997 3.3 0.0004531 3.3 0.0004532 0 0.00045312 0 0.00045322 3.3 0.00045314 3.3 0.00045324 0 0.00045316 0 0.00045326 3.3 0.00045317999999999997 3.3 0.00045327999999999997 0 0.0004532 0 0.0004533 3.3 0.00045322 3.3 0.00045332 0 0.00045324 0 0.00045334 3.3 0.00045326 3.3 0.00045336 0 0.00045327999999999997 0 0.00045337999999999997 3.3 0.0004533 3.3 0.0004534 0 0.00045332 0 0.00045342 3.3 0.00045334 3.3 0.00045344 0 0.00045336 0 0.00045346 3.3 0.00045337999999999997 3.3 0.00045348 0 0.00045339999999999996 0 0.00045349999999999996 3.3 0.00045342 3.3 0.00045352 0 0.00045344 0 0.00045354 3.3 0.00045346 3.3 0.00045356 0 0.00045348 0 0.00045358 3.3 0.00045349999999999996 3.3 0.00045359999999999997 0 0.00045352 0 0.00045362 3.3 0.00045354 3.3 0.00045364 0 0.00045356 0 0.00045366 3.3 0.00045358 3.3 0.00045368 0 0.00045359999999999997 0 0.00045369999999999997 3.3 0.00045362 3.3 0.00045372 0 0.00045364 0 0.00045374 3.3 0.00045366 3.3 0.00045376 0 0.00045368 0 0.00045378 3.3 0.00045369999999999997 3.3 0.00045379999999999997 0 0.00045372 0 0.00045382 3.3 0.00045374 3.3 0.00045384 0 0.00045376 0 0.00045386 3.3 0.00045378 3.3 0.00045388 0 0.00045379999999999997 0 0.0004539 3.3 0.00045382 3.3 0.00045392 0 0.00045384 0 0.00045394 3.3 0.00045386 3.3 0.00045396 0 0.00045388 0 0.00045398 3.3 0.0004539 3.3 0.000454 0 0.00045391999999999996 0 0.00045401999999999997 3.3 0.00045394 3.3 0.00045404 0 0.00045396 0 0.00045406 3.3 0.00045398 3.3 0.00045408 0 0.000454 0 0.0004541 3.3 0.00045401999999999997 3.3 0.00045411999999999997 0 0.00045404 0 0.00045414 3.3 0.00045406 3.3 0.00045416 0 0.00045408 0 0.00045418 3.3 0.0004541 3.3 0.0004542 0 0.00045411999999999997 0 0.00045421999999999997 3.3 0.00045414 3.3 0.00045424 0 0.00045416 0 0.00045426 3.3 0.00045418 3.3 0.00045428 0 0.0004542 0 0.0004543 3.3 0.00045421999999999997 3.3 0.00045432 0 0.00045424 0 0.00045434 3.3 0.00045426 3.3 0.00045436 0 0.00045428 0 0.00045438 3.3 0.0004543 3.3 0.0004544 0 0.00045432 0 0.00045442 3.3 0.00045433999999999996 3.3 0.00045443999999999997 0 0.00045436 0 0.00045446 3.3 0.00045438 3.3 0.00045448 0 0.0004544 0 0.0004545 3.3 0.00045442 3.3 0.00045452 0 0.00045443999999999997 0 0.00045453999999999997 3.3 0.00045446 3.3 0.00045456 0 0.00045448 0 0.00045458 3.3 0.0004545 3.3 0.0004546 0 0.00045452 0 0.00045462 3.3 0.00045453999999999997 3.3 0.00045463999999999997 0 0.00045456 0 0.00045466 3.3 0.00045458 3.3 0.00045468 0 0.0004546 0 0.0004547 3.3 0.00045462 3.3 0.00045472 0 0.00045463999999999997 0 0.00045473999999999997 3.3 0.00045466 3.3 0.00045476 0 0.00045468 0 0.00045478 3.3 0.0004547 3.3 0.0004548 0 0.00045472 0 0.00045482 3.3 0.00045473999999999997 3.3 0.00045484 0 0.00045475999999999996 0 0.00045485999999999996 3.3 0.00045478 3.3 0.00045488 0 0.0004548 0 0.0004549 3.3 0.00045482 3.3 0.00045492 0 0.00045484 0 0.00045494 3.3 0.00045485999999999996 3.3 0.00045495999999999997 0 0.00045488 0 0.00045498 3.3 0.0004549 3.3 0.000455 0 0.00045492 0 0.00045502 3.3 0.00045494 3.3 0.00045504 0 0.00045495999999999997 0 0.00045505999999999997 3.3 0.00045498 3.3 0.00045508 0 0.000455 0 0.0004551 3.3 0.00045502 3.3 0.00045512 0 0.00045504 0 0.00045514 3.3 0.00045505999999999997 3.3 0.00045515999999999997 0 0.00045508 0 0.00045518 3.3 0.0004551 3.3 0.0004552 0 0.00045512 0 0.00045522 3.3 0.00045514 3.3 0.00045524 0 0.00045515999999999997 0 0.00045526 3.3 0.00045517999999999996 3.3 0.00045527999999999996 0 0.0004552 0 0.0004553 3.3 0.00045522 3.3 0.00045532 0 0.00045524 0 0.00045534 3.3 0.00045526 3.3 0.00045536 0 0.00045527999999999996 0 0.00045537999999999997 3.3 0.0004553 3.3 0.0004554 0 0.00045532 0 0.00045542 3.3 0.00045534 3.3 0.00045544 0 0.00045536 0 0.00045546 3.3 0.00045537999999999997 3.3 0.00045547999999999997 0 0.0004554 0 0.0004555 3.3 0.00045542 3.3 0.00045552 0 0.00045544 0 0.00045554 3.3 0.00045546 3.3 0.00045556 0 0.00045547999999999997 0 0.00045557999999999997 3.3 0.0004555 3.3 0.0004556 0 0.00045552 0 0.00045562 3.3 0.00045554 3.3 0.00045564 0 0.00045556 0 0.00045566 3.3 0.00045557999999999997 3.3 0.00045568 0 0.0004556 0 0.0004557 3.3 0.00045562 3.3 0.00045572 0 0.00045564 0 0.00045574 3.3 0.00045566 3.3 0.00045576 0 0.00045568 0 0.00045578 3.3 0.00045569999999999996 3.3 0.00045579999999999997 0 0.00045572 0 0.00045582 3.3 0.00045574 3.3 0.00045584 0 0.00045576 0 0.00045586 3.3 0.00045578 3.3 0.00045588 0 0.00045579999999999997 0 0.00045589999999999997 3.3 0.00045582 3.3 0.00045592 0 0.00045584 0 0.00045594 3.3 0.00045586 3.3 0.00045596 0 0.00045588 0 0.00045598 3.3 0.00045589999999999997 3.3 0.00045599999999999997 0 0.00045592 0 0.00045602 3.3 0.00045594 3.3 0.00045604 0 0.00045596 0 0.00045606 3.3 0.00045598 3.3 0.00045608 0 0.00045599999999999997 0 0.0004561 3.3 0.00045602 3.3 0.00045612 0 0.00045604 0 0.00045614 3.3 0.00045606 3.3 0.00045616 0 0.00045608 0 0.00045618 3.3 0.0004561 3.3 0.0004562 0 0.00045611999999999996 0 0.00045621999999999997 3.3 0.00045614 3.3 0.00045624 0 0.00045616 0 0.00045626 3.3 0.00045618 3.3 0.00045628 0 0.0004562 0 0.0004563 3.3 0.00045621999999999997 3.3 0.00045631999999999997 0 0.00045624 0 0.00045634 3.3 0.00045626 3.3 0.00045636 0 0.00045628 0 0.00045638 3.3 0.0004563 3.3 0.0004564 0 0.00045631999999999997 0 0.00045641999999999997 3.3 0.00045634 3.3 0.00045644 0 0.00045636 0 0.00045646 3.3 0.00045638 3.3 0.00045648 0 0.0004564 0 0.0004565 3.3 0.00045641999999999997 3.3 0.00045651999999999997 0 0.00045644 0 0.00045654 3.3 0.00045646 3.3 0.00045656 0 0.00045648 0 0.00045658 3.3 0.0004565 3.3 0.0004566 0 0.00045651999999999997 0 0.00045662 3.3 0.00045653999999999996 3.3 0.00045663999999999996 0 0.00045656 0 0.00045666 3.3 0.00045658 3.3 0.00045668 0 0.0004566 0 0.0004567 3.3 0.00045662 3.3 0.00045672 0 0.00045663999999999996 0 0.00045673999999999997 3.3 0.00045666 3.3 0.00045676 0 0.00045668 0 0.00045678 3.3 0.0004567 3.3 0.0004568 0 0.00045672 0 0.00045682 3.3 0.00045673999999999997 3.3 0.00045683999999999997 0 0.00045676 0 0.00045686 3.3 0.00045678 3.3 0.00045688 0 0.0004568 0 0.0004569 3.3 0.00045682 3.3 0.00045692 0 0.00045683999999999997 0 0.00045693999999999997 3.3 0.00045686 3.3 0.00045696 0 0.00045688 0 0.00045698 3.3 0.0004569 3.3 0.000457 0 0.00045692 0 0.00045702 3.3 0.00045693999999999997 3.3 0.00045704 0 0.00045695999999999996 0 0.00045705999999999996 3.3 0.00045698 3.3 0.00045708 0 0.000457 0 0.0004571 3.3 0.00045702 3.3 0.00045712 0 0.00045704 0 0.00045714 3.3 0.00045705999999999996 3.3 0.00045715999999999997 0 0.00045708 0 0.00045718 3.3 0.0004571 3.3 0.0004572 0 0.00045712 0 0.00045722 3.3 0.00045714 3.3 0.00045724 0 0.00045715999999999997 0 0.00045725999999999997 3.3 0.00045718 3.3 0.00045728 0 0.0004572 0 0.0004573 3.3 0.00045722 3.3 0.00045732 0 0.00045724 0 0.00045734 3.3 0.00045725999999999997 3.3 0.00045735999999999997 0 0.00045728 0 0.00045738 3.3 0.0004573 3.3 0.0004574 0 0.00045732 0 0.00045742 3.3 0.00045734 3.3 0.00045744 0 0.00045735999999999997 0 0.00045746 3.3 0.00045738 3.3 0.00045748 0 0.0004574 0 0.0004575 3.3 0.00045742 3.3 0.00045752 0 0.00045744 0 0.00045754 3.3 0.00045746 3.3 0.00045756 0 0.00045747999999999996 0 0.00045757999999999997 3.3 0.0004575 3.3 0.0004576 0 0.00045752 0 0.00045762 3.3 0.00045754 3.3 0.00045764 0 0.00045756 0 0.00045766 3.3 0.00045757999999999997 3.3 0.00045767999999999997 0 0.0004576 0 0.0004577 3.3 0.00045762 3.3 0.00045772 0 0.00045764 0 0.00045774 3.3 0.00045766 3.3 0.00045776 0 0.00045767999999999997 0 0.00045777999999999997 3.3 0.0004577 3.3 0.0004578 0 0.00045772 0 0.00045782 3.3 0.00045774 3.3 0.00045784 0 0.00045776 0 0.00045786 3.3 0.00045777999999999997 3.3 0.00045788 0 0.0004578 0 0.0004579 3.3 0.00045782 3.3 0.00045792 0 0.00045784 0 0.00045794 3.3 0.00045786 3.3 0.00045796 0 0.00045788 0 0.00045798 3.3 0.00045789999999999996 3.3 0.00045799999999999997 0 0.00045792 0 0.00045802 3.3 0.00045794 3.3 0.00045804 0 0.00045796 0 0.00045806 3.3 0.00045798 3.3 0.00045808 0 0.00045799999999999997 0 0.00045809999999999997 3.3 0.00045802 3.3 0.00045812 0 0.00045804 0 0.00045814 3.3 0.00045806 3.3 0.00045816 0 0.00045808 0 0.00045818 3.3 0.00045809999999999997 3.3 0.00045819999999999997 0 0.00045812 0 0.00045822 3.3 0.00045814 3.3 0.00045824 0 0.00045816 0 0.00045826 3.3 0.00045818 3.3 0.00045828 0 0.00045819999999999997 0 0.00045829999999999997 3.3 0.00045822 3.3 0.00045832 0 0.00045824 0 0.00045834 3.3 0.00045826 3.3 0.00045836 0 0.00045828 0 0.00045838 3.3 0.00045829999999999997 3.3 0.0004584 0 0.00045831999999999996 0 0.00045841999999999996 3.3 0.00045834 3.3 0.00045844 0 0.00045836 0 0.00045846 3.3 0.00045838 3.3 0.00045848 0 0.0004584 0 0.0004585 3.3 0.00045841999999999996 3.3 0.00045851999999999997 0 0.00045844 0 0.00045854 3.3 0.00045846 3.3 0.00045856 0 0.00045848 0 0.00045858 3.3 0.0004585 3.3 0.0004586 0 0.00045851999999999997 0 0.00045861999999999997 3.3 0.00045854 3.3 0.00045864 0 0.00045856 0 0.00045866 3.3 0.00045858 3.3 0.00045868 0 0.0004586 0 0.0004587 3.3 0.00045861999999999997 3.3 0.00045871999999999997 0 0.00045864 0 0.00045874 3.3 0.00045866 3.3 0.00045876 0 0.00045868 0 0.00045878 3.3 0.0004587 3.3 0.0004588 0 0.00045871999999999997 0 0.00045882 3.3 0.00045873999999999996 3.3 0.00045883999999999996 0 0.00045876 0 0.00045886 3.3 0.00045878 3.3 0.00045888 0 0.0004588 0 0.0004589 3.3 0.00045882 3.3 0.00045892 0 0.00045883999999999996 0 0.00045893999999999997 3.3 0.00045886 3.3 0.00045896 0 0.00045888 0 0.00045898 3.3 0.0004589 3.3 0.000459 0 0.00045892 0 0.00045902 3.3 0.00045893999999999997 3.3 0.00045903999999999997 0 0.00045896 0 0.00045906 3.3 0.00045898 3.3 0.00045908 0 0.000459 0 0.0004591 3.3 0.00045902 3.3 0.00045912 0 0.00045903999999999997 0 0.00045913999999999997 3.3 0.00045906 3.3 0.00045916 0 0.00045908 0 0.00045918 3.3 0.0004591 3.3 0.0004592 0 0.00045912 0 0.00045922 3.3 0.00045913999999999997 3.3 0.00045924 0 0.00045916 0 0.00045926 3.3 0.00045918 3.3 0.00045928 0 0.0004592 0 0.0004593 3.3 0.00045922 3.3 0.00045932 0 0.00045924 0 0.00045934 3.3 0.00045925999999999996 3.3 0.00045935999999999997 0 0.00045928 0 0.00045938 3.3 0.0004593 3.3 0.0004594 0 0.00045932 0 0.00045942 3.3 0.00045934 3.3 0.00045944 0 0.00045935999999999997 0 0.00045945999999999997 3.3 0.00045938 3.3 0.00045948 0 0.0004594 0 0.0004595 3.3 0.00045942 3.3 0.00045952 0 0.00045944 0 0.00045954 3.3 0.00045945999999999997 3.3 0.00045955999999999997 0 0.00045948 0 0.00045958 3.3 0.0004595 3.3 0.0004596 0 0.00045952 0 0.00045962 3.3 0.00045954 3.3 0.00045964 0 0.00045955999999999997 0 0.00045966 3.3 0.00045958 3.3 0.00045968 0 0.0004596 0 0.0004597 3.3 0.00045962 3.3 0.00045972 0 0.00045964 0 0.00045974 3.3 0.00045966 3.3 0.00045976 0 0.00045967999999999996 0 0.00045977999999999997 3.3 0.0004597 3.3 0.0004598 0 0.00045972 0 0.00045982 3.3 0.00045974 3.3 0.00045984 0 0.00045976 0 0.00045986 3.3 0.00045977999999999997 3.3 0.00045987999999999997 0 0.0004598 0 0.0004599 3.3 0.00045982 3.3 0.00045992 0 0.00045984 0 0.00045994 3.3 0.00045986 3.3 0.00045996 0 0.00045987999999999997 0 0.00045997999999999997 3.3 0.0004599 3.3 0.00046 0 0.00045992 0 0.00046002 3.3 0.00045994 3.3 0.00046004 0 0.00045996 0 0.00046006 3.3 0.00045997999999999997 3.3 0.00046007999999999997 0 0.00046 0 0.0004601 3.3 0.00046002 3.3 0.00046012 0 0.00046004 0 0.00046014 3.3 0.00046006 3.3 0.00046016 0 0.00046007999999999997 0 0.00046018 3.3 0.00046009999999999996 3.3 0.00046019999999999996 0 0.00046012 0 0.00046022 3.3 0.00046014 3.3 0.00046024 0 0.00046016 0 0.00046026 3.3 0.00046018 3.3 0.00046028 0 0.00046019999999999996 0 0.00046029999999999997 3.3 0.00046022 3.3 0.00046032 0 0.00046024 0 0.00046034 3.3 0.00046026 3.3 0.00046036 0 0.00046028 0 0.00046038 3.3 0.00046029999999999997 3.3 0.00046039999999999997 0 0.00046032 0 0.00046042 3.3 0.00046034 3.3 0.00046044 0 0.00046036 0 0.00046046 3.3 0.00046038 3.3 0.00046048 0 0.00046039999999999997 0 0.00046049999999999997 3.3 0.00046042 3.3 0.00046052 0 0.00046044 0 0.00046054 3.3 0.00046046 3.3 0.00046056 0 0.00046048 0 0.00046058 3.3 0.00046049999999999997 3.3 0.0004606 0 0.00046051999999999996 0 0.00046061999999999996 3.3 0.00046054 3.3 0.00046064 0 0.00046056 0 0.00046066 3.3 0.00046058 3.3 0.00046068 0 0.0004606 0 0.0004607 3.3 0.00046061999999999996 3.3 0.00046071999999999997 0 0.00046064 0 0.00046074 3.3 0.00046066 3.3 0.00046076 0 0.00046068 0 0.00046078 3.3 0.0004607 3.3 0.0004608 0 0.00046071999999999997 0 0.00046081999999999997 3.3 0.00046074 3.3 0.00046084 0 0.00046076 0 0.00046086 3.3 0.00046078 3.3 0.00046088 0 0.0004608 0 0.0004609 3.3 0.00046081999999999997 3.3 0.00046091999999999997 0 0.00046084 0 0.00046094 3.3 0.00046086 3.3 0.00046096 0 0.00046088 0 0.00046098 3.3 0.0004609 3.3 0.000461 0 0.00046091999999999997 0 0.00046102 3.3 0.00046094 3.3 0.00046104 0 0.00046096 0 0.00046106 3.3 0.00046098 3.3 0.00046108 0 0.000461 0 0.0004611 3.3 0.00046102 3.3 0.00046112 0 0.00046103999999999996 0 0.00046113999999999997 3.3 0.00046106 3.3 0.00046116 0 0.00046108 0 0.00046118 3.3 0.0004611 3.3 0.0004612 0 0.00046112 0 0.00046122 3.3 0.00046113999999999997 3.3 0.00046123999999999997 0 0.00046116 0 0.00046126 3.3 0.00046118 3.3 0.00046128 0 0.0004612 0 0.0004613 3.3 0.00046122 3.3 0.00046132 0 0.00046123999999999997 0 0.00046133999999999997 3.3 0.00046126 3.3 0.00046136 0 0.00046128 0 0.00046138 3.3 0.0004613 3.3 0.0004614 0 0.00046132 0 0.00046142 3.3 0.00046133999999999997 3.3 0.00046144 0 0.00046136 0 0.00046146 3.3 0.00046138 3.3 0.00046148 0 0.0004614 0 0.0004615 3.3 0.00046142 3.3 0.00046152 0 0.00046144 0 0.00046154 3.3 0.00046145999999999996 3.3 0.00046155999999999997 0 0.00046148 0 0.00046158 3.3 0.0004615 3.3 0.0004616 0 0.00046152 0 0.00046162 3.3 0.00046154 3.3 0.00046164 0 0.00046155999999999997 0 0.00046165999999999997 3.3 0.00046158 3.3 0.00046168 0 0.0004616 0 0.0004617 3.3 0.00046162 3.3 0.00046172 0 0.00046164 0 0.00046174 3.3 0.00046165999999999997 3.3 0.00046175999999999997 0 0.00046168 0 0.00046178 3.3 0.0004617 3.3 0.0004618 0 0.00046172 0 0.00046182 3.3 0.00046174 3.3 0.00046184 0 0.00046175999999999997 0 0.00046185999999999997 3.3 0.00046178 3.3 0.00046188 0 0.0004618 0 0.0004619 3.3 0.00046182 3.3 0.00046192 0 0.00046184 0 0.00046194 3.3 0.00046185999999999997 3.3 0.00046196 0 0.00046187999999999996 0 0.00046197999999999996 3.3 0.0004619 3.3 0.000462 0 0.00046192 0 0.00046202 3.3 0.00046194 3.3 0.00046204 0 0.00046196 0 0.00046206 3.3 0.00046197999999999996 3.3 0.00046207999999999997 0 0.000462 0 0.0004621 3.3 0.00046202 3.3 0.00046212 0 0.00046204 0 0.00046214 3.3 0.00046206 3.3 0.00046216 0 0.00046207999999999997 0 0.00046217999999999997 3.3 0.0004621 3.3 0.0004622 0 0.00046212 0 0.00046222 3.3 0.00046214 3.3 0.00046224 0 0.00046216 0 0.00046226 3.3 0.00046217999999999997 3.3 0.00046227999999999997 0 0.0004622 0 0.0004623 3.3 0.00046222 3.3 0.00046232 0 0.00046224 0 0.00046234 3.3 0.00046226 3.3 0.00046236 0 0.00046227999999999997 0 0.00046238 3.3 0.00046229999999999996 3.3 0.00046239999999999996 0 0.00046232 0 0.00046242 3.3 0.00046234 3.3 0.00046244 0 0.00046236 0 0.00046246 3.3 0.00046238 3.3 0.00046248 0 0.00046239999999999996 0 0.00046249999999999997 3.3 0.00046242 3.3 0.00046252 0 0.00046244 0 0.00046254 3.3 0.00046246 3.3 0.00046256 0 0.00046248 0 0.00046258 3.3 0.00046249999999999997 3.3 0.00046259999999999997 0 0.00046252 0 0.00046262 3.3 0.00046254 3.3 0.00046264 0 0.00046256 0 0.00046266 3.3 0.00046258 3.3 0.00046268 0 0.00046259999999999997 0 0.00046269999999999997 3.3 0.00046262 3.3 0.00046272 0 0.00046264 0 0.00046274 3.3 0.00046266 3.3 0.00046276 0 0.00046268 0 0.00046278 3.3 0.00046269999999999997 3.3 0.0004628 0 0.00046272 0 0.00046282 3.3 0.00046274 3.3 0.00046284 0 0.00046276 0 0.00046286 3.3 0.00046278 3.3 0.00046288 0 0.0004628 0 0.0004629 3.3 0.00046281999999999996 3.3 0.00046291999999999997 0 0.00046284 0 0.00046294 3.3 0.00046286 3.3 0.00046296 0 0.00046288 0 0.00046298 3.3 0.0004629 3.3 0.000463 0 0.00046291999999999997 0 0.00046301999999999997 3.3 0.00046294 3.3 0.00046304 0 0.00046296 0 0.00046306 3.3 0.00046298 3.3 0.00046308 0 0.000463 0 0.0004631 3.3 0.00046301999999999997 3.3 0.00046311999999999997 0 0.00046304 0 0.00046314 3.3 0.00046306 3.3 0.00046316 0 0.00046308 0 0.00046318 3.3 0.0004631 3.3 0.0004632 0 0.00046311999999999997 0 0.00046322 3.3 0.00046314 3.3 0.00046324 0 0.00046316 0 0.00046326 3.3 0.00046318 3.3 0.00046328 0 0.0004632 0 0.0004633 3.3 0.00046322 3.3 0.00046332 0 0.00046323999999999996 0 0.00046333999999999996 3.3 0.00046326 3.3 0.00046336 0 0.00046328 0 0.00046338 3.3 0.0004633 3.3 0.0004634 0 0.00046332 0 0.00046342 3.3 0.00046333999999999996 3.3 0.00046343999999999997 0 0.00046336 0 0.00046346 3.3 0.00046338 3.3 0.00046348 0 0.0004634 0 0.0004635 3.3 0.00046342 3.3 0.00046352 0 0.00046343999999999997 0 0.00046353999999999997 3.3 0.00046346 3.3 0.00046356 0 0.00046348 0 0.00046358 3.3 0.0004635 3.3 0.0004636 0 0.00046352 0 0.00046362 3.3 0.00046353999999999997 3.3 0.00046363999999999997 0 0.00046356 0 0.00046366 3.3 0.00046358 3.3 0.00046368 0 0.0004636 0 0.0004637 3.3 0.00046362 3.3 0.00046372 0 0.00046363999999999997 0 0.00046374 3.3 0.00046365999999999996 3.3 0.00046375999999999996 0 0.00046368 0 0.00046378 3.3 0.0004637 3.3 0.0004638 0 0.00046372 0 0.00046382 3.3 0.00046374 3.3 0.00046384 0 0.00046375999999999996 0 0.00046385999999999997 3.3 0.00046378 3.3 0.00046388 0 0.0004638 0 0.0004639 3.3 0.00046382 3.3 0.00046392 0 0.00046384 0 0.00046394 3.3 0.00046385999999999997 3.3 0.00046395999999999997 0 0.00046388 0 0.00046398 3.3 0.0004639 3.3 0.000464 0 0.00046392 0 0.00046402 3.3 0.00046394 3.3 0.00046404 0 0.00046395999999999997 0 0.00046405999999999997 3.3 0.00046398 3.3 0.00046408 0 0.000464 0 0.0004641 3.3 0.00046402 3.3 0.00046412 0 0.00046404 0 0.00046414 3.3 0.00046405999999999997 3.3 0.00046416 0 0.00046407999999999996 0 0.00046417999999999996 3.3 0.0004641 3.3 0.0004642 0 0.00046412 0 0.00046422 3.3 0.00046414 3.3 0.00046424 0 0.00046416 0 0.00046426 3.3 0.00046417999999999996 3.3 0.00046427999999999997 0 0.0004642 0 0.0004643 3.3 0.00046422 3.3 0.00046432 0 0.00046424 0 0.00046434 3.3 0.00046426 3.3 0.00046436 0 0.00046427999999999997 0 0.00046437999999999997 3.3 0.0004643 3.3 0.0004644 0 0.00046432 0 0.00046442 3.3 0.00046434 3.3 0.00046444 0 0.00046436 0 0.00046446 3.3 0.00046437999999999997 3.3 0.00046447999999999997 0 0.0004644 0 0.0004645 3.3 0.00046442 3.3 0.00046452 0 0.00046444 0 0.00046454 3.3 0.00046446 3.3 0.00046456 0 0.00046447999999999997 0 0.00046458 3.3 0.0004645 3.3 0.0004646 0 0.00046452 0 0.00046462 3.3 0.00046454 3.3 0.00046464 0 0.00046456 0 0.00046466 3.3 0.00046458 3.3 0.00046468 0 0.00046459999999999996 0 0.00046469999999999997 3.3 0.00046462 3.3 0.00046472 0 0.00046464 0 0.00046474 3.3 0.00046466 3.3 0.00046476 0 0.00046468 0 0.00046478 3.3 0.00046469999999999997 3.3 0.00046479999999999997 0 0.00046472 0 0.00046482 3.3 0.00046474 3.3 0.00046484 0 0.00046476 0 0.00046486 3.3 0.00046478 3.3 0.00046488 0 0.00046479999999999997 0 0.00046489999999999997 3.3 0.00046482 3.3 0.00046492 0 0.00046484 0 0.00046494 3.3 0.00046486 3.3 0.00046496 0 0.00046488 0 0.00046498 3.3 0.00046489999999999997 3.3 0.00046499999999999997 0 0.00046492 0 0.00046502 3.3 0.00046494 3.3 0.00046504 0 0.00046496 0 0.00046506 3.3 0.00046498 3.3 0.00046508 0 0.00046499999999999997 0 0.0004651 3.3 0.00046501999999999996 3.3 0.00046511999999999996 0 0.00046504 0 0.00046514 3.3 0.00046506 3.3 0.00046516 0 0.00046508 0 0.00046518 3.3 0.0004651 3.3 0.0004652 0 0.00046511999999999996 0 0.00046521999999999997 3.3 0.00046514 3.3 0.00046524 0 0.00046516 0 0.00046526 3.3 0.00046518 3.3 0.00046528 0 0.0004652 0 0.0004653 3.3 0.00046521999999999997 3.3 0.00046531999999999997 0 0.00046524 0 0.00046534 3.3 0.00046526 3.3 0.00046536 0 0.00046528 0 0.00046538 3.3 0.0004653 3.3 0.0004654 0 0.00046531999999999997 0 0.00046541999999999997 3.3 0.00046534 3.3 0.00046544 0 0.00046536 0 0.00046546 3.3 0.00046538 3.3 0.00046548 0 0.0004654 0 0.0004655 3.3 0.00046541999999999997 3.3 0.00046552 0 0.00046543999999999996 0 0.00046553999999999996 3.3 0.00046546 3.3 0.00046556 0 0.00046548 0 0.00046558 3.3 0.0004655 3.3 0.0004656 0 0.00046552 0 0.00046562 3.3 0.00046553999999999996 3.3 0.00046563999999999997 0 0.00046556 0 0.00046566 3.3 0.00046558 3.3 0.00046568 0 0.0004656 0 0.0004657 3.3 0.00046562 3.3 0.00046572 0 0.00046563999999999997 0 0.00046573999999999997 3.3 0.00046566 3.3 0.00046576 0 0.00046568 0 0.00046578 3.3 0.0004657 3.3 0.0004658 0 0.00046572 0 0.00046582 3.3 0.00046573999999999997 3.3 0.00046583999999999997 0 0.00046576 0 0.00046586 3.3 0.00046578 3.3 0.00046588 0 0.0004658 0 0.0004659 3.3 0.00046582 3.3 0.00046592 0 0.00046583999999999997 0 0.00046594 3.3 0.00046585999999999996 3.3 0.00046595999999999996 0 0.00046588 0 0.00046598 3.3 0.0004659 3.3 0.000466 0 0.00046592 0 0.00046602 3.3 0.00046594 3.3 0.00046604 0 0.00046595999999999996 0 0.00046605999999999997 3.3 0.00046598 3.3 0.00046608 0 0.000466 0 0.0004661 3.3 0.00046602 3.3 0.00046612 0 0.00046604 0 0.00046614 3.3 0.00046605999999999997 3.3 0.00046615999999999997 0 0.00046608 0 0.00046618 3.3 0.0004661 3.3 0.0004662 0 0.00046612 0 0.00046622 3.3 0.00046614 3.3 0.00046624 0 0.00046615999999999997 0 0.00046625999999999997 3.3 0.00046618 3.3 0.00046628 0 0.0004662 0 0.0004663 3.3 0.00046622 3.3 0.00046632 0 0.00046624 0 0.00046634 3.3 0.00046625999999999997 3.3 0.00046636 0 0.00046628 0 0.00046638 3.3 0.0004663 3.3 0.0004664 0 0.00046632 0 0.00046642 3.3 0.00046634 3.3 0.00046644 0 0.00046636 0 0.00046646 3.3 0.00046637999999999996 3.3 0.00046647999999999997 0 0.0004664 0 0.0004665 3.3 0.00046642 3.3 0.00046652 0 0.00046644 0 0.00046654 3.3 0.00046646 3.3 0.00046656 0 0.00046647999999999997 0 0.00046657999999999997 3.3 0.0004665 3.3 0.0004666 0 0.00046652 0 0.00046662 3.3 0.00046654 3.3 0.00046664 0 0.00046656 0 0.00046666 3.3 0.00046657999999999997 3.3 0.00046667999999999997 0 0.0004666 0 0.0004667 3.3 0.00046662 3.3 0.00046672 0 0.00046664 0 0.00046674 3.3 0.00046666 3.3 0.00046676 0 0.00046667999999999997 0 0.00046677999999999997 3.3 0.0004667 3.3 0.0004668 0 0.00046672 0 0.00046682 3.3 0.00046674 3.3 0.00046684 0 0.00046676 0 0.00046686 3.3 0.00046677999999999997 3.3 0.00046688 0 0.00046679999999999996 0 0.00046689999999999996 3.3 0.00046682 3.3 0.00046692 0 0.00046684 0 0.00046694 3.3 0.00046686 3.3 0.00046696 0 0.00046688 0 0.00046698 3.3 0.00046689999999999996 3.3 0.00046699999999999997 0 0.00046692 0 0.00046702 3.3 0.00046694 3.3 0.00046704 0 0.00046696 0 0.00046706 3.3 0.00046698 3.3 0.00046708 0 0.00046699999999999997 0 0.00046709999999999997 3.3 0.00046702 3.3 0.00046712 0 0.00046704 0 0.00046714 3.3 0.00046706 3.3 0.00046716 0 0.00046708 0 0.00046718 3.3 0.00046709999999999997 3.3 0.00046719999999999997 0 0.00046712 0 0.00046722 3.3 0.00046714 3.3 0.00046724 0 0.00046716 0 0.00046726 3.3 0.00046718 3.3 0.00046728 0 0.00046719999999999997 0 0.0004673 3.3 0.00046721999999999996 3.3 0.00046731999999999996 0 0.00046724 0 0.00046734 3.3 0.00046726 3.3 0.00046736 0 0.00046728 0 0.00046738 3.3 0.0004673 3.3 0.0004674 0 0.00046731999999999996 0 0.00046741999999999997 3.3 0.00046734 3.3 0.00046744 0 0.00046736 0 0.00046746 3.3 0.00046738 3.3 0.00046748 0 0.0004674 0 0.0004675 3.3 0.00046741999999999997 3.3 0.00046751999999999997 0 0.00046744 0 0.00046754 3.3 0.00046746 3.3 0.00046756 0 0.00046748 0 0.00046758 3.3 0.0004675 3.3 0.0004676 0 0.00046751999999999997 0 0.00046761999999999997 3.3 0.00046754 3.3 0.00046764 0 0.00046756 0 0.00046766 3.3 0.00046758 3.3 0.00046768 0 0.0004676 0 0.0004677 3.3 0.00046761999999999997 3.3 0.00046772 0 0.00046763999999999996 0 0.00046773999999999996 3.3 0.00046766 3.3 0.00046776 0 0.00046768 0 0.00046778 3.3 0.0004677 3.3 0.0004678 0 0.00046772 0 0.00046782 3.3 0.00046773999999999996 3.3 0.00046783999999999997 0 0.00046776 0 0.00046786 3.3 0.00046778 3.3 0.00046788 0 0.0004678 0 0.0004679 3.3 0.00046782 3.3 0.00046792 0 0.00046783999999999997 0 0.00046793999999999997 3.3 0.00046786 3.3 0.00046796 0 0.00046788 0 0.00046798 3.3 0.0004679 3.3 0.000468 0 0.00046792 0 0.00046802 3.3 0.00046793999999999997 3.3 0.00046803999999999997 0 0.00046796 0 0.00046806 3.3 0.00046798 3.3 0.00046808 0 0.000468 0 0.0004681 3.3 0.00046802 3.3 0.00046812 0 0.00046803999999999997 0 0.00046814 3.3 0.00046806 3.3 0.00046816 0 0.00046808 0 0.00046818 3.3 0.0004681 3.3 0.0004682 0 0.00046812 0 0.00046822 3.3 0.00046814 3.3 0.00046824 0 0.00046815999999999996 0 0.00046825999999999997 3.3 0.00046818 3.3 0.00046828 0 0.0004682 0 0.0004683 3.3 0.00046822 3.3 0.00046832 0 0.00046824 0 0.00046834 3.3 0.00046825999999999997 3.3 0.00046835999999999997 0 0.00046828 0 0.00046838 3.3 0.0004683 3.3 0.0004684 0 0.00046832 0 0.00046842 3.3 0.00046834 3.3 0.00046844 0 0.00046835999999999997 0 0.00046845999999999997 3.3 0.00046838 3.3 0.00046848 0 0.0004684 0 0.0004685 3.3 0.00046842 3.3 0.00046852 0 0.00046844 0 0.00046854 3.3 0.00046845999999999997 3.3 0.00046855999999999997 0 0.00046848 0 0.00046858 3.3 0.0004685 3.3 0.0004686 0 0.00046852 0 0.00046862 3.3 0.00046854 3.3 0.00046864 0 0.00046855999999999997 0 0.00046866 3.3 0.00046857999999999996 3.3 0.00046867999999999996 0 0.0004686 0 0.0004687 3.3 0.00046862 3.3 0.00046872 0 0.00046864 0 0.00046874 3.3 0.00046866 3.3 0.00046876 0 0.00046867999999999996 0 0.00046877999999999997 3.3 0.0004687 3.3 0.0004688 0 0.00046872 0 0.00046882 3.3 0.00046874 3.3 0.00046884 0 0.00046876 0 0.00046886 3.3 0.00046877999999999997 3.3 0.00046887999999999997 0 0.0004688 0 0.0004689 3.3 0.00046882 3.3 0.00046892 0 0.00046884 0 0.00046894 3.3 0.00046886 3.3 0.00046896 0 0.00046887999999999997 0 0.00046897999999999997 3.3 0.0004689 3.3 0.000469 0 0.00046892 0 0.00046902 3.3 0.00046894 3.3 0.00046904 0 0.00046896 0 0.00046906 3.3 0.00046897999999999997 3.3 0.00046908 0 0.00046899999999999996 0 0.00046909999999999996 3.3 0.00046902 3.3 0.00046912 0 0.00046904 0 0.00046914 3.3 0.00046906 3.3 0.00046916 0 0.00046908 0 0.00046918 3.3 0.00046909999999999996 3.3 0.00046919999999999997 0 0.00046912 0 0.00046922 3.3 0.00046914 3.3 0.00046924 0 0.00046916 0 0.00046926 3.3 0.00046918 3.3 0.00046928 0 0.00046919999999999997 0 0.00046929999999999997 3.3 0.00046922 3.3 0.00046932 0 0.00046924 0 0.00046934 3.3 0.00046926 3.3 0.00046936 0 0.00046928 0 0.00046938 3.3 0.00046929999999999997 3.3 0.00046939999999999997 0 0.00046932 0 0.00046942 3.3 0.00046934 3.3 0.00046944 0 0.00046936 0 0.00046946 3.3 0.00046938 3.3 0.00046948 0 0.00046939999999999997 0 0.0004695 3.3 0.00046942 3.3 0.00046952 0 0.00046944 0 0.00046954 3.3 0.00046946 3.3 0.00046956 0 0.00046948 0 0.00046958 3.3 0.0004695 3.3 0.0004696 0 0.00046951999999999996 0 0.00046961999999999997 3.3 0.00046954 3.3 0.00046964 0 0.00046956 0 0.00046966 3.3 0.00046958 3.3 0.00046968 0 0.0004696 0 0.0004697 3.3 0.00046961999999999997 3.3 0.00046971999999999997 0 0.00046964 0 0.00046974 3.3 0.00046966 3.3 0.00046976 0 0.00046968 0 0.00046978 3.3 0.0004697 3.3 0.0004698 0 0.00046971999999999997 0 0.00046981999999999997 3.3 0.00046974 3.3 0.00046984 0 0.00046976 0 0.00046986 3.3 0.00046978 3.3 0.00046988 0 0.0004698 0 0.0004699 3.3 0.00046981999999999997 3.3 0.00046992 0 0.00046984 0 0.00046994 3.3 0.00046986 3.3 0.00046996 0 0.00046988 0 0.00046998 3.3 0.0004699 3.3 0.00047 0 0.00046992 0 0.00047002 3.3 0.00046993999999999996 3.3 0.00047003999999999997 0 0.00046996 0 0.00047006 3.3 0.00046998 3.3 0.00047008 0 0.00047 0 0.0004701 3.3 0.00047002 3.3 0.00047012 0 0.00047003999999999997 0 0.00047013999999999997 3.3 0.00047006 3.3 0.00047016 0 0.00047008 0 0.00047018 3.3 0.0004701 3.3 0.0004702 0 0.00047012 0 0.00047022 3.3 0.00047013999999999997 3.3 0.00047023999999999997 0 0.00047016 0 0.00047026 3.3 0.00047018 3.3 0.00047028 0 0.0004702 0 0.0004703 3.3 0.00047022 3.3 0.00047032 0 0.00047023999999999997 0 0.00047033999999999997 3.3 0.00047026 3.3 0.00047036 0 0.00047028 0 0.00047038 3.3 0.0004703 3.3 0.0004704 0 0.00047032 0 0.00047042 3.3 0.00047033999999999997 3.3 0.00047044 0 0.00047035999999999996 0 0.00047045999999999996 3.3 0.00047038 3.3 0.00047048 0 0.0004704 0 0.0004705 3.3 0.00047042 3.3 0.00047052 0 0.00047044 0 0.00047054 3.3 0.00047045999999999996 3.3 0.00047055999999999997 0 0.00047048 0 0.00047058 3.3 0.0004705 3.3 0.0004706 0 0.00047052 0 0.00047062 3.3 0.00047054 3.3 0.00047064 0 0.00047055999999999997 0 0.00047065999999999997 3.3 0.00047058 3.3 0.00047068 0 0.0004706 0 0.0004707 3.3 0.00047062 3.3 0.00047072 0 0.00047064 0 0.00047074 3.3 0.00047065999999999997 3.3 0.00047075999999999997 0 0.00047068 0 0.00047078 3.3 0.0004707 3.3 0.0004708 0 0.00047072 0 0.00047082 3.3 0.00047074 3.3 0.00047084 0 0.00047075999999999997 0 0.00047086 3.3 0.00047077999999999996 3.3 0.00047087999999999996 0 0.0004708 0 0.0004709 3.3 0.00047082 3.3 0.00047092 0 0.00047084 0 0.00047094 3.3 0.00047086 3.3 0.00047096 0 0.00047087999999999996 0 0.00047097999999999997 3.3 0.0004709 3.3 0.000471 0 0.00047092 0 0.00047102 3.3 0.00047094 3.3 0.00047104 0 0.00047096 0 0.00047106 3.3 0.00047097999999999997 3.3 0.00047107999999999997 0 0.000471 0 0.0004711 3.3 0.00047102 3.3 0.00047112 0 0.00047104 0 0.00047114 3.3 0.00047106 3.3 0.00047116 0 0.00047107999999999997 0 0.00047117999999999997 3.3 0.0004711 3.3 0.0004712 0 0.00047112 0 0.00047122 3.3 0.00047114 3.3 0.00047124 0 0.00047116 0 0.00047126 3.3 0.00047117999999999997 3.3 0.00047128 0 0.0004712 0 0.0004713 3.3 0.00047122 3.3 0.00047132 0 0.00047124 0 0.00047134 3.3 0.00047126 3.3 0.00047136 0 0.00047128 0 0.00047138 3.3 0.00047129999999999996 3.3 0.00047139999999999997 0 0.00047132 0 0.00047142 3.3 0.00047134 3.3 0.00047144 0 0.00047136 0 0.00047146 3.3 0.00047138 3.3 0.00047148 0 0.00047139999999999997 0 0.00047149999999999997 3.3 0.00047142 3.3 0.00047152 0 0.00047144 0 0.00047154 3.3 0.00047146 3.3 0.00047156 0 0.00047148 0 0.00047158 3.3 0.00047149999999999997 3.3 0.00047159999999999997 0 0.00047152 0 0.00047162 3.3 0.00047154 3.3 0.00047164 0 0.00047156 0 0.00047166 3.3 0.00047158 3.3 0.00047168 0 0.00047159999999999997 0 0.0004717 3.3 0.00047162 3.3 0.00047172 0 0.00047164 0 0.00047174 3.3 0.00047166 3.3 0.00047176 0 0.00047168 0 0.00047178 3.3 0.0004717 3.3 0.0004718 0 0.00047171999999999996 0 0.00047181999999999997 3.3 0.00047174 3.3 0.00047184 0 0.00047176 0 0.00047186 3.3 0.00047178 3.3 0.00047188 0 0.0004718 0 0.0004719 3.3 0.00047181999999999997 3.3 0.00047191999999999997 0 0.00047184 0 0.00047194 3.3 0.00047186 3.3 0.00047196 0 0.00047188 0 0.00047198 3.3 0.0004719 3.3 0.000472 0 0.00047191999999999997 0 0.00047201999999999997 3.3 0.00047194 3.3 0.00047204 0 0.00047196 0 0.00047206 3.3 0.00047198 3.3 0.00047208 0 0.000472 0 0.0004721 3.3 0.00047201999999999997 3.3 0.00047211999999999997 0 0.00047204 0 0.00047214 3.3 0.00047206 3.3 0.00047216 0 0.00047208 0 0.00047218 3.3 0.0004721 3.3 0.0004722 0 0.00047211999999999997 0 0.00047222 3.3 0.00047213999999999996 3.3 0.00047223999999999996 0 0.00047216 0 0.00047226 3.3 0.00047218 3.3 0.00047228 0 0.0004722 0 0.0004723 3.3 0.00047222 3.3 0.00047232 0 0.00047223999999999996 0 0.00047233999999999997 3.3 0.00047226 3.3 0.00047236 0 0.00047228 0 0.00047238 3.3 0.0004723 3.3 0.0004724 0 0.00047232 0 0.00047242 3.3 0.00047233999999999997 3.3 0.00047243999999999997 0 0.00047236 0 0.00047246 3.3 0.00047238 3.3 0.00047248 0 0.0004724 0 0.0004725 3.3 0.00047242 3.3 0.00047252 0 0.00047243999999999997 0 0.00047253999999999997 3.3 0.00047246 3.3 0.00047256 0 0.00047248 0 0.00047258 3.3 0.0004725 3.3 0.0004726 0 0.00047252 0 0.00047262 3.3 0.00047253999999999997 3.3 0.00047264 0 0.00047255999999999996 0 0.00047265999999999996 3.3 0.00047258 3.3 0.00047268 0 0.0004726 0 0.0004727 3.3 0.00047262 3.3 0.00047272 0 0.00047264 0 0.00047274 3.3 0.00047265999999999996 3.3 0.00047275999999999997 0 0.00047268 0 0.00047278 3.3 0.0004727 3.3 0.0004728 0 0.00047272 0 0.00047282 3.3 0.00047274 3.3 0.00047284 0 0.00047275999999999997 0 0.00047285999999999997 3.3 0.00047278 3.3 0.00047288 0 0.0004728 0 0.0004729 3.3 0.00047282 3.3 0.00047292 0 0.00047284 0 0.00047294 3.3 0.00047285999999999997 3.3 0.00047295999999999997 0 0.00047288 0 0.00047298 3.3 0.0004729 3.3 0.000473 0 0.00047292 0 0.00047302 3.3 0.00047294 3.3 0.00047304 0 0.00047295999999999997 0 0.00047306 3.3 0.00047298 3.3 0.00047308 0 0.000473 0 0.0004731 3.3 0.00047302 3.3 0.00047312 0 0.00047304 0 0.00047314 3.3 0.00047306 3.3 0.00047316 0 0.00047307999999999996 0 0.00047317999999999997 3.3 0.0004731 3.3 0.0004732 0 0.00047312 0 0.00047322 3.3 0.00047314 3.3 0.00047324 0 0.00047316 0 0.00047326 3.3 0.00047317999999999997 3.3 0.00047327999999999997 0 0.0004732 0 0.0004733 3.3 0.00047322 3.3 0.00047332 0 0.00047324 0 0.00047334 3.3 0.00047326 3.3 0.00047336 0 0.00047327999999999997 0 0.00047337999999999997 3.3 0.0004733 3.3 0.0004734 0 0.00047332 0 0.00047342 3.3 0.00047334 3.3 0.00047344 0 0.00047336 0 0.00047346 3.3 0.00047337999999999997 3.3 0.00047348 0 0.0004734 0 0.0004735 3.3 0.00047342 3.3 0.00047352 0 0.00047344 0 0.00047354 3.3 0.00047346 3.3 0.00047356 0 0.00047348 0 0.00047358 3.3 0.00047349999999999996 3.3 0.00047359999999999997 0 0.00047352 0 0.00047362 3.3 0.00047354 3.3 0.00047364 0 0.00047356 0 0.00047366 3.3 0.00047358 3.3 0.00047368 0 0.00047359999999999997 0 0.00047369999999999997 3.3 0.00047362 3.3 0.00047372 0 0.00047364 0 0.00047374 3.3 0.00047366 3.3 0.00047376 0 0.00047368 0 0.00047378 3.3 0.00047369999999999997 3.3 0.00047379999999999997 0 0.00047372 0 0.00047382 3.3 0.00047374 3.3 0.00047384 0 0.00047376 0 0.00047386 3.3 0.00047378 3.3 0.00047388 0 0.00047379999999999997 0 0.00047389999999999997 3.3 0.00047382 3.3 0.00047392 0 0.00047384 0 0.00047394 3.3 0.00047386 3.3 0.00047396 0 0.00047388 0 0.00047398 3.3 0.00047389999999999997 3.3 0.000474 0 0.00047391999999999996 0 0.00047401999999999996 3.3 0.00047394 3.3 0.00047404 0 0.00047396 0 0.00047406 3.3 0.00047398 3.3 0.00047408 0 0.000474 0 0.0004741 3.3 0.00047401999999999996 3.3 0.00047411999999999997 0 0.00047404 0 0.00047414 3.3 0.00047406 3.3 0.00047416 0 0.00047408 0 0.00047418 3.3 0.0004741 3.3 0.0004742 0 0.00047411999999999997 0 0.00047421999999999997 3.3 0.00047414 3.3 0.00047424 0 0.00047416 0 0.00047426 3.3 0.00047418 3.3 0.00047428 0 0.0004742 0 0.0004743 3.3 0.00047421999999999997 3.3 0.00047431999999999997 0 0.00047424 0 0.00047434 3.3 0.00047426 3.3 0.00047436 0 0.00047428 0 0.00047438 3.3 0.0004743 3.3 0.0004744 0 0.00047431999999999997 0 0.00047442 3.3 0.00047433999999999996 3.3 0.00047443999999999996 0 0.00047436 0 0.00047446 3.3 0.00047438 3.3 0.00047448 0 0.0004744 0 0.0004745 3.3 0.00047442 3.3 0.00047452 0 0.00047443999999999996 0 0.00047453999999999997 3.3 0.00047446 3.3 0.00047456 0 0.00047448 0 0.00047458 3.3 0.0004745 3.3 0.0004746 0 0.00047452 0 0.00047462 3.3 0.00047453999999999997 3.3 0.00047463999999999997 0 0.00047456 0 0.00047466 3.3 0.00047458 3.3 0.00047468 0 0.0004746 0 0.0004747 3.3 0.00047462 3.3 0.00047472 0 0.00047463999999999997 0 0.00047473999999999997 3.3 0.00047466 3.3 0.00047476 0 0.00047468 0 0.00047478 3.3 0.0004747 3.3 0.0004748 0 0.00047472 0 0.00047482 3.3 0.00047473999999999997 3.3 0.00047484 0 0.00047476 0 0.00047486 3.3 0.00047478 3.3 0.00047488 0 0.0004748 0 0.0004749 3.3 0.00047482 3.3 0.00047492 0 0.00047484 0 0.00047494 3.3 0.00047485999999999996 3.3 0.00047495999999999997 0 0.00047488 0 0.00047498 3.3 0.0004749 3.3 0.000475 0 0.00047492 0 0.00047502 3.3 0.00047494 3.3 0.00047504 0 0.00047495999999999997 0 0.00047505999999999997 3.3 0.00047498 3.3 0.00047508 0 0.000475 0 0.0004751 3.3 0.00047502 3.3 0.00047512 0 0.00047504 0 0.00047514 3.3 0.00047505999999999997 3.3 0.00047515999999999997 0 0.00047508 0 0.00047518 3.3 0.0004751 3.3 0.0004752 0 0.00047512 0 0.00047522 3.3 0.00047514 3.3 0.00047524 0 0.00047515999999999997 0 0.00047525999999999997 3.3 0.00047518 3.3 0.00047528 0 0.0004752 0 0.0004753 3.3 0.00047522 3.3 0.00047532 0 0.00047524 0 0.00047534 3.3 0.00047525999999999997 3.3 0.00047536 0 0.00047527999999999996 0 0.00047537999999999996 3.3 0.0004753 3.3 0.0004754 0 0.00047532 0 0.00047542 3.3 0.00047534 3.3 0.00047544 0 0.00047536 0 0.00047546 3.3 0.00047537999999999996 3.3 0.00047547999999999997 0 0.0004754 0 0.0004755 3.3 0.00047542 3.3 0.00047552 0 0.00047544 0 0.00047554 3.3 0.00047546 3.3 0.00047556 0 0.00047547999999999997 0 0.00047557999999999997 3.3 0.0004755 3.3 0.0004756 0 0.00047552 0 0.00047562 3.3 0.00047554 3.3 0.00047564 0 0.00047556 0 0.00047566 3.3 0.00047557999999999997 3.3 0.00047567999999999997 0 0.0004756 0 0.0004757 3.3 0.00047562 3.3 0.00047572 0 0.00047564 0 0.00047574 3.3 0.00047566 3.3 0.00047576 0 0.00047567999999999997 0 0.00047578 3.3 0.00047569999999999996 3.3 0.00047579999999999996 0 0.00047572 0 0.00047582 3.3 0.00047574 3.3 0.00047584 0 0.00047576 0 0.00047586 3.3 0.00047578 3.3 0.00047588 0 0.00047579999999999996 0 0.00047589999999999997 3.3 0.00047582 3.3 0.00047592 0 0.00047584 0 0.00047594 3.3 0.00047586 3.3 0.00047596 0 0.00047588 0 0.00047598 3.3 0.00047589999999999997 3.3 0.00047599999999999997 0 0.00047592 0 0.00047602 3.3 0.00047594 3.3 0.00047604 0 0.00047596 0 0.00047606 3.3 0.00047598 3.3 0.00047608 0 0.00047599999999999997 0 0.00047609999999999997 3.3 0.00047602 3.3 0.00047612 0 0.00047604 0 0.00047614 3.3 0.00047606 3.3 0.00047616 0 0.00047608 0 0.00047618 3.3 0.00047609999999999997 3.3 0.0004762 0 0.00047611999999999996 0 0.00047621999999999996 3.3 0.00047614 3.3 0.00047624 0 0.00047616 0 0.00047626 3.3 0.00047618 3.3 0.00047628 0 0.0004762 0 0.0004763 3.3 0.00047621999999999996 3.3 0.00047631999999999997 0 0.00047624 0 0.00047634 3.3 0.00047626 3.3 0.00047636 0 0.00047628 0 0.00047638 3.3 0.0004763 3.3 0.0004764 0 0.00047631999999999997 0 0.00047641999999999997 3.3 0.00047634 3.3 0.00047644 0 0.00047636 0 0.00047646 3.3 0.00047638 3.3 0.00047648 0 0.0004764 0 0.0004765 3.3 0.00047641999999999997 3.3 0.00047651999999999997 0 0.00047644 0 0.00047654 3.3 0.00047646 3.3 0.00047656 0 0.00047648 0 0.00047658 3.3 0.0004765 3.3 0.0004766 0 0.00047651999999999997 0 0.00047662 3.3 0.00047654 3.3 0.00047664 0 0.00047656 0 0.00047666 3.3 0.00047658 3.3 0.00047668 0 0.0004766 0 0.0004767 3.3 0.00047662 3.3 0.00047672 0 0.00047663999999999996 0 0.00047673999999999997 3.3 0.00047666 3.3 0.00047676 0 0.00047668 0 0.00047678 3.3 0.0004767 3.3 0.0004768 0 0.00047672 0 0.00047682 3.3 0.00047673999999999997 3.3 0.00047683999999999997 0 0.00047676 0 0.00047686 3.3 0.00047678 3.3 0.00047688 0 0.0004768 0 0.0004769 3.3 0.00047682 3.3 0.00047692 0 0.00047683999999999997 0 0.00047693999999999997 3.3 0.00047686 3.3 0.00047696 0 0.00047688 0 0.00047698 3.3 0.0004769 3.3 0.000477 0 0.00047692 0 0.00047702 3.3 0.00047693999999999997 3.3 0.00047703999999999997 0 0.00047696 0 0.00047706 3.3 0.00047698 3.3 0.00047708 0 0.000477 0 0.0004771 3.3 0.00047702 3.3 0.00047712 0 0.00047703999999999997 0 0.00047714 3.3 0.00047705999999999996 3.3 0.00047715999999999996 0 0.00047708 0 0.00047718 3.3 0.0004771 3.3 0.0004772 0 0.00047712 0 0.00047722 3.3 0.00047714 3.3 0.00047724 0 0.00047715999999999996 0 0.00047725999999999997 3.3 0.00047718 3.3 0.00047728 0 0.0004772 0 0.0004773 3.3 0.00047722 3.3 0.00047732 0 0.00047724 0 0.00047734 3.3 0.00047725999999999997 3.3 0.00047735999999999997 0 0.00047728 0 0.00047738 3.3 0.0004773 3.3 0.0004774 0 0.00047732 0 0.00047742 3.3 0.00047734 3.3 0.00047744 0 0.00047735999999999997 0 0.00047745999999999997 3.3 0.00047738 3.3 0.00047748 0 0.0004774 0 0.0004775 3.3 0.00047742 3.3 0.00047752 0 0.00047744 0 0.00047754 3.3 0.00047745999999999997 3.3 0.00047756 0 0.00047747999999999996 0 0.00047757999999999996 3.3 0.0004775 3.3 0.0004776 0 0.00047752 0 0.00047762 3.3 0.00047754 3.3 0.00047764 0 0.00047756 0 0.00047766 3.3 0.00047757999999999996 3.3 0.00047767999999999997 0 0.0004776 0 0.0004777 3.3 0.00047762 3.3 0.00047772 0 0.00047764 0 0.00047774 3.3 0.00047766 3.3 0.00047776 0 0.00047767999999999997 0 0.00047777999999999997 3.3 0.0004777 3.3 0.0004778 0 0.00047772 0 0.00047782 3.3 0.00047774 3.3 0.00047784 0 0.00047776 0 0.00047786 3.3 0.00047777999999999997 3.3 0.00047787999999999997 0 0.0004778 0 0.0004779 3.3 0.00047782 3.3 0.00047792 0 0.00047784 0 0.00047794 3.3 0.00047786 3.3 0.00047796 0 0.00047787999999999997 0 0.00047798 3.3 0.00047789999999999996 3.3 0.00047799999999999996 0 0.00047792 0 0.00047802 3.3 0.00047794 3.3 0.00047804 0 0.00047796 0 0.00047806 3.3 0.00047798 3.3 0.00047808 0 0.00047799999999999996 0 0.00047809999999999997 3.3 0.00047802 3.3 0.00047812 0 0.00047804 0 0.00047814 3.3 0.00047806 3.3 0.00047816 0 0.00047808 0 0.00047818 3.3 0.00047809999999999997 3.3 0.00047819999999999997 0 0.00047812 0 0.00047822 3.3 0.00047814 3.3 0.00047824 0 0.00047816 0 0.00047826 3.3 0.00047818 3.3 0.00047828 0 0.00047819999999999997 0 0.00047829999999999997 3.3 0.00047822 3.3 0.00047832 0 0.00047824 0 0.00047834 3.3 0.00047826 3.3 0.00047836 0 0.00047828 0 0.00047838 3.3 0.00047829999999999997 3.3 0.0004784 0 0.00047832 0 0.00047842 3.3 0.00047834 3.3 0.00047844 0 0.00047836 0 0.00047846 3.3 0.00047838 3.3 0.00047848 0 0.0004784 0 0.0004785 3.3 0.00047841999999999996 3.3 0.00047851999999999997 0 0.00047844 0 0.00047854 3.3 0.00047846 3.3 0.00047856 0 0.00047848 0 0.00047858 3.3 0.0004785 3.3 0.0004786 0 0.00047851999999999997 0 0.00047861999999999997 3.3 0.00047854 3.3 0.00047864 0 0.00047856 0 0.00047866 3.3 0.00047858 3.3 0.00047868 0 0.0004786 0 0.0004787 3.3 0.00047861999999999997 3.3 0.00047871999999999997 0 0.00047864 0 0.00047874 3.3 0.00047866 3.3 0.00047876 0 0.00047868 0 0.00047878 3.3 0.0004787 3.3 0.0004788 0 0.00047871999999999997 0 0.00047881999999999997 3.3 0.00047874 3.3 0.00047884 0 0.00047876 0 0.00047886 3.3 0.00047878 3.3 0.00047888 0 0.0004788 0 0.0004789 3.3 0.00047881999999999997 3.3 0.00047892 0 0.00047883999999999996 0 0.00047893999999999996 3.3 0.00047886 3.3 0.00047896 0 0.00047888 0 0.00047898 3.3 0.0004789 3.3 0.000479 0 0.00047892 0 0.00047902 3.3 0.00047893999999999996 3.3 0.00047903999999999997 0 0.00047896 0 0.00047906 3.3 0.00047898 3.3 0.00047908 0 0.000479 0 0.0004791 3.3 0.00047902 3.3 0.00047912 0 0.00047903999999999997 0 0.00047913999999999997 3.3 0.00047906 3.3 0.00047916 0 0.00047908 0 0.00047918 3.3 0.0004791 3.3 0.0004792 0 0.00047912 0 0.00047922 3.3 0.00047913999999999997 3.3 0.00047923999999999997 0 0.00047916 0 0.00047926 3.3 0.00047918 3.3 0.00047928 0 0.0004792 0 0.0004793 3.3 0.00047922 3.3 0.00047932 0 0.00047923999999999997 0 0.00047934 3.3 0.00047925999999999996 3.3 0.00047935999999999996 0 0.00047928 0 0.00047938 3.3 0.0004793 3.3 0.0004794 0 0.00047932 0 0.00047942 3.3 0.00047934 3.3 0.00047944 0 0.00047935999999999996 0 0.00047945999999999997 3.3 0.00047938 3.3 0.00047948 0 0.0004794 0 0.0004795 3.3 0.00047942 3.3 0.00047952 0 0.00047944 0 0.00047954 3.3 0.00047945999999999997 3.3 0.00047955999999999997 0 0.00047948 0 0.00047958 3.3 0.0004795 3.3 0.0004796 0 0.00047952 0 0.00047962 3.3 0.00047954 3.3 0.00047964 0 0.00047955999999999997 0 0.00047965999999999997 3.3 0.00047958 3.3 0.00047968 0 0.0004796 0 0.0004797 3.3 0.00047962 3.3 0.00047972 0 0.00047964 0 0.00047974 3.3 0.00047965999999999997 3.3 0.00047976 0 0.00047967999999999996 0 0.00047977999999999996 3.3 0.0004797 3.3 0.0004798 0 0.00047972 0 0.00047982 3.3 0.00047974 3.3 0.00047984 0 0.00047976 0 0.00047986 3.3 0.00047977999999999996 3.3 0.00047987999999999997 0 0.0004798 0 0.0004799 3.3 0.00047982 3.3 0.00047992 0 0.00047984 0 0.00047994 3.3 0.00047986 3.3 0.00047996 0 0.00047987999999999997 0 0.00047997999999999997 3.3 0.0004799 3.3 0.00048 0 0.00047992 0 0.00048002 3.3 0.00047994 3.3 0.00048004 0 0.00047996 0 0.00048006 3.3 0.00047997999999999997 3.3 0.00048007999999999997 0 0.00048 0 0.0004801 3.3 0.00048002 3.3 0.00048012 0 0.00048004 0 0.00048014 3.3 0.00048006 3.3 0.00048016 0 0.00048007999999999997 0 0.00048018 3.3 0.0004801 3.3 0.0004802 0 0.00048012 0 0.00048022 3.3 0.00048014 3.3 0.00048024 0 0.00048016 0 0.00048026 3.3 0.00048018 3.3 0.00048028 0 0.00048019999999999996 0 0.00048029999999999997 3.3 0.00048022 3.3 0.00048032 0 0.00048024 0 0.00048034 3.3 0.00048026 3.3 0.00048036 0 0.00048028 0 0.00048038 3.3 0.00048029999999999997 3.3 0.00048039999999999997 0 0.00048032 0 0.00048042 3.3 0.00048034 3.3 0.00048044 0 0.00048036 0 0.00048046 3.3 0.00048038 3.3 0.00048048 0 0.00048039999999999997 0 0.00048049999999999997 3.3 0.00048042 3.3 0.00048052 0 0.00048044 0 0.00048054 3.3 0.00048046 3.3 0.00048056 0 0.00048048 0 0.00048058 3.3 0.00048049999999999997 3.3 0.00048059999999999997 0 0.00048052 0 0.00048062 3.3 0.00048054 3.3 0.00048064 0 0.00048056 0 0.00048066 3.3 0.00048058 3.3 0.00048068 0 0.00048059999999999997 0 0.0004807 3.3 0.00048061999999999996 3.3 0.00048071999999999996 0 0.00048064 0 0.00048074 3.3 0.00048066 3.3 0.00048076 0 0.00048068 0 0.00048078 3.3 0.0004807 3.3 0.0004808 0 0.00048071999999999996 0 0.00048081999999999997 3.3 0.00048074 3.3 0.00048084 0 0.00048076 0 0.00048086 3.3 0.00048078 3.3 0.00048088 0 0.0004808 0 0.0004809 3.3 0.00048081999999999997 3.3 0.00048091999999999997 0 0.00048084 0 0.00048094 3.3 0.00048086 3.3 0.00048096 0 0.00048088 0 0.00048098 3.3 0.0004809 3.3 0.000481 0 0.00048091999999999997 0 0.00048101999999999997 3.3 0.00048094 3.3 0.00048104 0 0.00048096 0 0.00048106 3.3 0.00048098 3.3 0.00048108 0 0.000481 0 0.0004811 3.3 0.00048101999999999997 3.3 0.00048112 0 0.00048103999999999996 0 0.00048113999999999996 3.3 0.00048106 3.3 0.00048116 0 0.00048108 0 0.00048118 3.3 0.0004811 3.3 0.0004812 0 0.00048112 0 0.00048122 3.3 0.00048113999999999996 3.3 0.00048123999999999997 0 0.00048116 0 0.00048126 3.3 0.00048118 3.3 0.00048128 0 0.0004812 0 0.0004813 3.3 0.00048122 3.3 0.00048132 0 0.00048123999999999997 0 0.00048133999999999997 3.3 0.00048126 3.3 0.00048136 0 0.00048128 0 0.00048138 3.3 0.0004813 3.3 0.0004814 0 0.00048132 0 0.00048142 3.3 0.00048133999999999997 3.3 0.00048143999999999997 0 0.00048136 0 0.00048146 3.3 0.00048138 3.3 0.00048148 0 0.0004814 0 0.0004815 3.3 0.00048142 3.3 0.00048152 0 0.00048143999999999997 0 0.00048154 3.3 0.00048145999999999996 3.3 0.00048155999999999996 0 0.00048148 0 0.00048158 3.3 0.0004815 3.3 0.0004816 0 0.00048152 0 0.00048162 3.3 0.00048154 3.3 0.00048164 0 0.00048155999999999996 0 0.00048165999999999997 3.3 0.00048158 3.3 0.00048168 0 0.0004816 0 0.0004817 3.3 0.00048162 3.3 0.00048172 0 0.00048164 0 0.00048174 3.3 0.00048165999999999997 3.3 0.00048175999999999997 0 0.00048168 0 0.00048178 3.3 0.0004817 3.3 0.0004818 0 0.00048172 0 0.00048182 3.3 0.00048174 3.3 0.00048184 0 0.00048175999999999997 0 0.00048185999999999997 3.3 0.00048178 3.3 0.00048188 0 0.0004818 0 0.0004819 3.3 0.00048182 3.3 0.00048192 0 0.00048184 0 0.00048194 3.3 0.00048185999999999997 3.3 0.00048196 0 0.00048188 0 0.00048198 3.3 0.0004819 3.3 0.000482 0 0.00048192 0 0.00048202 3.3 0.00048194 3.3 0.00048204 0 0.00048196 0 0.00048206 3.3 0.00048197999999999996 3.3 0.00048207999999999997 0 0.000482 0 0.0004821 3.3 0.00048202 3.3 0.00048212 0 0.00048204 0 0.00048214 3.3 0.00048206 3.3 0.00048216 0 0.00048207999999999997 0 0.00048217999999999997 3.3 0.0004821 3.3 0.0004822 0 0.00048212 0 0.00048222 3.3 0.00048214 3.3 0.00048224 0 0.00048216 0 0.00048226 3.3 0.00048217999999999997 3.3 0.00048227999999999997 0 0.0004822 0 0.0004823 3.3 0.00048222 3.3 0.00048232 0 0.00048224 0 0.00048234 3.3 0.00048226 3.3 0.00048236 0 0.00048227999999999997 0 0.00048237999999999997 3.3 0.0004823 3.3 0.0004824 0 0.00048232 0 0.00048242 3.3 0.00048234 3.3 0.00048244 0 0.00048236 0 0.00048246 3.3 0.00048237999999999997 3.3 0.00048248 0 0.00048239999999999996 0 0.00048249999999999996 3.3 0.00048242 3.3 0.00048252 0 0.00048244 0 0.00048254 3.3 0.00048246 3.3 0.00048256 0 0.00048248 0 0.00048258 3.3 0.00048249999999999996 3.3 0.00048259999999999997 0 0.00048252 0 0.00048262 3.3 0.00048254 3.3 0.00048264 0 0.00048256 0 0.00048266 3.3 0.00048258 3.3 0.00048268 0 0.00048259999999999997 0 0.00048269999999999997 3.3 0.00048262 3.3 0.00048272 0 0.00048264 0 0.00048274 3.3 0.00048266 3.3 0.00048276 0 0.00048268 0 0.00048278 3.3 0.00048269999999999997 3.3 0.00048279999999999997 0 0.00048272 0 0.00048282 3.3 0.00048274 3.3 0.00048284 0 0.00048276 0 0.00048286 3.3 0.00048278 3.3 0.00048288 0 0.00048279999999999997 0 0.0004829 3.3 0.00048281999999999996 3.3 0.00048291999999999996 0 0.00048284 0 0.00048294 3.3 0.00048286 3.3 0.00048296 0 0.00048288 0 0.00048298 3.3 0.0004829 3.3 0.000483 0 0.00048291999999999996 0 0.00048301999999999997 3.3 0.00048294 3.3 0.00048304 0 0.00048296 0 0.00048306 3.3 0.00048298 3.3 0.00048308 0 0.000483 0 0.0004831 3.3 0.00048301999999999997 3.3 0.00048311999999999997 0 0.00048304 0 0.00048314 3.3 0.00048306 3.3 0.00048316 0 0.00048308 0 0.00048318 3.3 0.0004831 3.3 0.0004832 0 0.00048311999999999997 0 0.00048321999999999997 3.3 0.00048314 3.3 0.00048324 0 0.00048316 0 0.00048326 3.3 0.00048318 3.3 0.00048328 0 0.0004832 0 0.0004833 3.3 0.00048321999999999997 3.3 0.00048332 0 0.00048323999999999996 0 0.00048333999999999996 3.3 0.00048326 3.3 0.00048336 0 0.00048328 0 0.00048338 3.3 0.0004833 3.3 0.0004834 0 0.00048332 0 0.00048342 3.3 0.00048333999999999996 3.3 0.00048343999999999997 0 0.00048336 0 0.00048346 3.3 0.00048338 3.3 0.00048348 0 0.0004834 0 0.0004835 3.3 0.00048342 3.3 0.00048352 0 0.00048343999999999997 0 0.00048353999999999997 3.3 0.00048346 3.3 0.00048356 0 0.00048348 0 0.00048358 3.3 0.0004835 3.3 0.0004836 0 0.00048352 0 0.00048362 3.3 0.00048353999999999997 3.3 0.00048363999999999997 0 0.00048356 0 0.00048366 3.3 0.00048358 3.3 0.00048368 0 0.0004836 0 0.0004837 3.3 0.00048362 3.3 0.00048372 0 0.00048363999999999997 0 0.00048374 3.3 0.00048366 3.3 0.00048376 0 0.00048368 0 0.00048378 3.3 0.0004837 3.3 0.0004838 0 0.00048372 0 0.00048382 3.3 0.00048374 3.3 0.00048384 0 0.00048375999999999996 0 0.00048385999999999997 3.3 0.00048378 3.3 0.00048388 0 0.0004838 0 0.0004839 3.3 0.00048382 3.3 0.00048392 0 0.00048384 0 0.00048394 3.3 0.00048385999999999997 3.3 0.00048395999999999997 0 0.00048388 0 0.00048398 3.3 0.0004839 3.3 0.000484 0 0.00048392 0 0.00048402 3.3 0.00048394 3.3 0.00048404 0 0.00048395999999999997 0 0.00048405999999999997 3.3 0.00048398 3.3 0.00048408 0 0.000484 0 0.0004841 3.3 0.00048402 3.3 0.00048412 0 0.00048404 0 0.00048414 3.3 0.00048405999999999997 3.3 0.00048415999999999997 0 0.00048408 0 0.00048418 3.3 0.0004841 3.3 0.0004842 0 0.00048412 0 0.00048422 3.3 0.00048414 3.3 0.00048424 0 0.00048415999999999997 0 0.00048426 3.3 0.00048417999999999996 3.3 0.00048427999999999996 0 0.0004842 0 0.0004843 3.3 0.00048422 3.3 0.00048432 0 0.00048424 0 0.00048434 3.3 0.00048426 3.3 0.00048436 0 0.00048427999999999996 0 0.00048437999999999997 3.3 0.0004843 3.3 0.0004844 0 0.00048432 0 0.00048442 3.3 0.00048434 3.3 0.00048444 0 0.00048436 0 0.00048446 3.3 0.00048437999999999997 3.3 0.00048447999999999997 0 0.0004844 0 0.0004845 3.3 0.00048442 3.3 0.00048452 0 0.00048444 0 0.00048454 3.3 0.00048446 3.3 0.00048456 0 0.00048447999999999997 0 0.00048457999999999997 3.3 0.0004845 3.3 0.0004846 0 0.00048452 0 0.00048462 3.3 0.00048454 3.3 0.00048464 0 0.00048456 0 0.00048466 3.3 0.00048457999999999997 3.3 0.00048468 0 0.00048459999999999996 0 0.00048469999999999996 3.3 0.00048462 3.3 0.00048472 0 0.00048464 0 0.00048474 3.3 0.00048466 3.3 0.00048476 0 0.00048468 0 0.00048478 3.3 0.00048469999999999996 3.3 0.00048479999999999997 0 0.00048472 0 0.00048482 3.3 0.00048474 3.3 0.00048484 0 0.00048476 0 0.00048486 3.3 0.00048478 3.3 0.00048488 0 0.00048479999999999997 0 0.00048489999999999997 3.3 0.00048482 3.3 0.00048492 0 0.00048484 0 0.00048494 3.3 0.00048486 3.3 0.00048496 0 0.00048488 0 0.00048498 3.3 0.00048489999999999997 3.3 0.00048499999999999997 0 0.00048492 0 0.00048502 3.3 0.00048494 3.3 0.00048504 0 0.00048496 0 0.00048506 3.3 0.00048498 3.3 0.00048508 0 0.00048499999999999997 0 0.0004851 3.3 0.00048501999999999996 3.3 0.00048511999999999996 0 0.00048504 0 0.00048514 3.3 0.00048506 3.3 0.00048516 0 0.00048508 0 0.00048518 3.3 0.0004851 3.3 0.0004852 0 0.00048511999999999996 0 0.00048521999999999997 3.3 0.00048514 3.3 0.00048524 0 0.00048516 0 0.00048526 3.3 0.00048518 3.3 0.00048528 0 0.0004852 0 0.0004853 3.3 0.00048521999999999997 3.3 0.00048531999999999997 0 0.00048524 0 0.00048534 3.3 0.00048526 3.3 0.00048536 0 0.00048528 0 0.00048538 3.3 0.0004853 3.3 0.0004854 0 0.00048531999999999997 0 0.00048541999999999997 3.3 0.00048534 3.3 0.00048544 0 0.00048536 0 0.00048546 3.3 0.00048538 3.3 0.00048548 0 0.0004854 0 0.0004855 3.3 0.00048541999999999997 3.3 0.00048551999999999997 0 0.00048544 0 0.00048554 3.3 0.00048546 3.3 0.00048556 0 0.00048548 0 0.00048558 3.3 0.0004855 3.3 0.0004856 0 0.00048551999999999997 0 0.00048562 3.3 0.00048553999999999996 3.3 0.00048563999999999996 0 0.00048556 0 0.00048566 3.3 0.00048558 3.3 0.00048568 0 0.0004856 0 0.0004857 3.3 0.00048562 3.3 0.00048572 0 0.00048563999999999996 0 0.00048573999999999997 3.3 0.00048566 3.3 0.00048576 0 0.00048568 0 0.00048578 3.3 0.0004857 3.3 0.0004858 0 0.00048572 0 0.00048582 3.3 0.00048573999999999997 3.3 0.00048583999999999997 0 0.00048576 0 0.00048586 3.3 0.00048578 3.3 0.00048588 0 0.0004858 0 0.0004859 3.3 0.00048582 3.3 0.00048592 0 0.00048583999999999997 0 0.00048593999999999997 3.3 0.00048586 3.3 0.00048596 0 0.00048588 0 0.00048598 3.3 0.0004859 3.3 0.000486 0 0.00048592 0 0.00048602 3.3 0.00048593999999999997 3.3 0.00048604 0 0.00048595999999999996 0 0.00048605999999999996 3.3 0.00048598 3.3 0.00048608 0 0.000486 0 0.0004861 3.3 0.00048602 3.3 0.00048612 0 0.00048604 0 0.00048614 3.3 0.00048605999999999996 3.3 0.00048615999999999997 0 0.00048608 0 0.00048618 3.3 0.0004861 3.3 0.0004862 0 0.00048612 0 0.00048622 3.3 0.00048614 3.3 0.00048624 0 0.00048615999999999997 0 0.00048625999999999997 3.3 0.00048618 3.3 0.00048628 0 0.0004862 0 0.0004863 3.3 0.00048622 3.3 0.00048632 0 0.00048624 0 0.00048634 3.3 0.00048625999999999997 3.3 0.00048635999999999997 0 0.00048628 0 0.00048638 3.3 0.0004863 3.3 0.0004864 0 0.00048632 0 0.00048642 3.3 0.00048634 3.3 0.00048644 0 0.00048635999999999997 0 0.00048646 3.3 0.00048637999999999996 3.3 0.00048647999999999996 0 0.0004864 0 0.0004865 3.3 0.00048642 3.3 0.00048652 0 0.00048644 0 0.00048654 3.3 0.00048646 3.3 0.00048656 0 0.00048647999999999996 0 0.00048657999999999997 3.3 0.0004865 3.3 0.0004866 0 0.00048652 0 0.00048662 3.3 0.00048654 3.3 0.00048664 0 0.00048656 0 0.00048666 3.3 0.00048657999999999997 3.3 0.00048667999999999997 0 0.0004866 0 0.0004867 3.3 0.00048662 3.3 0.00048672 0 0.00048664 0 0.00048674 3.3 0.00048666 3.3 0.00048676 0 0.00048667999999999997 0 0.00048677999999999997 3.3 0.0004867 3.3 0.0004868 0 0.00048672 0 0.00048682 3.3 0.00048674 3.3 0.00048684 0 0.00048676 0 0.00048686 3.3 0.00048677999999999997 3.3 0.00048688 0 0.0004868 0 0.0004869 3.3 0.00048682 3.3 0.00048692 0 0.00048684 0 0.00048694 3.3 0.00048686 3.3 0.00048696 0 0.00048688 0 0.00048698 3.3 0.00048689999999999996 3.3 0.00048699999999999997 0 0.00048692 0 0.00048702 3.3 0.00048694 3.3 0.00048704 0 0.00048696 0 0.00048706 3.3 0.00048698 3.3 0.00048708 0 0.00048699999999999997 0 0.00048709999999999997 3.3 0.00048702 3.3 0.00048712 0 0.00048704 0 0.00048714 3.3 0.00048706 3.3 0.00048716 0 0.00048708 0 0.00048718 3.3 0.00048709999999999997 3.3 0.00048719999999999997 0 0.00048712 0 0.00048722 3.3 0.00048714 3.3 0.00048724 0 0.00048716 0 0.00048726 3.3 0.00048718 3.3 0.00048728 0 0.00048719999999999997 0 0.00048729999999999997 3.3 0.00048722 3.3 0.00048732 0 0.00048724 0 0.00048734 3.3 0.00048726 3.3 0.00048736 0 0.00048728 0 0.00048738 3.3 0.00048729999999999997 3.3 0.0004874 0 0.00048731999999999996 0 0.00048741999999999996 3.3 0.00048734 3.3 0.00048744 0 0.00048736 0 0.00048746 3.3 0.00048738 3.3 0.00048748 0 0.0004874 0 0.0004875 3.3 0.00048741999999999996 3.3 0.00048751999999999997 0 0.00048744 0 0.00048754 3.3 0.00048746 3.3 0.00048756 0 0.00048748 0 0.00048758 3.3 0.0004875 3.3 0.0004876 0 0.00048751999999999997 0 0.00048761999999999997 3.3 0.00048754 3.3 0.00048764 0 0.00048756 0 0.00048766 3.3 0.00048758 3.3 0.00048768 0 0.0004876 0 0.0004877 3.3 0.00048761999999999997 3.3 0.00048771999999999997 0 0.00048764 0 0.00048774 3.3 0.00048766 3.3 0.00048776 0 0.00048768 0 0.00048778 3.3 0.0004877 3.3 0.0004878 0 0.00048771999999999997 0 0.00048782 3.3 0.00048773999999999996 3.3 0.00048783999999999996 0 0.00048776 0 0.00048786 3.3 0.00048778 3.3 0.00048788 0 0.0004878 0 0.0004879 3.3 0.00048782 3.3 0.00048792 0 0.00048783999999999996 0 0.00048793999999999997 3.3 0.00048786 3.3 0.00048796 0 0.00048788 0 0.00048798 3.3 0.0004879 3.3 0.000488 0 0.00048792 0 0.00048802 3.3 0.00048793999999999997 3.3 0.00048803999999999997 0 0.00048796 0 0.00048806 3.3 0.00048798 3.3 0.00048808 0 0.000488 0 0.0004881 3.3 0.00048802 3.3 0.00048812 0 0.00048803999999999997 0 0.00048813999999999997 3.3 0.00048806 3.3 0.00048816 0 0.00048808 0 0.00048818 3.3 0.0004881 3.3 0.0004882 0 0.00048812 0 0.00048822 3.3 0.00048813999999999997 3.3 0.00048824 0 0.00048815999999999996 0 0.00048825999999999996 3.3 0.00048818 3.3 0.00048828 0 0.0004882 0 0.0004883 3.3 0.00048822 3.3 0.00048832 0 0.00048824 0 0.00048834 3.3 0.00048825999999999996 3.3 0.00048836 0 0.00048827999999999995 0 0.00048838 3.3 0.0004883 3.3 0.0004883999999999999 0 0.0004883200000000001 0 0.00048842 3.3 0.0004883400000000001 3.3 0.00048844 0 0.0004883600000000001 0 0.00048846 3.3 0.0004883800000000001 3.3 0.00048848 0 0.0004884 0 0.0004885 3.3 0.00048842 3.3 0.00048852 0 0.00048844 0 0.00048854 3.3 0.00048846 3.3 0.00048856 0 0.00048848 0 0.00048858 3.3 0.0004885 3.3 0.0004886 0 0.00048852 0 0.0004886199999999999 3.3 0.0004885400000000001 3.3 0.00048864 0 0.0004885600000000001 0 0.00048866 3.3 0.0004885800000000001 3.3 0.00048868 0 0.0004886000000000001 0 0.0004887 3.3 0.00048862 3.3 0.00048872 0 0.00048864 0 0.00048874 3.3 0.00048866 3.3 0.00048876 0 0.00048868 0 0.00048878 3.3 0.0004887 3.3 0.0004888 0 0.00048872 0 0.0004888199999999999 3.3 0.0004887400000000001 3.3 0.00048884 0 0.0004887600000000001 0 0.00048886 3.3 0.0004887800000000001 3.3 0.00048888 0 0.0004888000000000001 0 0.0004889 3.3 0.00048882 3.3 0.00048892 0 0.00048884 0 0.00048894 3.3 0.00048886 3.3 0.00048896 0 0.00048888 0 0.00048898 3.3 0.0004889 3.3 0.000489 0 0.00048892 0 0.00048902 3.3 0.00048894 3.3 0.0004890399999999999 0 0.0004889600000000001 0 0.00048906 3.3 0.0004889800000000001 3.3 0.00048908 0 0.0004890000000000001 0 0.0004891 3.3 0.0004890200000000001 3.3 0.00048912 0 0.00048904 0 0.00048914 3.3 0.00048906 3.3 0.00048916 0 0.00048908 0 0.00048918 3.3 0.0004891 3.3 0.0004892 0 0.00048912 0 0.00048922 3.3 0.00048914 3.3 0.0004892399999999999 0 0.0004891600000000001 0 0.00048926 3.3 0.0004891800000000001 3.3 0.00048928 0 0.0004892000000000001 0 0.0004893 3.3 0.0004892200000000001 3.3 0.00048932 0 0.00048924 0 0.00048934 3.3 0.00048926 3.3 0.00048936 0 0.00048928 0 0.00048938 3.3 0.0004893 3.3 0.0004894 0 0.00048932 0 0.00048942 3.3 0.00048934 3.3 0.00048944 0 0.00048936 0 0.0004894599999999999 3.3 0.0004893800000000001 3.3 0.00048948 0 0.0004894000000000001 0 0.0004895 3.3 0.0004894200000000001 3.3 0.00048952 0 0.0004894400000000001 0 0.00048954 3.3 0.00048946 3.3 0.00048956 0 0.00048948 0 0.00048958 3.3 0.0004895 3.3 0.0004896 0 0.00048952 0 0.00048962 3.3 0.00048954 3.3 0.00048964 0 0.00048956 0 0.0004896599999999999 3.3 0.0004895800000000001 3.3 0.00048968 0 0.0004896000000000001 0 0.0004897 3.3 0.0004896200000000001 3.3 0.00048972 0 0.0004896400000000001 0 0.00048974 3.3 0.00048966 3.3 0.00048976 0 0.00048968 0 0.00048978 3.3 0.0004897 3.3 0.0004898 0 0.00048972 0 0.00048982 3.3 0.00048974 3.3 0.00048984 0 0.00048976 0 0.00048986 3.3 0.00048978 3.3 0.0004898799999999999 0 0.0004898000000000001 0 0.0004899 3.3 0.0004898200000000001 3.3 0.00048992 0 0.0004898400000000001 0 0.00048994 3.3 0.0004898600000000001 3.3 0.00048996 0 0.00048988 0 0.00048998 3.3 0.0004899 3.3 0.00049 0 0.00048992 0 0.00049002 3.3 0.00048994 3.3 0.00049004 0 0.00048996 0 0.00049006 3.3 0.00048998 3.3 0.0004900799999999999 0 0.0004900000000000001 0 0.0004901 3.3 0.0004900200000000001 3.3 0.00049012 0 0.0004900400000000001 0 0.00049014 3.3 0.0004900600000000001 3.3 0.00049016 0 0.00049008 0 0.00049018 3.3 0.0004901 3.3 0.0004902 0 0.00049012 0 0.00049022 3.3 0.00049014 3.3 0.00049024 0 0.00049016 0 0.00049026 3.3 0.00049018 3.3 0.00049028 0 0.0004902 0 0.0004902999999999999 3.3 0.0004902200000000001 3.3 0.00049032 0 0.0004902400000000001 0 0.00049034 3.3 0.0004902600000000001 3.3 0.00049036 0 0.0004902800000000001 0 0.00049038 3.3 0.0004903 3.3 0.0004904 0 0.00049032 0 0.00049042 3.3 0.00049034 3.3 0.00049044 0 0.00049036 0 0.00049046 3.3 0.00049038 3.3 0.00049048 0 0.0004904 0 0.0004904999999999999 3.3 0.0004904200000000001 3.3 0.00049052 0 0.0004904400000000001 0 0.00049054 3.3 0.0004904600000000001 3.3 0.00049056 0 0.0004904800000000001 0 0.00049058 3.3 0.0004905 3.3 0.0004906 0 0.00049052 0 0.00049062 3.3 0.00049054 3.3 0.00049064 0 0.00049056 0 0.00049066 3.3 0.00049058 3.3 0.00049068 0 0.0004906 0 0.0004907 3.3 0.00049062 3.3 0.0004907199999999999 0 0.0004906400000000001 0 0.00049074 3.3 0.0004906600000000001 3.3 0.00049076 0 0.0004906800000000001 0 0.00049078 3.3 0.0004907000000000001 3.3 0.0004908 0 0.00049072 0 0.00049082 3.3 0.00049074 3.3 0.00049084 0 0.00049076 0 0.00049086 3.3 0.00049078 3.3 0.00049088 0 0.0004908 0 0.0004909 3.3 0.00049082 3.3 0.0004909199999999999 0 0.0004908400000000001 0 0.00049094 3.3 0.0004908600000000001 3.3 0.00049096 0 0.0004908800000000001 0 0.00049098 3.3 0.0004909000000000001 3.3 0.000491 0 0.00049092 0 0.00049102 3.3 0.00049094 3.3 0.00049104 0 0.00049096 0 0.00049106 3.3 0.00049098 3.3 0.00049108 0 0.000491 0 0.0004911 3.3 0.00049102 3.3 0.00049112 0 0.00049104 0 0.0004911399999999999 3.3 0.0004910600000000001 3.3 0.00049116 0 0.0004910800000000001 0 0.00049118 3.3 0.0004911000000000001 3.3 0.0004912 0 0.0004911200000000001 0 0.00049122 3.3 0.00049114 3.3 0.00049124 0 0.00049116 0 0.00049126 3.3 0.00049118 3.3 0.00049128 0 0.0004912 0 0.0004913 3.3 0.00049122 3.3 0.00049132 0 0.00049124 0 0.0004913399999999999 3.3 0.0004912600000000001 3.3 0.00049136 0 0.0004912800000000001 0 0.00049138 3.3 0.0004913000000000001 3.3 0.0004914 0 0.0004913200000000001 0 0.00049142 3.3 0.00049134 3.3 0.00049144 0 0.00049136 0 0.00049146 3.3 0.00049138 3.3 0.00049148 0 0.0004914 0 0.0004915 3.3 0.00049142 3.3 0.00049152 0 0.00049144 0 0.0004915399999999999 3.3 0.0004914600000000001 3.3 0.00049156 0 0.0004914800000000001 0 0.00049158 3.3 0.0004915000000000001 3.3 0.0004916 0 0.0004915200000000001 0 0.00049162 3.3 0.00049154 3.3 0.00049164 0 0.00049156 0 0.00049166 3.3 0.00049158 3.3 0.00049168 0 0.0004916 0 0.0004917 3.3 0.00049162 3.3 0.00049172 0 0.00049164 0 0.00049174 3.3 0.00049166 3.3 0.0004917599999999999 0 0.0004916800000000001 0 0.00049178 3.3 0.0004917000000000001 3.3 0.0004918 0 0.0004917200000000001 0 0.00049182 3.3 0.0004917400000000001 3.3 0.00049184 0 0.00049176 0 0.00049186 3.3 0.00049178 3.3 0.00049188 0 0.0004918 0 0.0004919 3.3 0.00049182 3.3 0.00049192 0 0.00049184 0 0.00049194 3.3 0.00049186 3.3 0.0004919599999999999 0 0.0004918800000000001 0 0.00049198 3.3 0.0004919000000000001 3.3 0.000492 0 0.0004919200000000001 0 0.00049202 3.3 0.0004919400000000001 3.3 0.00049204 0 0.00049196 0 0.00049206 3.3 0.00049198 3.3 0.00049208 0 0.000492 0 0.0004921 3.3 0.00049202 3.3 0.00049212 0 0.00049204 0 0.00049214 3.3 0.00049206 3.3 0.00049216 0 0.00049208 0 0.0004921799999999999 3.3 0.0004921000000000001 3.3 0.0004922 0 0.0004921200000000001 0 0.00049222 3.3 0.0004921400000000001 3.3 0.00049224 0 0.0004921600000000001 0 0.00049226 3.3 0.00049218 3.3 0.00049228 0 0.0004922 0 0.0004923 3.3 0.00049222 3.3 0.00049232 0 0.00049224 0 0.00049234 3.3 0.00049226 3.3 0.00049236 0 0.00049228 0 0.0004923799999999999 3.3 0.0004923000000000001 3.3 0.0004924 0 0.0004923200000000001 0 0.00049242 3.3 0.0004923400000000001 3.3 0.00049244 0 0.0004923600000000001 0 0.00049246 3.3 0.00049238 3.3 0.00049248 0 0.0004924 0 0.0004925 3.3 0.00049242 3.3 0.00049252 0 0.00049244 0 0.00049254 3.3 0.00049246 3.3 0.00049256 0 0.00049248 0 0.00049258 3.3 0.0004925 3.3 0.0004925999999999999 0 0.0004925200000000001 0 0.00049262 3.3 0.0004925400000000001 3.3 0.00049264 0 0.0004925600000000001 0 0.00049266 3.3 0.0004925800000000001 3.3 0.00049268 0 0.0004926 0 0.0004927 3.3 0.00049262 3.3 0.00049272 0 0.00049264 0 0.00049274 3.3 0.00049266 3.3 0.00049276 0 0.00049268 0 0.00049278 3.3 0.0004927 3.3 0.0004927999999999999 0 0.0004927200000000001 0 0.00049282 3.3 0.0004927400000000001 3.3 0.00049284 0 0.0004927600000000001 0 0.00049286 3.3 0.0004927800000000001 3.3 0.00049288 0 0.0004928 0 0.0004929 3.3 0.00049282 3.3 0.00049292 0 0.00049284 0 0.00049294 3.3 0.00049286 3.3 0.00049296 0 0.00049288 0 0.00049298 3.3 0.0004929 3.3 0.000493 0 0.00049292 0 0.0004930199999999999 3.3 0.0004929400000000001 3.3 0.00049304 0 0.0004929600000000001 0 0.00049306 3.3 0.0004929800000000001 3.3 0.00049308 0 0.0004930000000000001 0 0.0004931 3.3 0.00049302 3.3 0.00049312 0 0.00049304 0 0.00049314 3.3 0.00049306 3.3 0.00049316 0 0.00049308 0 0.00049318 3.3 0.0004931 3.3 0.0004932 0 0.00049312 0 0.0004932199999999999 3.3 0.0004931400000000001 3.3 0.00049324 0 0.0004931600000000001 0 0.00049326 3.3 0.0004931800000000001 3.3 0.00049328 0 0.0004932000000000001 0 0.0004933 3.3 0.00049322 3.3 0.00049332 0 0.00049324 0 0.00049334 3.3 0.00049326 3.3 0.00049336 0 0.00049328 0 0.00049338 3.3 0.0004933 3.3 0.0004934 0 0.00049332 0 0.00049342 3.3 0.00049334 3.3 0.0004934399999999999 0 0.0004933600000000001 0 0.00049346 3.3 0.0004933800000000001 3.3 0.00049348 0 0.0004934000000000001 0 0.0004935 3.3 0.0004934200000000001 3.3 0.00049352 0 0.00049344 0 0.00049354 3.3 0.00049346 3.3 0.00049356 0 0.00049348 0 0.00049358 3.3 0.0004935 3.3 0.0004936 0 0.00049352 0 0.00049362 3.3 0.00049354 3.3 0.0004936399999999999 0 0.0004935600000000001 0 0.00049366 3.3 0.0004935800000000001 3.3 0.00049368 0 0.0004936000000000001 0 0.0004937 3.3 0.0004936200000000001 3.3 0.00049372 0 0.00049364 0 0.00049374 3.3 0.00049366 3.3 0.00049376 0 0.00049368 0 0.00049378 3.3 0.0004937 3.3 0.0004938 0 0.00049372 0 0.00049382 3.3 0.00049374 3.3 0.00049384 0 0.00049376 0 0.0004938599999999999 3.3 0.0004937800000000001 3.3 0.00049388 0 0.0004938000000000001 0 0.0004939 3.3 0.0004938200000000001 3.3 0.00049392 0 0.0004938400000000001 0 0.00049394 3.3 0.00049386 3.3 0.00049396 0 0.00049388 0 0.00049398 3.3 0.0004939 3.3 0.000494 0 0.00049392 0 0.00049402 3.3 0.00049394 3.3 0.00049404 0 0.00049396 0 0.0004940599999999999 3.3 0.0004939800000000001 3.3 0.00049408 0 0.0004940000000000001 0 0.0004941 3.3 0.0004940200000000001 3.3 0.00049412 0 0.0004940400000000001 0 0.00049414 3.3 0.00049406 3.3 0.00049416 0 0.00049408 0 0.00049418 3.3 0.0004941 3.3 0.0004942 0 0.00049412 0 0.00049422 3.3 0.00049414 3.3 0.00049424 0 0.00049416 0 0.00049426 3.3 0.00049418 3.3 0.0004942799999999999 0 0.0004942000000000001 0 0.0004943 3.3 0.0004942200000000001 3.3 0.00049432 0 0.0004942400000000001 0 0.00049434 3.3 0.0004942600000000001 3.3 0.00049436 0 0.00049428 0 0.00049438 3.3 0.0004943 3.3 0.0004944 0 0.00049432 0 0.00049442 3.3 0.00049434 3.3 0.00049444 0 0.00049436 0 0.00049446 3.3 0.00049438 3.3 0.0004944799999999999 0 0.0004944000000000001 0 0.0004945 3.3 0.0004944200000000001 3.3 0.00049452 0 0.0004944400000000001 0 0.00049454 3.3 0.0004944600000000001 3.3 0.00049456 0 0.00049448 0 0.00049458 3.3 0.0004945 3.3 0.0004946 0 0.00049452 0 0.00049462 3.3 0.00049454 3.3 0.00049464 0 0.00049456 0 0.00049466 3.3 0.00049458 3.3 0.00049468 0 0.0004946000000000001 0 0.0004947 3.3 0.0004946200000000001 3.3 0.00049472 0 0.0004946400000000001 0 0.00049474 3.3 0.0004946600000000001 3.3 0.00049476 0 0.0004946800000000001 0 0.00049478 3.3 0.0004947 3.3 0.0004948 0 0.00049472 0 0.00049482 3.3 0.00049474 3.3 0.00049484 0 0.00049476 0 0.00049486 3.3 0.00049478 3.3 0.00049488 0 0.0004948 0 0.0004948999999999999 3.3 0.0004948200000000001 3.3 0.00049492 0 0.0004948400000000001 0 0.00049494 3.3 0.0004948600000000001 3.3 0.00049496 0 0.0004948800000000001 0 0.00049498 3.3 0.0004949 3.3 0.000495 0 0.00049492 0 0.00049502 3.3 0.00049494 3.3 0.00049504 0 0.00049496 0 0.00049506 3.3 0.00049498 3.3 0.00049508 0 0.000495 0 0.0004950999999999999 3.3 0.0004950200000000001 3.3 0.00049512 0 0.0004950400000000001 0 0.00049514 3.3 0.0004950600000000001 3.3 0.00049516 0 0.0004950800000000001 0 0.00049518 3.3 0.0004951 3.3 0.0004952 0 0.00049512 0 0.00049522 3.3 0.00049514 3.3 0.00049524 0 0.00049516 0 0.00049526 3.3 0.00049518 3.3 0.00049528 0 0.0004952 0 0.0004953 3.3 0.00049522 3.3 0.0004953199999999999 0 0.0004952400000000001 0 0.00049534 3.3 0.0004952600000000001 3.3 0.00049536 0 0.0004952800000000001 0 0.00049538 3.3 0.0004953000000000001 3.3 0.0004954 0 0.00049532 0 0.00049542 3.3 0.00049534 3.3 0.00049544 0 0.00049536 0 0.00049546 3.3 0.00049538 3.3 0.00049548 0 0.0004954 0 0.0004955 3.3 0.00049542 3.3 0.0004955199999999999 0 0.0004954400000000001 0 0.00049554 3.3 0.0004954600000000001 3.3 0.00049556 0 0.0004954800000000001 0 0.00049558 3.3 0.0004955000000000001 3.3 0.0004956 0 0.00049552 0 0.00049562 3.3 0.00049554 3.3 0.00049564 0 0.00049556 0 0.00049566 3.3 0.00049558 3.3 0.00049568 0 0.0004956 0 0.0004957 3.3 0.00049562 3.3 0.00049572 0 0.00049564 0 0.0004957399999999999 3.3 0.0004956600000000001 3.3 0.00049576 0 0.0004956800000000001 0 0.00049578 3.3 0.0004957000000000001 3.3 0.0004958 0 0.0004957200000000001 0 0.00049582 3.3 0.00049574 3.3 0.00049584 0 0.00049576 0 0.00049586 3.3 0.00049578 3.3 0.00049588 0 0.0004958 0 0.0004959 3.3 0.00049582 3.3 0.00049592 0 0.00049584 0 0.0004959399999999999 3.3 0.0004958600000000001 3.3 0.00049596 0 0.0004958800000000001 0 0.00049598 3.3 0.0004959000000000001 3.3 0.000496 0 0.0004959200000000001 0 0.00049602 3.3 0.00049594 3.3 0.00049604 0 0.00049596 0 0.00049606 3.3 0.00049598 3.3 0.00049608 0 0.000496 0 0.0004961 3.3 0.00049602 3.3 0.00049612 0 0.00049604 0 0.00049614 3.3 0.00049606 3.3 0.0004961599999999999 0 0.0004960800000000001 0 0.00049618 3.3 0.0004961000000000001 3.3 0.0004962 0 0.0004961200000000001 0 0.00049622 3.3 0.0004961400000000001 3.3 0.00049624 0 0.00049616 0 0.00049626 3.3 0.00049618 3.3 0.00049628 0 0.0004962 0 0.0004963 3.3 0.00049622 3.3 0.00049632 0 0.00049624 0 0.00049634 3.3 0.00049626 3.3 0.0004963599999999999 0 0.0004962800000000001 0 0.00049638 3.3 0.0004963000000000001 3.3 0.0004964 0 0.0004963200000000001 0 0.00049642 3.3 0.0004963400000000001 3.3 0.00049644 0 0.00049636 0 0.00049646 3.3 0.00049638 3.3 0.00049648 0 0.0004964 0 0.0004965 3.3 0.00049642 3.3 0.00049652 0 0.00049644 0 0.00049654 3.3 0.00049646 3.3 0.00049656 0 0.00049648 0 0.0004965799999999999 3.3 0.0004965000000000001 3.3 0.0004966 0 0.0004965200000000001 0 0.00049662 3.3 0.0004965400000000001 3.3 0.00049664 0 0.0004965600000000001 0 0.00049666 3.3 0.00049658 3.3 0.00049668 0 0.0004966 0 0.0004967 3.3 0.00049662 3.3 0.00049672 0 0.00049664 0 0.00049674 3.3 0.00049666 3.3 0.00049676 0 0.00049668 0 0.0004967799999999999 3.3 0.0004967000000000001 3.3 0.0004968 0 0.0004967200000000001 0 0.00049682 3.3 0.0004967400000000001 3.3 0.00049684 0 0.0004967600000000001 0 0.00049686 3.3 0.00049678 3.3 0.00049688 0 0.0004968 0 0.0004969 3.3 0.00049682 3.3 0.00049692 0 0.00049684 0 0.00049694 3.3 0.00049686 3.3 0.00049696 0 0.00049688 0 0.00049698 3.3 0.0004969 3.3 0.0004969999999999999 0 0.0004969200000000001 0 0.00049702 3.3 0.0004969400000000001 3.3 0.00049704 0 0.0004969600000000001 0 0.00049706 3.3 0.0004969800000000001 3.3 0.00049708 0 0.000497 0 0.0004971 3.3 0.00049702 3.3 0.00049712 0 0.00049704 0 0.00049714 3.3 0.00049706 3.3 0.00049716 0 0.00049708 0 0.00049718 3.3 0.0004971 3.3 0.0004971999999999999 0 0.0004971200000000001 0 0.00049722 3.3 0.0004971400000000001 3.3 0.00049724 0 0.0004971600000000001 0 0.00049726 3.3 0.0004971800000000001 3.3 0.00049728 0 0.0004972 0 0.0004973 3.3 0.00049722 3.3 0.00049732 0 0.00049724 0 0.00049734 3.3 0.00049726 3.3 0.00049736 0 0.00049728 0 0.00049738 3.3 0.0004973 3.3 0.0004974 0 0.00049732 0 0.0004974199999999999 3.3 0.0004973400000000001 3.3 0.00049744 0 0.0004973600000000001 0 0.00049746 3.3 0.0004973800000000001 3.3 0.00049748 0 0.0004974000000000001 0 0.0004975 3.3 0.00049742 3.3 0.00049752 0 0.00049744 0 0.00049754 3.3 0.00049746 3.3 0.00049756 0 0.00049748 0 0.00049758 3.3 0.0004975 3.3 0.0004976 0 0.00049752 0 0.0004976199999999999 3.3 0.0004975400000000001 3.3 0.00049764 0 0.0004975600000000001 0 0.00049766 3.3 0.0004975800000000001 3.3 0.00049768 0 0.0004976000000000001 0 0.0004977 3.3 0.00049762 3.3 0.00049772 0 0.00049764 0 0.00049774 3.3 0.00049766 3.3 0.00049776 0 0.00049768 0 0.00049778 3.3 0.0004977 3.3 0.0004978 0 0.00049772 0 0.00049782 3.3 0.00049774 3.3 0.0004978399999999999 0 0.0004977600000000001 0 0.00049786 3.3 0.0004977800000000001 3.3 0.00049788 0 0.0004978000000000001 0 0.0004979 3.3 0.0004978200000000001 3.3 0.00049792 0 0.00049784 0 0.00049794 3.3 0.00049786 3.3 0.00049796 0 0.00049788 0 0.00049798 3.3 0.0004979 3.3 0.000498 0 0.00049792 0 0.00049802 3.3 0.00049794 3.3 0.0004980399999999999 0 0.0004979600000000001 0 0.00049806 3.3 0.0004979800000000001 3.3 0.00049808 0 0.0004980000000000001 0 0.0004981 3.3 0.0004980200000000001 3.3 0.00049812 0 0.00049804 0 0.00049814 3.3 0.00049806 3.3 0.00049816 0 0.00049808 0 0.00049818 3.3 0.0004981 3.3 0.0004982 0 0.00049812 0 0.00049822 3.3 0.00049814 3.3 0.00049824 0 0.0004981600000000001 0 0.00049826 3.3 0.0004981800000000001 3.3 0.00049828 0 0.0004982000000000001 0 0.0004983 3.3 0.0004982200000000001 3.3 0.00049832 0 0.0004982400000000001 0 0.00049834 3.3 0.00049826 3.3 0.00049836 0 0.00049828 0 0.00049838 3.3 0.0004983 3.3 0.0004984 0 0.00049832 0 0.00049842 3.3 0.00049834 3.3 0.00049844 0 0.00049836 0 0.0004984599999999999 3.3 0.0004983800000000001 3.3 0.00049848 0 0.0004984000000000001 0 0.0004985 3.3 0.0004984200000000001 3.3 0.00049852 0 0.0004984400000000001 0 0.00049854 3.3 0.00049846 3.3 0.00049856 0 0.00049848 0 0.00049858 3.3 0.0004985 3.3 0.0004986 0 0.00049852 0 0.00049862 3.3 0.00049854 3.3 0.00049864 0 0.00049856 0 0.0004986599999999999 3.3 0.0004985800000000001 3.3 0.00049868 0 0.0004986000000000001 0 0.0004987 3.3 0.0004986200000000001 3.3 0.00049872 0 0.0004986400000000001 0 0.00049874 3.3 0.00049866 3.3 0.00049876 0 0.00049868 0 0.00049878 3.3 0.0004987 3.3 0.0004988 0 0.00049872 0 0.00049882 3.3 0.00049874 3.3 0.00049884 0 0.00049876 0 0.00049886 3.3 0.00049878 3.3 0.0004988799999999999 0 0.0004988000000000001 0 0.0004989 3.3 0.0004988200000000001 3.3 0.00049892 0 0.0004988400000000001 0 0.00049894 3.3 0.0004988600000000001 3.3 0.00049896 0 0.00049888 0 0.00049898 3.3 0.0004989 3.3 0.000499 0 0.00049892 0 0.00049902 3.3 0.00049894 3.3 0.00049904 0 0.00049896 0 0.00049906 3.3 0.00049898 3.3 0.0004990799999999999 0 0.0004990000000000001 0 0.0004991 3.3 0.0004990200000000001 3.3 0.00049912 0 0.0004990400000000001 0 0.00049914 3.3 0.0004990600000000001 3.3 0.00049916 0 0.00049908 0 0.00049918 3.3 0.0004991 3.3 0.0004992 0 0.00049912 0 0.00049922 3.3 0.00049914 3.3 0.00049924 0 0.00049916 0 0.00049926 3.3 0.00049918 3.3 0.00049928 0 0.0004992 0 0.0004992999999999999 3.3 0.0004992200000000001 3.3 0.00049932 0 0.0004992400000000001 0 0.00049934 3.3 0.0004992600000000001 3.3 0.00049936 0 0.0004992800000000001 0 0.00049938 3.3 0.0004993 3.3 0.0004994 0 0.00049932 0 0.00049942 3.3 0.00049934 3.3 0.00049944 0 0.00049936 0 0.00049946 3.3 0.00049938 3.3 0.00049948 0 0.0004994 0 0.0004994999999999999 3.3 0.0004994200000000001 3.3 0.00049952 0 0.0004994400000000001 0 0.00049954 3.3 0.0004994600000000001 3.3 0.00049956 0 0.0004994800000000001 0 0.00049958 3.3 0.0004995 3.3 0.0004996 0 0.00049952 0 0.00049962 3.3 0.00049954 3.3 0.00049964 0 0.00049956 0 0.00049966 3.3 0.00049958 3.3 0.00049968 0 0.0004996 0 0.0004997 3.3 0.00049962 3.3 0.0004997199999999999 0 0.0004996400000000001 0 0.00049974 3.3 0.0004996600000000001 3.3 0.00049976 0 0.0004996800000000001 0 0.00049978 3.3 0.0004997000000000001 3.3 0.0004998 0 0.00049972 0 0.00049982 3.3 0.00049974 3.3 0.00049984 0 0.00049976 0 0.00049986 3.3 0.00049978 3.3 0.00049988 0 0.0004998 0 0.0004999 3.3 0.00049982 3.3 0.0004999199999999999 0 0.0004998400000000001 0 0.00049994 3.3 0.0004998600000000001 3.3 0.00049996 0 0.0004998800000000001 0 0.00049998 3.3 0.0004999000000000001 3.3 0.0005 0 0.00049992 0 0.00050002 3.3 0.00049994 3.3 0.00050004 0 0.00049996 0 0.00050006 3.3 0.00049998 3.3 0.00050008 0 0.0005 0 0.0005001 3.3 0.00050002 3.3 0.00050012 0 0.00050004 0 0.0005001399999999999 3.3 0.0005000600000000001 3.3 0.00050016 0 0.0005000800000000001 0 0.00050018 3.3 0.0005001000000000001 3.3 0.0005002 0 0.0005001200000000001 0 0.00050022 3.3 0.00050014 3.3 0.00050024 0 0.00050016 0 0.00050026 3.3 0.00050018 3.3 0.00050028 0 0.0005002 0 0.0005003 3.3 0.00050022 3.3 0.00050032 0 0.00050024 0 0.0005003399999999999 3.3 0.0005002600000000001 3.3 0.00050036 0 0.0005002800000000001 0 0.00050038 3.3 0.0005003000000000001 3.3 0.0005004 0 0.0005003200000000001 0 0.00050042 3.3 0.00050034 3.3 0.00050044 0 0.00050036 0 0.00050046 3.3 0.00050038 3.3 0.00050048 0 0.0005004 0 0.0005005 3.3 0.00050042 3.3 0.00050052 0 0.00050044 0 0.00050054 3.3 0.00050046 3.3 0.0005005599999999999 0 0.0005004800000000001 0 0.00050058 3.3 0.0005005000000000001 3.3 0.0005006 0 0.0005005200000000001 0 0.00050062 3.3 0.0005005400000000001 3.3 0.00050064 0 0.00050056 0 0.00050066 3.3 0.00050058 3.3 0.00050068 0 0.0005006 0 0.0005007 3.3 0.00050062 3.3 0.00050072 0 0.00050064 0 0.00050074 3.3 0.00050066 3.3 0.0005007599999999999 0 0.0005006800000000001 0 0.00050078 3.3 0.0005007000000000001 3.3 0.0005008 0 0.0005007200000000001 0 0.00050082 3.3 0.0005007400000000001 3.3 0.00050084 0 0.00050076 0 0.00050086 3.3 0.00050078 3.3 0.00050088 0 0.0005008 0 0.0005009 3.3 0.00050082 3.3 0.00050092 0 0.00050084 0 0.00050094 3.3 0.00050086 3.3 0.00050096 0 0.00050088 0 0.0005009799999999999 3.3 0.0005009000000000001 3.3 0.000501 0 0.0005009200000000001 0 0.00050102 3.3 0.0005009400000000001 3.3 0.00050104 0 0.0005009600000000001 0 0.00050106 3.3 0.00050098 3.3 0.00050108 0 0.000501 0 0.0005011 3.3 0.00050102 3.3 0.00050112 0 0.00050104 0 0.00050114 3.3 0.00050106 3.3 0.00050116 0 0.00050108 0 0.0005011799999999999 3.3 0.0005011000000000001 3.3 0.0005012 0 0.0005011200000000001 0 0.00050122 3.3 0.0005011400000000001 3.3 0.00050124 0 0.0005011600000000001 0 0.00050126 3.3 0.00050118 3.3 0.00050128 0 0.0005012 0 0.0005013 3.3 0.00050122 3.3 0.00050132 0 0.00050124 0 0.00050134 3.3 0.00050126 3.3 0.00050136 0 0.00050128 0 0.00050138 3.3 0.0005013 3.3 0.0005013999999999999 0 0.0005013200000000001 0 0.00050142 3.3 0.0005013400000000001 3.3 0.00050144 0 0.0005013600000000001 0 0.00050146 3.3 0.0005013800000000001 3.3 0.00050148 0 0.0005014 0 0.0005015 3.3 0.00050142 3.3 0.00050152 0 0.00050144 0 0.00050154 3.3 0.00050146 3.3 0.00050156 0 0.00050148 0 0.00050158 3.3 0.0005015 3.3 0.0005015999999999999 0 0.0005015200000000001 0 0.00050162 3.3 0.0005015400000000001 3.3 0.00050164 0 0.0005015600000000001 0 0.00050166 3.3 0.0005015800000000001 3.3 0.00050168 0 0.0005016 0 0.0005017 3.3 0.00050162 3.3 0.00050172 0 0.00050164 0 0.00050174 3.3 0.00050166 3.3 0.00050176 0 0.00050168 0 0.00050178 3.3 0.0005017 3.3 0.0005017999999999999 0 0.0005017200000000001 0 0.00050182 3.3 0.0005017400000000001 3.3 0.00050184 0 0.0005017600000000001 0 0.00050186 3.3 0.0005017800000000001 3.3 0.00050188 0 0.0005018 0 0.0005019 3.3 0.00050182 3.3 0.00050192 0 0.00050184 0 0.00050194 3.3 0.00050186 3.3 0.00050196 0 0.00050188 0 0.00050198 3.3 0.0005019 3.3 0.000502 0 0.00050192 0 0.0005020199999999999 3.3 0.0005019400000000001 3.3 0.00050204 0 0.0005019600000000001 0 0.00050206 3.3 0.0005019800000000001 3.3 0.00050208 0 0.0005020000000000001 0 0.0005021 3.3 0.00050202 3.3 0.00050212 0 0.00050204 0 0.00050214 3.3 0.00050206 3.3 0.00050216 0 0.00050208 0 0.00050218 3.3 0.0005021 3.3 0.0005022 0 0.00050212 0 0.0005022199999999999 3.3 0.0005021400000000001 3.3 0.00050224 0 0.0005021600000000001 0 0.00050226 3.3 0.0005021800000000001 3.3 0.00050228 0 0.0005022000000000001 0 0.0005023 3.3 0.00050222 3.3 0.00050232 0 0.00050224 0 0.00050234 3.3 0.00050226 3.3 0.00050236 0 0.00050228 0 0.00050238 3.3 0.0005023 3.3 0.0005024 0 0.00050232 0 0.00050242 3.3 0.00050234 3.3 0.0005024399999999999 0 0.0005023600000000001 0 0.00050246 3.3 0.0005023800000000001 3.3 0.00050248 0 0.0005024000000000001 0 0.0005025 3.3 0.0005024200000000001 3.3 0.00050252 0 0.00050244 0 0.00050254 3.3 0.00050246 3.3 0.00050256 0 0.00050248 0 0.00050258 3.3 0.0005025 3.3 0.0005026 0 0.00050252 0 0.00050262 3.3 0.00050254 3.3 0.0005026399999999999 0 0.0005025600000000001 0 0.00050266 3.3 0.0005025800000000001 3.3 0.00050268 0 0.0005026000000000001 0 0.0005027 3.3 0.0005026200000000001 3.3 0.00050272 0 0.00050264 0 0.00050274 3.3 0.00050266 3.3 0.00050276 0 0.00050268 0 0.00050278 3.3 0.0005027 3.3 0.0005028 0 0.00050272 0 0.00050282 3.3 0.00050274 3.3 0.00050284 0 0.00050276 0 0.0005028599999999999 3.3 0.0005027800000000001 3.3 0.00050288 0 0.0005028000000000001 0 0.0005029 3.3 0.0005028200000000001 3.3 0.00050292 0 0.0005028400000000001 0 0.00050294 3.3 0.00050286 3.3 0.00050296 0 0.00050288 0 0.00050298 3.3 0.0005029 3.3 0.000503 0 0.00050292 0 0.00050302 3.3 0.00050294 3.3 0.00050304 0 0.00050296 0 0.0005030599999999999 3.3 0.0005029800000000001 3.3 0.00050308 0 0.0005030000000000001 0 0.0005031 3.3 0.0005030200000000001 3.3 0.00050312 0 0.0005030400000000001 0 0.00050314 3.3 0.00050306 3.3 0.00050316 0 0.00050308 0 0.00050318 3.3 0.0005031 3.3 0.0005032 0 0.00050312 0 0.00050322 3.3 0.00050314 3.3 0.00050324 0 0.00050316 0 0.00050326 3.3 0.00050318 3.3 0.0005032799999999999 0 0.0005032000000000001 0 0.0005033 3.3 0.0005032200000000001 3.3 0.00050332 0 0.0005032400000000001 0 0.00050334 3.3 0.0005032600000000001 3.3 0.00050336 0 0.00050328 0 0.00050338 3.3 0.0005033 3.3 0.0005034 0 0.00050332 0 0.00050342 3.3 0.00050334 3.3 0.00050344 0 0.00050336 0 0.00050346 3.3 0.00050338 3.3 0.0005034799999999999 0 0.0005034000000000001 0 0.0005035 3.3 0.0005034200000000001 3.3 0.00050352 0 0.0005034400000000001 0 0.00050354 3.3 0.0005034600000000001 3.3 0.00050356 0 0.00050348 0 0.00050358 3.3 0.0005035 3.3 0.0005036 0 0.00050352 0 0.00050362 3.3 0.00050354 3.3 0.00050364 0 0.00050356 0 0.00050366 3.3 0.00050358 3.3 0.00050368 0 0.0005036 0 0.0005036999999999999 3.3 0.0005036200000000001 3.3 0.00050372 0 0.0005036400000000001 0 0.00050374 3.3 0.0005036600000000001 3.3 0.00050376 0 0.0005036800000000001 0 0.00050378 3.3 0.0005037 3.3 0.0005038 0 0.00050372 0 0.00050382 3.3 0.00050374 3.3 0.00050384 0 0.00050376 0 0.00050386 3.3 0.00050378 3.3 0.00050388 0 0.0005038 0 0.0005038999999999999 3.3 0.0005038200000000001 3.3 0.00050392 0 0.0005038400000000001 0 0.00050394 3.3 0.0005038600000000001 3.3 0.00050396 0 0.0005038800000000001 0 0.00050398 3.3 0.0005039 3.3 0.000504 0 0.00050392 0 0.00050402 3.3 0.00050394 3.3 0.00050404 0 0.00050396 0 0.00050406 3.3 0.00050398 3.3 0.00050408 0 0.000504 0 0.0005041 3.3 0.00050402 3.3 0.0005041199999999999 0 0.0005040400000000001 0 0.00050414 3.3 0.0005040600000000001 3.3 0.00050416 0 0.0005040800000000001 0 0.00050418 3.3 0.0005041000000000001 3.3 0.0005042 0 0.00050412 0 0.00050422 3.3 0.00050414 3.3 0.00050424 0 0.00050416 0 0.00050426 3.3 0.00050418 3.3 0.00050428 0 0.0005042 0 0.0005043 3.3 0.00050422 3.3 0.0005043199999999999 0 0.0005042400000000001 0 0.00050434 3.3 0.0005042600000000001 3.3 0.00050436 0 0.0005042800000000001 0 0.00050438 3.3 0.0005043000000000001 3.3 0.0005044 0 0.00050432 0 0.00050442 3.3 0.00050434 3.3 0.00050444 0 0.00050436 0 0.00050446 3.3 0.00050438 3.3 0.00050448 0 0.0005044 0 0.0005045 3.3 0.00050442 3.3 0.00050452 0 0.00050444 0 0.0005045399999999999 3.3 0.0005044600000000001 3.3 0.00050456 0 0.0005044800000000001 0 0.00050458 3.3 0.0005045000000000001 3.3 0.0005046 0 0.0005045200000000001 0 0.00050462 3.3 0.00050454 3.3 0.00050464 0 0.00050456 0 0.00050466 3.3 0.00050458 3.3 0.00050468 0 0.0005046 0 0.0005047 3.3 0.00050462 3.3 0.00050472 0 0.00050464 0 0.0005047399999999999 3.3 0.0005046600000000001 3.3 0.00050476 0 0.0005046800000000001 0 0.00050478 3.3 0.0005047000000000001 3.3 0.0005048 0 0.0005047200000000001 0 0.00050482 3.3 0.00050474 3.3 0.00050484 0 0.00050476 0 0.00050486 3.3 0.00050478 3.3 0.00050488 0 0.0005048 0 0.0005049 3.3 0.00050482 3.3 0.00050492 0 0.00050484 0 0.00050494 3.3 0.00050486 3.3 0.0005049599999999999 0 0.0005048800000000001 0 0.00050498 3.3 0.0005049000000000001 3.3 0.000505 0 0.0005049200000000001 0 0.00050502 3.3 0.0005049400000000001 3.3 0.00050504 0 0.00050496 0 0.00050506 3.3 0.00050498 3.3 0.00050508 0 0.000505 0 0.0005051 3.3 0.00050502 3.3 0.00050512 0 0.00050504 0 0.00050514 3.3 0.00050506 3.3 0.0005051599999999999 0 0.0005050800000000001 0 0.00050518 3.3 0.0005051000000000001 3.3 0.0005052 0 0.0005051200000000001 0 0.00050522 3.3 0.0005051400000000001 3.3 0.00050524 0 0.00050516 0 0.00050526 3.3 0.00050518 3.3 0.00050528 0 0.0005052 0 0.0005053 3.3 0.00050522 3.3 0.00050532 0 0.00050524 0 0.00050534 3.3 0.00050526 3.3 0.0005053599999999999 0 0.0005052800000000001 0 0.00050538 3.3 0.0005053000000000001 3.3 0.0005054 0 0.0005053200000000001 0 0.00050542 3.3 0.0005053400000000001 3.3 0.00050544 0 0.00050536 0 0.00050546 3.3 0.00050538 3.3 0.00050548 0 0.0005054 0 0.0005055 3.3 0.00050542 3.3 0.00050552 0 0.00050544 0 0.00050554 3.3 0.00050546 3.3 0.00050556 0 0.00050548 0 0.0005055799999999999 3.3 0.0005055000000000001 3.3 0.0005056 0 0.0005055200000000001 0 0.00050562 3.3 0.0005055400000000001 3.3 0.00050564 0 0.0005055600000000001 0 0.00050566 3.3 0.00050558 3.3 0.00050568 0 0.0005056 0 0.0005057 3.3 0.00050562 3.3 0.00050572 0 0.00050564 0 0.00050574 3.3 0.00050566 3.3 0.00050576 0 0.00050568 0 0.0005057799999999999 3.3 0.0005057000000000001 3.3 0.0005058 0 0.0005057200000000001 0 0.00050582 3.3 0.0005057400000000001 3.3 0.00050584 0 0.0005057600000000001 0 0.00050586 3.3 0.00050578 3.3 0.00050588 0 0.0005058 0 0.0005059 3.3 0.00050582 3.3 0.00050592 0 0.00050584 0 0.00050594 3.3 0.00050586 3.3 0.00050596 0 0.00050588 0 0.00050598 3.3 0.0005059 3.3 0.0005059999999999999 0 0.0005059200000000001 0 0.00050602 3.3 0.0005059400000000001 3.3 0.00050604 0 0.0005059600000000001 0 0.00050606 3.3 0.0005059800000000001 3.3 0.00050608 0 0.000506 0 0.0005061 3.3 0.00050602 3.3 0.00050612 0 0.00050604 0 0.00050614 3.3 0.00050606 3.3 0.00050616 0 0.00050608 0 0.00050618 3.3 0.0005061 3.3 0.0005061999999999999 0 0.0005061200000000001 0 0.00050622 3.3 0.0005061400000000001 3.3 0.00050624 0 0.0005061600000000001 0 0.00050626 3.3 0.0005061800000000001 3.3 0.00050628 0 0.0005062 0 0.0005063 3.3 0.00050622 3.3 0.00050632 0 0.00050624 0 0.00050634 3.3 0.00050626 3.3 0.00050636 0 0.00050628 0 0.00050638 3.3 0.0005063 3.3 0.0005064 0 0.00050632 0 0.0005064199999999999 3.3 0.0005063400000000001 3.3 0.00050644 0 0.0005063600000000001 0 0.00050646 3.3 0.0005063800000000001 3.3 0.00050648 0 0.0005064000000000001 0 0.0005065 3.3 0.00050642 3.3 0.00050652 0 0.00050644 0 0.00050654 3.3 0.00050646 3.3 0.00050656 0 0.00050648 0 0.00050658 3.3 0.0005065 3.3 0.0005066 0 0.00050652 0 0.0005066199999999999 3.3 0.0005065400000000001 3.3 0.00050664 0 0.0005065600000000001 0 0.00050666 3.3 0.0005065800000000001 3.3 0.00050668 0 0.0005066000000000001 0 0.0005067 3.3 0.00050662 3.3 0.00050672 0 0.00050664 0 0.00050674 3.3 0.00050666 3.3 0.00050676 0 0.00050668 0 0.00050678 3.3 0.0005067 3.3 0.0005068 0 0.00050672 0 0.00050682 3.3 0.00050674 3.3 0.0005068399999999999 0 0.0005067600000000001 0 0.00050686 3.3 0.0005067800000000001 3.3 0.00050688 0 0.0005068000000000001 0 0.0005069 3.3 0.0005068200000000001 3.3 0.00050692 0 0.00050684 0 0.00050694 3.3 0.00050686 3.3 0.00050696 0 0.00050688 0 0.00050698 3.3 0.0005069 3.3 0.000507 0 0.00050692 0 0.00050702 3.3 0.00050694 3.3 0.0005070399999999999 0 0.0005069600000000001 0 0.00050706 3.3 0.0005069800000000001 3.3 0.00050708 0 0.0005070000000000001 0 0.0005071 3.3 0.0005070200000000001 3.3 0.00050712 0 0.00050704 0 0.00050714 3.3 0.00050706 3.3 0.00050716 0 0.00050708 0 0.00050718 3.3 0.0005071 3.3 0.0005072 0 0.00050712 0 0.00050722 3.3 0.00050714 3.3 0.00050724 0 0.00050716 0 0.0005072599999999999 3.3 0.0005071800000000001 3.3 0.00050728 0 0.0005072000000000001 0 0.0005073 3.3 0.0005072200000000001 3.3 0.00050732 0 0.0005072400000000001 0 0.00050734 3.3 0.00050726 3.3 0.00050736 0 0.00050728 0 0.00050738 3.3 0.0005073 3.3 0.0005074 0 0.00050732 0 0.00050742 3.3 0.00050734 3.3 0.00050744 0 0.00050736 0 0.0005074599999999999 3.3 0.0005073800000000001 3.3 0.00050748 0 0.0005074000000000001 0 0.0005075 3.3 0.0005074200000000001 3.3 0.00050752 0 0.0005074400000000001 0 0.00050754 3.3 0.00050746 3.3 0.00050756 0 0.00050748 0 0.00050758 3.3 0.0005075 3.3 0.0005076 0 0.00050752 0 0.00050762 3.3 0.00050754 3.3 0.00050764 0 0.00050756 0 0.00050766 3.3 0.00050758 3.3 0.0005076799999999999 0 0.0005076000000000001 0 0.0005077 3.3 0.0005076200000000001 3.3 0.00050772 0 0.0005076400000000001 0 0.00050774 3.3 0.0005076600000000001 3.3 0.00050776 0 0.00050768 0 0.00050778 3.3 0.0005077 3.3 0.0005078 0 0.00050772 0 0.00050782 3.3 0.00050774 3.3 0.00050784 0 0.00050776 0 0.00050786 3.3 0.00050778 3.3 0.0005078799999999999 0 0.0005078000000000001 0 0.0005079 3.3 0.0005078200000000001 3.3 0.00050792 0 0.0005078400000000001 0 0.00050794 3.3 0.0005078600000000001 3.3 0.00050796 0 0.00050788 0 0.00050798 3.3 0.0005079 3.3 0.000508 0 0.00050792 0 0.00050802 3.3 0.00050794 3.3 0.00050804 0 0.00050796 0 0.00050806 3.3 0.00050798 3.3 0.00050808 0 0.000508 0 0.0005080999999999999 3.3 0.0005080200000000001 3.3 0.00050812 0 0.0005080400000000001 0 0.00050814 3.3 0.0005080600000000001 3.3 0.00050816 0 0.0005080800000000001 0 0.00050818 3.3 0.0005081 3.3 0.0005082 0 0.00050812 0 0.00050822 3.3 0.00050814 3.3 0.00050824 0 0.00050816 0 0.00050826 3.3 0.00050818 3.3 0.00050828 0 0.0005082 0 0.0005082999999999999 3.3 0.0005082200000000001 3.3 0.00050832 0 0.0005082400000000001 0 0.00050834 3.3 0.0005082600000000001 3.3 0.00050836 0 0.0005082800000000001 0 0.00050838 3.3 0.0005083 3.3 0.0005084 0 0.00050832 0 0.00050842 3.3 0.00050834 3.3 0.00050844 0 0.00050836 0 0.00050846 3.3 0.00050838 3.3 0.00050848 0 0.0005084 0 0.0005085 3.3 0.00050842 3.3 0.0005085199999999999 0 0.0005084400000000001 0 0.00050854 3.3 0.0005084600000000001 3.3 0.00050856 0 0.0005084800000000001 0 0.00050858 3.3 0.0005085000000000001 3.3 0.0005086 0 0.00050852 0 0.00050862 3.3 0.00050854 3.3 0.00050864 0 0.00050856 0 0.00050866 3.3 0.00050858 3.3 0.00050868 0 0.0005086 0 0.0005087 3.3 0.00050862 3.3 0.0005087199999999999 0 0.0005086400000000001 0 0.00050874 3.3 0.0005086600000000001 3.3 0.00050876 0 0.0005086800000000001 0 0.00050878 3.3 0.0005087000000000001 3.3 0.0005088 0 0.00050872 0 0.00050882 3.3 0.00050874 3.3 0.00050884 0 0.00050876 0 0.00050886 3.3 0.00050878 3.3 0.00050888 0 0.0005088 0 0.0005089 3.3 0.00050882 3.3 0.0005089199999999999 0 0.0005088400000000001 0 0.00050894 3.3 0.0005088600000000001 3.3 0.00050896 0 0.0005088800000000001 0 0.00050898 3.3 0.0005089000000000001 3.3 0.000509 0 0.00050892 0 0.00050902 3.3 0.00050894 3.3 0.00050904 0 0.00050896 0 0.00050906 3.3 0.00050898 3.3 0.00050908 0 0.000509 0 0.0005091 3.3 0.00050902 3.3 0.00050912 0 0.00050904 0 0.0005091399999999999 3.3 0.0005090600000000001 3.3 0.00050916 0 0.0005090800000000001 0 0.00050918 3.3 0.0005091000000000001 3.3 0.0005092 0 0.0005091200000000001 0 0.00050922 3.3 0.00050914 3.3 0.00050924 0 0.00050916 0 0.00050926 3.3 0.00050918 3.3 0.00050928 0 0.0005092 0 0.0005093 3.3 0.00050922 3.3 0.00050932 0 0.00050924 0 0.0005093399999999999 3.3 0.0005092600000000001 3.3 0.00050936 0 0.0005092800000000001 0 0.00050938 3.3 0.0005093000000000001 3.3 0.0005094 0 0.0005093200000000001 0 0.00050942 3.3 0.00050934 3.3 0.00050944 0 0.00050936 0 0.00050946 3.3 0.00050938 3.3 0.00050948 0 0.0005094 0 0.0005095 3.3 0.00050942 3.3 0.00050952 0 0.00050944 0 0.00050954 3.3 0.00050946 3.3 0.0005095599999999999 0 0.0005094800000000001 0 0.00050958 3.3 0.0005095000000000001 3.3 0.0005096 0 0.0005095200000000001 0 0.00050962 3.3 0.0005095400000000001 3.3 0.00050964 0 0.00050956 0 0.00050966 3.3 0.00050958 3.3 0.00050968 0 0.0005096 0 0.0005097 3.3 0.00050962 3.3 0.00050972 0 0.00050964 0 0.00050974 3.3 0.00050966 3.3 0.0005097599999999999 0 0.0005096800000000001 0 0.00050978 3.3 0.0005097000000000001 3.3 0.0005098 0 0.0005097200000000001 0 0.00050982 3.3 0.0005097400000000001 3.3 0.00050984 0 0.00050976 0 0.00050986 3.3 0.00050978 3.3 0.00050988 0 0.0005098 0 0.0005099 3.3 0.00050982 3.3 0.00050992 0 0.00050984 0 0.00050994 3.3 0.00050986 3.3 0.00050996 0 0.00050988 0 0.0005099799999999999 3.3 0.0005099000000000001 3.3 0.00051 0 0.0005099200000000001 0 0.00051002 3.3 0.0005099400000000001 3.3 0.00051004 0 0.0005099600000000001 0 0.00051006 3.3 0.00050998 3.3 0.00051008 0 0.00051 0 0.0005101 3.3 0.00051002 3.3 0.00051012 0 0.00051004 0 0.00051014 3.3 0.00051006 3.3 0.00051016 0 0.00051008 0 0.0005101799999999999 3.3 0.0005101000000000001 3.3 0.0005102 0 0.0005101200000000001 0 0.00051022 3.3 0.0005101400000000001 3.3 0.00051024 0 0.0005101600000000001 0 0.00051026 3.3 0.00051018 3.3 0.00051028 0 0.0005102 0 0.0005103 3.3 0.00051022 3.3 0.00051032 0 0.00051024 0 0.00051034 3.3 0.00051026 3.3 0.00051036 0 0.00051028 0 0.00051038 3.3 0.0005103 3.3 0.0005103999999999999 0 0.0005103200000000001 0 0.00051042 3.3 0.0005103400000000001 3.3 0.00051044 0 0.0005103600000000001 0 0.00051046 3.3 0.0005103800000000001 3.3 0.00051048 0 0.0005104 0 0.0005105 3.3 0.00051042 3.3 0.00051052 0 0.00051044 0 0.00051054 3.3 0.00051046 3.3 0.00051056 0 0.00051048 0 0.00051058 3.3 0.0005105 3.3 0.0005105999999999999 0 0.0005105200000000001 0 0.00051062 3.3 0.0005105400000000001 3.3 0.00051064 0 0.0005105600000000001 0 0.00051066 3.3 0.0005105800000000001 3.3 0.00051068 0 0.0005106 0 0.0005107 3.3 0.00051062 3.3 0.00051072 0 0.00051064 0 0.00051074 3.3 0.00051066 3.3 0.00051076 0 0.00051068 0 0.00051078 3.3 0.0005107 3.3 0.0005108 0 0.00051072 0 0.0005108199999999999 3.3 0.0005107400000000001 3.3 0.00051084 0 0.0005107600000000001 0 0.00051086 3.3 0.0005107800000000001 3.3 0.00051088 0 0.0005108000000000001 0 0.0005109 3.3 0.00051082 3.3 0.00051092 0 0.00051084 0 0.00051094 3.3 0.00051086 3.3 0.00051096 0 0.00051088 0 0.00051098 3.3 0.0005109 3.3 0.000511 0 0.00051092 0 0.0005110199999999999 3.3 0.0005109400000000001 3.3 0.00051104 0 0.0005109600000000001 0 0.00051106 3.3 0.0005109800000000001 3.3 0.00051108 0 0.0005110000000000001 0 0.0005111 3.3 0.00051102 3.3 0.00051112 0 0.00051104 0 0.00051114 3.3 0.00051106 3.3 0.00051116 0 0.00051108 0 0.00051118 3.3 0.0005111 3.3 0.0005112 0 0.00051112 0 0.00051122 3.3 0.00051114 3.3 0.0005112399999999999 0 0.0005111600000000001 0 0.00051126 3.3 0.0005111800000000001 3.3 0.00051128 0 0.0005112000000000001 0 0.0005113 3.3 0.0005112200000000001 3.3 0.00051132 0 0.00051124 0 0.00051134 3.3 0.00051126 3.3 0.00051136 0 0.00051128 0 0.00051138 3.3 0.0005113 3.3 0.0005114 0 0.00051132 0 0.00051142 3.3 0.00051134 3.3 0.0005114399999999999 0 0.0005113600000000001 0 0.00051146 3.3 0.0005113800000000001 3.3 0.00051148 0 0.0005114000000000001 0 0.0005115 3.3 0.0005114200000000001 3.3 0.00051152 0 0.00051144 0 0.00051154 3.3 0.00051146 3.3 0.00051156 0 0.00051148 0 0.00051158 3.3 0.0005115 3.3 0.0005116 0 0.00051152 0 0.00051162 3.3 0.00051154 3.3 0.00051164 0 0.00051156 0 0.0005116599999999999 3.3 0.0005115800000000001 3.3 0.00051168 0 0.0005116000000000001 0 0.0005117 3.3 0.0005116200000000001 3.3 0.00051172 0 0.0005116400000000001 0 0.00051174 3.3 0.00051166 3.3 0.00051176 0 0.00051168 0 0.00051178 3.3 0.0005117 3.3 0.0005118 0 0.00051172 0 0.00051182 3.3 0.00051174 3.3 0.00051184 0 0.00051176 0 0.0005118599999999999 3.3 0.0005117800000000001 3.3 0.00051188 0 0.0005118000000000001 0 0.0005119 3.3 0.0005118200000000001 3.3 0.00051192 0 0.0005118400000000001 0 0.00051194 3.3 0.00051186 3.3 0.00051196 0 0.00051188 0 0.00051198 3.3 0.0005119 3.3 0.000512 0 0.00051192 0 0.00051202 3.3 0.00051194 3.3 0.00051204 0 0.00051196 0 0.0005120599999999999 3.3 0.0005119800000000001 3.3 0.00051208 0 0.0005120000000000001 0 0.0005121 3.3 0.0005120200000000001 3.3 0.00051212 0 0.0005120400000000001 0 0.00051214 3.3 0.00051206 3.3 0.00051216 0 0.00051208 0 0.00051218 3.3 0.0005121 3.3 0.0005122 0 0.00051212 0 0.00051222 3.3 0.00051214 3.3 0.00051224 0 0.00051216 0 0.00051226 3.3 0.00051218 3.3 0.0005122799999999999 0 0.0005122000000000001 0 0.0005123 3.3 0.0005122200000000001 3.3 0.00051232 0 0.0005122400000000001 0 0.00051234 3.3 0.0005122600000000001 3.3 0.00051236 0 0.00051228 0 0.00051238 3.3 0.0005123 3.3 0.0005124 0 0.00051232 0 0.00051242 3.3 0.00051234 3.3 0.00051244 0 0.00051236 0 0.00051246 3.3 0.00051238 3.3 0.0005124799999999999 0 0.0005124000000000001 0 0.0005125 3.3 0.0005124200000000001 3.3 0.00051252 0 0.0005124400000000001 0 0.00051254 3.3 0.0005124600000000001 3.3 0.00051256 0 0.00051248 0 0.00051258 3.3 0.0005125 3.3 0.0005126 0 0.00051252 0 0.00051262 3.3 0.00051254 3.3 0.00051264 0 0.00051256 0 0.00051266 3.3 0.00051258 3.3 0.00051268 0 0.0005126 0 0.0005126999999999999 3.3 0.0005126200000000001 3.3 0.00051272 0 0.0005126400000000001 0 0.00051274 3.3 0.0005126600000000001 3.3 0.00051276 0 0.0005126800000000001 0 0.00051278 3.3 0.0005127 3.3 0.0005128 0 0.00051272 0 0.00051282 3.3 0.00051274 3.3 0.00051284 0 0.00051276 0 0.00051286 3.3 0.00051278 3.3 0.00051288 0 0.0005128 0 0.0005128999999999999 3.3 0.0005128200000000001 3.3 0.00051292 0 0.0005128400000000001 0 0.00051294 3.3 0.0005128600000000001 3.3 0.00051296 0 0.0005128800000000001 0 0.00051298 3.3 0.0005129 3.3 0.000513 0 0.00051292 0 0.00051302 3.3 0.00051294 3.3 0.00051304 0 0.00051296 0 0.00051306 3.3 0.00051298 3.3 0.00051308 0 0.000513 0 0.0005131 3.3 0.00051302 3.3 0.0005131199999999999 0 0.0005130400000000001 0 0.00051314 3.3 0.0005130600000000001 3.3 0.00051316 0 0.0005130800000000001 0 0.00051318 3.3 0.0005131000000000001 3.3 0.0005132 0 0.00051312 0 0.00051322 3.3 0.00051314 3.3 0.00051324 0 0.00051316 0 0.00051326 3.3 0.00051318 3.3 0.00051328 0 0.0005132 0 0.0005133 3.3 0.00051322 3.3 0.0005133199999999999 0 0.0005132400000000001 0 0.00051334 3.3 0.0005132600000000001 3.3 0.00051336 0 0.0005132800000000001 0 0.00051338 3.3 0.0005133000000000001 3.3 0.0005134 0 0.00051332 0 0.00051342 3.3 0.00051334 3.3 0.00051344 0 0.00051336 0 0.00051346 3.3 0.00051338 3.3 0.00051348 0 0.0005134 0 0.0005135 3.3 0.00051342 3.3 0.00051352 0 0.00051344 0 0.0005135399999999999 3.3 0.0005134600000000001 3.3 0.00051356 0 0.0005134800000000001 0 0.00051358 3.3 0.0005135000000000001 3.3 0.0005136 0 0.0005135200000000001 0 0.00051362 3.3 0.00051354 3.3 0.00051364 0 0.00051356 0 0.00051366 3.3 0.00051358 3.3 0.00051368 0 0.0005136 0 0.0005137 3.3 0.00051362 3.3 0.00051372 0 0.00051364 0 0.0005137399999999999 3.3 0.0005136600000000001 3.3 0.00051376 0 0.0005136800000000001 0 0.00051378 3.3 0.0005137000000000001 3.3 0.0005138 0 0.0005137200000000001 0 0.00051382 3.3 0.00051374 3.3 0.00051384 0 0.00051376 0 0.00051386 3.3 0.00051378 3.3 0.00051388 0 0.0005138 0 0.0005139 3.3 0.00051382 3.3 0.00051392 0 0.00051384 0 0.00051394 3.3 0.00051386 3.3 0.0005139599999999999 0 0.0005138800000000001 0 0.00051398 3.3 0.0005139000000000001 3.3 0.000514 0 0.0005139200000000001 0 0.00051402 3.3 0.0005139400000000001 3.3 0.00051404 0 0.00051396 0 0.00051406 3.3 0.00051398 3.3 0.00051408 0 0.000514 0 0.0005141 3.3 0.00051402 3.3 0.00051412 0 0.00051404 0 0.00051414 3.3 0.00051406 3.3 0.0005141599999999999 0 0.0005140800000000001 0 0.00051418 3.3 0.0005141000000000001 3.3 0.0005142 0 0.0005141200000000001 0 0.00051422 3.3 0.0005141400000000001 3.3 0.00051424 0 0.00051416 0 0.00051426 3.3 0.00051418 3.3 0.00051428 0 0.0005142 0 0.0005143 3.3 0.00051422 3.3 0.00051432 0 0.00051424 0 0.00051434 3.3 0.00051426 3.3 0.00051436 0 0.00051428 0 0.0005143799999999999 3.3 0.0005143000000000001 3.3 0.0005144 0 0.0005143200000000001 0 0.00051442 3.3 0.0005143400000000001 3.3 0.00051444 0 0.0005143600000000001 0 0.00051446 3.3 0.00051438 3.3 0.00051448 0 0.0005144 0 0.0005145 3.3 0.00051442 3.3 0.00051452 0 0.00051444 0 0.00051454 3.3 0.00051446 3.3 0.00051456 0 0.00051448 0 0.0005145799999999999 3.3 0.0005145000000000001 3.3 0.0005146 0 0.0005145200000000001 0 0.00051462 3.3 0.0005145400000000001 3.3 0.00051464 0 0.0005145600000000001 0 0.00051466 3.3 0.00051458 3.3 0.00051468 0 0.0005146 0 0.0005147 3.3 0.00051462 3.3 0.00051472 0 0.00051464 0 0.00051474 3.3 0.00051466 3.3 0.00051476 0 0.00051468 0 0.00051478 3.3 0.0005147 3.3 0.0005147999999999999 0 0.0005147200000000001 0 0.00051482 3.3 0.0005147400000000001 3.3 0.00051484 0 0.0005147600000000001 0 0.00051486 3.3 0.0005147800000000001 3.3 0.00051488 0 0.0005148 0 0.0005149 3.3 0.00051482 3.3 0.00051492 0 0.00051484 0 0.00051494 3.3 0.00051486 3.3 0.00051496 0 0.00051488 0 0.00051498 3.3 0.0005149 3.3 0.0005149999999999999 0 0.0005149200000000001 0 0.00051502 3.3 0.0005149400000000001 3.3 0.00051504 0 0.0005149600000000001 0 0.00051506 3.3 0.0005149800000000001 3.3 0.00051508 0 0.000515 0 0.0005151 3.3 0.00051502 3.3 0.00051512 0 0.00051504 0 0.00051514 3.3 0.00051506 3.3 0.00051516 0 0.00051508 0 0.00051518 3.3 0.0005151 3.3 0.0005152 0 0.00051512 0 0.0005152199999999999 3.3 0.0005151400000000001 3.3 0.00051524 0 0.0005151600000000001 0 0.00051526 3.3 0.0005151800000000001 3.3 0.00051528 0 0.0005152000000000001 0 0.0005153 3.3 0.00051522 3.3 0.00051532 0 0.00051524 0 0.00051534 3.3 0.00051526 3.3 0.00051536 0 0.00051528 0 0.00051538 3.3 0.0005153 3.3 0.0005154 0 0.00051532 0 0.0005154199999999999 3.3 0.0005153400000000001 3.3 0.00051544 0 0.0005153600000000001 0 0.00051546 3.3 0.0005153800000000001 3.3 0.00051548 0 0.0005154000000000001 0 0.0005155 3.3 0.00051542 3.3 0.00051552 0 0.00051544 0 0.00051554 3.3 0.00051546 3.3 0.00051556 0 0.00051548 0 0.00051558 3.3 0.0005155 3.3 0.0005156 0 0.00051552 0 0.0005156199999999999 3.3 0.0005155400000000001 3.3 0.00051564 0 0.0005155600000000001 0 0.00051566 3.3 0.0005155800000000001 3.3 0.00051568 0 0.0005156000000000001 0 0.0005157 3.3 0.00051562 3.3 0.00051572 0 0.00051564 0 0.00051574 3.3 0.00051566 3.3 0.00051576 0 0.00051568 0 0.00051578 3.3 0.0005157 3.3 0.0005158 0 0.00051572 0 0.00051582 3.3 0.00051574 3.3 0.0005158399999999999 0 0.0005157600000000001 0 0.00051586 3.3 0.0005157800000000001 3.3 0.00051588 0 0.0005158000000000001 0 0.0005159 3.3 0.0005158200000000001 3.3 0.00051592 0 0.00051584 0 0.00051594 3.3 0.00051586 3.3 0.00051596 0 0.00051588 0 0.00051598 3.3 0.0005159 3.3 0.000516 0 0.00051592 0 0.00051602 3.3 0.00051594 3.3 0.0005160399999999999 0 0.0005159600000000001 0 0.00051606 3.3 0.0005159800000000001 3.3 0.00051608 0 0.0005160000000000001 0 0.0005161 3.3 0.0005160200000000001 3.3 0.00051612 0 0.00051604 0 0.00051614 3.3 0.00051606 3.3 0.00051616 0 0.00051608 0 0.00051618 3.3 0.0005161 3.3 0.0005162 0 0.00051612 0 0.00051622 3.3 0.00051614 3.3 0.00051624 0 0.00051616 0 0.0005162599999999999 3.3 0.0005161800000000001 3.3 0.00051628 0 0.0005162000000000001 0 0.0005163 3.3 0.0005162200000000001 3.3 0.00051632 0 0.0005162400000000001 0 0.00051634 3.3 0.00051626 3.3 0.00051636 0 0.00051628 0 0.00051638 3.3 0.0005163 3.3 0.0005164 0 0.00051632 0 0.00051642 3.3 0.00051634 3.3 0.00051644 0 0.00051636 0 0.0005164599999999999 3.3 0.0005163800000000001 3.3 0.00051648 0 0.0005164000000000001 0 0.0005165 3.3 0.0005164200000000001 3.3 0.00051652 0 0.0005164400000000001 0 0.00051654 3.3 0.00051646 3.3 0.00051656 0 0.00051648 0 0.00051658 3.3 0.0005165 3.3 0.0005166 0 0.00051652 0 0.00051662 3.3 0.00051654 3.3 0.00051664 0 0.00051656 0 0.00051666 3.3 0.00051658 3.3 0.0005166799999999999 0 0.0005166000000000001 0 0.0005167 3.3 0.0005166200000000001 3.3 0.00051672 0 0.0005166400000000001 0 0.00051674 3.3 0.0005166600000000001 3.3 0.00051676 0 0.00051668 0 0.00051678 3.3 0.0005167 3.3 0.0005168 0 0.00051672 0 0.00051682 3.3 0.00051674 3.3 0.00051684 0 0.00051676 0 0.00051686 3.3 0.00051678 3.3 0.0005168799999999999 0 0.0005168000000000001 0 0.0005169 3.3 0.0005168200000000001 3.3 0.00051692 0 0.0005168400000000001 0 0.00051694 3.3 0.0005168600000000001 3.3 0.00051696 0 0.00051688 0 0.00051698 3.3 0.0005169 3.3 0.000517 0 0.00051692 0 0.00051702 3.3 0.00051694 3.3 0.00051704 0 0.00051696 0 0.00051706 3.3 0.00051698 3.3 0.00051708 0 0.000517 0 0.0005170999999999999 3.3 0.0005170200000000001 3.3 0.00051712 0 0.0005170400000000001 0 0.00051714 3.3 0.0005170600000000001 3.3 0.00051716 0 0.0005170800000000001 0 0.00051718 3.3 0.0005171 3.3 0.0005172 0 0.00051712 0 0.00051722 3.3 0.00051714 3.3 0.00051724 0 0.00051716 0 0.00051726 3.3 0.00051718 3.3 0.00051728 0 0.0005172 0 0.0005172999999999999 3.3 0.0005172200000000001 3.3 0.00051732 0 0.0005172400000000001 0 0.00051734 3.3 0.0005172600000000001 3.3 0.00051736 0 0.0005172800000000001 0 0.00051738 3.3 0.0005173 3.3 0.0005174 0 0.00051732 0 0.00051742 3.3 0.00051734 3.3 0.00051744 0 0.00051736 0 0.00051746 3.3 0.00051738 3.3 0.00051748 0 0.0005174 0 0.0005175 3.3 0.00051742 3.3 0.0005175199999999999 0 0.0005174400000000001 0 0.00051754 3.3 0.0005174600000000001 3.3 0.00051756 0 0.0005174800000000001 0 0.00051758 3.3 0.0005175000000000001 3.3 0.0005176 0 0.00051752 0 0.00051762 3.3 0.00051754 3.3 0.00051764 0 0.00051756 0 0.00051766 3.3 0.00051758 3.3 0.00051768 0 0.0005176 0 0.0005177 3.3 0.00051762 3.3 0.0005177199999999999 0 0.0005176400000000001 0 0.00051774 3.3 0.0005176600000000001 3.3 0.00051776 0 0.0005176800000000001 0 0.00051778 3.3 0.0005177000000000001 3.3 0.0005178 0 0.00051772 0 0.00051782 3.3 0.00051774 3.3 0.00051784 0 0.00051776 0 0.00051786 3.3 0.00051778 3.3 0.00051788 0 0.0005178 0 0.0005179 3.3 0.00051782 3.3 0.00051792 0 0.00051784 0 0.0005179399999999999 3.3 0.0005178600000000001 3.3 0.00051796 0 0.0005178800000000001 0 0.00051798 3.3 0.0005179000000000001 3.3 0.000518 0 0.0005179200000000001 0 0.00051802 3.3 0.00051794 3.3 0.00051804 0 0.00051796 0 0.00051806 3.3 0.00051798 3.3 0.00051808 0 0.000518 0 0.0005181 3.3 0.00051802 3.3 0.00051812 0 0.00051804 0 0.0005181399999999999 3.3 0.0005180600000000001 3.3 0.00051816 0 0.0005180800000000001 0 0.00051818 3.3 0.0005181000000000001 3.3 0.0005182 0 0.0005181200000000001 0 0.00051822 3.3 0.00051814 3.3 0.00051824 0 0.00051816 0 0.00051826 3.3 0.00051818 3.3 0.00051828 0 0.0005182 0 0.0005183 3.3 0.00051822 3.3 0.00051832 0 0.00051824 0 0.00051834 3.3 0.00051826 3.3 0.0005183599999999999 0 0.0005182800000000001 0 0.00051838 3.3 0.0005183000000000001 3.3 0.0005184 0 0.0005183200000000001 0 0.00051842 3.3 0.0005183400000000001 3.3 0.00051844 0 0.00051836 0 0.00051846 3.3 0.00051838 3.3 0.00051848 0 0.0005184 0 0.0005185 3.3 0.00051842 3.3 0.00051852 0 0.00051844 0 0.00051854 3.3 0.00051846 3.3 0.0005185599999999999 0 0.0005184800000000001 0 0.00051858 3.3 0.0005185000000000001 3.3 0.0005186 0 0.0005185200000000001 0 0.00051862 3.3 0.0005185400000000001 3.3 0.00051864 0 0.00051856 0 0.00051866 3.3 0.00051858 3.3 0.00051868 0 0.0005186 0 0.0005187 3.3 0.00051862 3.3 0.00051872 0 0.00051864 0 0.00051874 3.3 0.00051866 3.3 0.00051876 0 0.00051868 0 0.0005187799999999999 3.3 0.0005187000000000001 3.3 0.0005188 0 0.0005187200000000001 0 0.00051882 3.3 0.0005187400000000001 3.3 0.00051884 0 0.0005187600000000001 0 0.00051886 3.3 0.00051878 3.3 0.00051888 0 0.0005188 0 0.0005189 3.3 0.00051882 3.3 0.00051892 0 0.00051884 0 0.00051894 3.3 0.00051886 3.3 0.00051896 0 0.00051888 0 0.0005189799999999999 3.3 0.0005189000000000001 3.3 0.000519 0 0.0005189200000000001 0 0.00051902 3.3 0.0005189400000000001 3.3 0.00051904 0 0.0005189600000000001 0 0.00051906 3.3 0.00051898 3.3 0.00051908 0 0.000519 0 0.0005191 3.3 0.00051902 3.3 0.00051912 0 0.00051904 0 0.00051914 3.3 0.00051906 3.3 0.00051916 0 0.00051908 0 0.0005191799999999999 3.3 0.0005191000000000001 3.3 0.0005192 0 0.0005191200000000001 0 0.00051922 3.3 0.0005191400000000001 3.3 0.00051924 0 0.0005191600000000001 0 0.00051926 3.3 0.00051918 3.3 0.00051928 0 0.0005192 0 0.0005193 3.3 0.00051922 3.3 0.00051932 0 0.00051924 0 0.00051934 3.3 0.00051926 3.3 0.00051936 0 0.00051928 0 0.00051938 3.3 0.0005193 3.3 0.0005193999999999999 0 0.0005193200000000001 0 0.00051942 3.3 0.0005193400000000001 3.3 0.00051944 0 0.0005193600000000001 0 0.00051946 3.3 0.0005193800000000001 3.3 0.00051948 0 0.0005194 0 0.0005195 3.3 0.00051942 3.3 0.00051952 0 0.00051944 0 0.00051954 3.3 0.00051946 3.3 0.00051956 0 0.00051948 0 0.00051958 3.3 0.0005195 3.3 0.0005195999999999999 0 0.0005195200000000001 0 0.00051962 3.3 0.0005195400000000001 3.3 0.00051964 0 0.0005195600000000001 0 0.00051966 3.3 0.0005195800000000001 3.3 0.00051968 0 0.0005196 0 0.0005197 3.3 0.00051962 3.3 0.00051972 0 0.00051964 0 0.00051974 3.3 0.00051966 3.3 0.00051976 0 0.00051968 0 0.00051978 3.3 0.0005197 3.3 0.0005198 0 0.00051972 0 0.0005198199999999999 3.3 0.0005197400000000001 3.3 0.00051984 0 0.0005197600000000001 0 0.00051986 3.3 0.0005197800000000001 3.3 0.00051988 0 0.0005198000000000001 0 0.0005199 3.3 0.00051982 3.3 0.00051992 0 0.00051984 0 0.00051994 3.3 0.00051986 3.3 0.00051996 0 0.00051988 0 0.00051998 3.3 0.0005199 3.3 0.00052 0 0.00051992 0 0.0005200199999999999 3.3 0.0005199400000000001 3.3 0.00052004 0 0.0005199600000000001 0 0.00052006 3.3 0.0005199800000000001 3.3 0.00052008 0 0.0005200000000000001 0 0.0005201 3.3 0.00052002 3.3 0.00052012 0 0.00052004 0 0.00052014 3.3 0.00052006 3.3 0.00052016 0 0.00052008 0 0.00052018 3.3 0.0005201 3.3 0.0005202 0 0.00052012 0 0.00052022 3.3 0.00052014 3.3 0.0005202399999999999 0 0.0005201600000000001 0 0.00052026 3.3 0.0005201800000000001 3.3 0.00052028 0 0.0005202000000000001 0 0.0005203 3.3 0.0005202200000000001 3.3 0.00052032 0 0.00052024 0 0.00052034 3.3 0.00052026 3.3 0.00052036 0 0.00052028 0 0.00052038 3.3 0.0005203 3.3 0.0005204 0 0.00052032 0 0.00052042 3.3 0.00052034 3.3 0.0005204399999999999 0 0.0005203600000000001 0 0.00052046 3.3 0.0005203800000000001 3.3 0.00052048 0 0.0005204000000000001 0 0.0005205 3.3 0.0005204200000000001 3.3 0.00052052 0 0.00052044 0 0.00052054 3.3 0.00052046 3.3 0.00052056 0 0.00052048 0 0.00052058 3.3 0.0005205 3.3 0.0005206 0 0.00052052 0 0.00052062 3.3 0.00052054 3.3 0.00052064 0 0.00052056 0 0.0005206599999999999 3.3 0.0005205800000000001 3.3 0.00052068 0 0.0005206000000000001 0 0.0005207 3.3 0.0005206200000000001 3.3 0.00052072 0 0.0005206400000000001 0 0.00052074 3.3 0.00052066 3.3 0.00052076 0 0.00052068 0 0.00052078 3.3 0.0005207 3.3 0.0005208 0 0.00052072 0 0.00052082 3.3 0.00052074 3.3 0.00052084 0 0.00052076 0 0.0005208599999999999 3.3 0.0005207800000000001 3.3 0.00052088 0 0.0005208000000000001 0 0.0005209 3.3 0.0005208200000000001 3.3 0.00052092 0 0.0005208400000000001 0 0.00052094 3.3 0.00052086 3.3 0.00052096 0 0.00052088 0 0.00052098 3.3 0.0005209 3.3 0.000521 0 0.00052092 0 0.00052102 3.3 0.00052094 3.3 0.00052104 0 0.00052096 0 0.00052106 3.3 0.00052098 3.3 0.0005210799999999999 0 0.0005210000000000001 0 0.0005211 3.3 0.0005210200000000001 3.3 0.00052112 0 0.0005210400000000001 0 0.00052114 3.3 0.0005210600000000001 3.3 0.00052116 0 0.00052108 0 0.00052118 3.3 0.0005211 3.3 0.0005212 0 0.00052112 0 0.00052122 3.3 0.00052114 3.3 0.00052124 0 0.00052116 0 0.00052126 3.3 0.00052118 3.3 0.0005212799999999999 0 0.0005212000000000001 0 0.0005213 3.3 0.0005212200000000001 3.3 0.00052132 0 0.0005212400000000001 0 0.00052134 3.3 0.0005212600000000001 3.3 0.00052136 0 0.00052128 0 0.00052138 3.3 0.0005213 3.3 0.0005214 0 0.00052132 0 0.00052142 3.3 0.00052134 3.3 0.00052144 0 0.00052136 0 0.00052146 3.3 0.00052138 3.3 0.00052148 0 0.0005214 0 0.0005214999999999999 3.3 0.0005214200000000001 3.3 0.00052152 0 0.0005214400000000001 0 0.00052154 3.3 0.0005214600000000001 3.3 0.00052156 0 0.0005214800000000001 0 0.00052158 3.3 0.0005215 3.3 0.0005216 0 0.00052152 0 0.00052162 3.3 0.00052154 3.3 0.00052164 0 0.00052156 0 0.00052166 3.3 0.00052158 3.3 0.00052168 0 0.0005216 0 0.0005216999999999999 3.3 0.0005216200000000001 3.3 0.00052172 0 0.0005216400000000001 0 0.00052174 3.3 0.0005216600000000001 3.3 0.00052176 0 0.0005216800000000001 0 0.00052178 3.3 0.0005217 3.3 0.0005218 0 0.00052172 0 0.00052182 3.3 0.00052174 3.3 0.00052184 0 0.00052176 0 0.00052186 3.3 0.00052178 3.3 0.00052188 0 0.0005218 0 0.0005219 3.3 0.00052182 3.3 0.0005219199999999999 0 0.0005218400000000001 0 0.00052194 3.3 0.0005218600000000001 3.3 0.00052196 0 0.0005218800000000001 0 0.00052198 3.3 0.0005219000000000001 3.3 0.000522 0 0.00052192 0 0.00052202 3.3 0.00052194 3.3 0.00052204 0 0.00052196 0 0.00052206 3.3 0.00052198 3.3 0.00052208 0 0.000522 0 0.0005221 3.3 0.00052202 3.3 0.0005221199999999999 0 0.0005220400000000001 0 0.00052214 3.3 0.0005220600000000001 3.3 0.00052216 0 0.0005220800000000001 0 0.00052218 3.3 0.0005221000000000001 3.3 0.0005222 0 0.00052212 0 0.00052222 3.3 0.00052214 3.3 0.00052224 0 0.00052216 0 0.00052226 3.3 0.00052218 3.3 0.00052228 0 0.0005222 0 0.0005223 3.3 0.00052222 3.3 0.0005223199999999999 0 0.00052224 0 0.0005223399999999999 3.3 0.0005222600000000001 3.3 0.00052236 0 0.0005222800000000001 0 0.00052238 3.3 0.0005223000000000001 3.3 0.0005224 0 0.00052232 0 0.00052242 3.3 0.00052234 3.3 0.00052244 0 0.00052236 0 0.00052246 3.3 0.00052238 3.3 0.00052248 0 0.0005224 0 0.0005225 3.3 0.00052242 3.3 0.00052252 0 0.00052244 0 0.0005225399999999999 3.3 0.0005224600000000001 3.3 0.00052256 0 0.0005224800000000001 0 0.00052258 3.3 0.0005225000000000001 3.3 0.0005226 0 0.0005225200000000001 0 0.00052262 3.3 0.00052254 3.3 0.00052264 0 0.00052256 0 0.00052266 3.3 0.00052258 3.3 0.00052268 0 0.0005226 0 0.0005227 3.3 0.00052262 3.3 0.00052272 0 0.00052264 0 0.0005227399999999999 3.3 0.0005226600000000001 3.3 0.00052276 0 0.0005226800000000001 0 0.00052278 3.3 0.0005227000000000001 3.3 0.0005228 0 0.0005227200000000001 0 0.00052282 3.3 0.00052274 3.3 0.00052284 0 0.00052276 0 0.00052286 3.3 0.00052278 3.3 0.00052288 0 0.0005228 0 0.0005229 3.3 0.00052282 3.3 0.00052292 0 0.00052284 0 0.00052294 3.3 0.00052286 3.3 0.0005229599999999999 0 0.0005228800000000001 0 0.00052298 3.3 0.0005229000000000001 3.3 0.000523 0 0.0005229200000000001 0 0.00052302 3.3 0.0005229400000000001 3.3 0.00052304 0 0.00052296 0 0.00052306 3.3 0.00052298 3.3 0.00052308 0 0.000523 0 0.0005231 3.3 0.00052302 3.3 0.00052312 0 0.00052304 0 0.00052314 3.3 0.00052306 3.3 0.0005231599999999999 0 0.0005230800000000001 0 0.00052318 3.3 0.0005231000000000001 3.3 0.0005232 0 0.0005231200000000001 0 0.00052322 3.3 0.0005231400000000001 3.3 0.00052324 0 0.00052316 0 0.00052326 3.3 0.00052318 3.3 0.00052328 0 0.0005232 0 0.0005233 3.3 0.00052322 3.3 0.00052332 0 0.00052324 0 0.00052334 3.3 0.00052326 3.3 0.00052336 0 0.00052328 0 0.0005233799999999999 3.3 0.0005233000000000001 3.3 0.0005234 0 0.0005233200000000001 0 0.00052342 3.3 0.0005233400000000001 3.3 0.00052344 0 0.0005233600000000001 0 0.00052346 3.3 0.00052338 3.3 0.00052348 0 0.0005234 0 0.0005235 3.3 0.00052342 3.3 0.00052352 0 0.00052344 0 0.00052354 3.3 0.00052346 3.3 0.00052356 0 0.00052348 0 0.0005235799999999999 3.3 0.0005235000000000001 3.3 0.0005236 0 0.0005235200000000001 0 0.00052362 3.3 0.0005235400000000001 3.3 0.00052364 0 0.0005235600000000001 0 0.00052366 3.3 0.00052358 3.3 0.00052368 0 0.0005236 0 0.0005237 3.3 0.00052362 3.3 0.00052372 0 0.00052364 0 0.00052374 3.3 0.00052366 3.3 0.00052376 0 0.00052368 0 0.00052378 3.3 0.0005237 3.3 0.0005237999999999999 0 0.0005237200000000001 0 0.00052382 3.3 0.0005237400000000001 3.3 0.00052384 0 0.0005237600000000001 0 0.00052386 3.3 0.0005237800000000001 3.3 0.00052388 0 0.0005238 0 0.0005239 3.3 0.00052382 3.3 0.00052392 0 0.00052384 0 0.00052394 3.3 0.00052386 3.3 0.00052396 0 0.00052388 0 0.00052398 3.3 0.0005239 3.3 0.0005239999999999999 0 0.0005239200000000001 0 0.00052402 3.3 0.0005239400000000001 3.3 0.00052404 0 0.0005239600000000001 0 0.00052406 3.3 0.0005239800000000001 3.3 0.00052408 0 0.000524 0 0.0005241 3.3 0.00052402 3.3 0.00052412 0 0.00052404 0 0.00052414 3.3 0.00052406 3.3 0.00052416 0 0.00052408 0 0.00052418 3.3 0.0005241 3.3 0.0005242 0 0.00052412 0 0.0005242199999999999 3.3 0.0005241400000000001 3.3 0.00052424 0 0.0005241600000000001 0 0.00052426 3.3 0.0005241800000000001 3.3 0.00052428 0 0.0005242000000000001 0 0.0005243 3.3 0.00052422 3.3 0.00052432 0 0.00052424 0 0.00052434 3.3 0.00052426 3.3 0.00052436 0 0.00052428 0 0.00052438 3.3 0.0005243 3.3 0.0005244 0 0.00052432 0 0.0005244199999999999 3.3 0.0005243400000000001 3.3 0.00052444 0 0.0005243600000000001 0 0.00052446 3.3 0.0005243800000000001 3.3 0.00052448 0 0.0005244000000000001 0 0.0005245 3.3 0.00052442 3.3 0.00052452 0 0.00052444 0 0.00052454 3.3 0.00052446 3.3 0.00052456 0 0.00052448 0 0.00052458 3.3 0.0005245 3.3 0.0005246 0 0.00052452 0 0.00052462 3.3 0.00052454 3.3 0.0005246399999999999 0 0.0005245600000000001 0 0.00052466 3.3 0.0005245800000000001 3.3 0.00052468 0 0.0005246000000000001 0 0.0005247 3.3 0.0005246200000000001 3.3 0.00052472 0 0.00052464 0 0.00052474 3.3 0.00052466 3.3 0.00052476 0 0.00052468 0 0.00052478 3.3 0.0005247 3.3 0.0005248 0 0.00052472 0 0.00052482 3.3 0.00052474 3.3 0.0005248399999999999 0 0.0005247600000000001 0 0.00052486 3.3 0.0005247800000000001 3.3 0.00052488 0 0.0005248000000000001 0 0.0005249 3.3 0.0005248200000000001 3.3 0.00052492 0 0.00052484 0 0.00052494 3.3 0.00052486 3.3 0.00052496 0 0.00052488 0 0.00052498 3.3 0.0005249 3.3 0.000525 0 0.00052492 0 0.00052502 3.3 0.00052494 3.3 0.00052504 0 0.00052496 0 0.0005250599999999999 3.3 0.0005249800000000001 3.3 0.00052508 0 0.0005250000000000001 0 0.0005251 3.3 0.0005250200000000001 3.3 0.00052512 0 0.0005250400000000001 0 0.00052514 3.3 0.00052506 3.3 0.00052516 0 0.00052508 0 0.00052518 3.3 0.0005251 3.3 0.0005252 0 0.00052512 0 0.00052522 3.3 0.00052514 3.3 0.00052524 0 0.00052516 0 0.0005252599999999999 3.3 0.0005251800000000001 3.3 0.00052528 0 0.0005252000000000001 0 0.0005253 3.3 0.0005252200000000001 3.3 0.00052532 0 0.0005252400000000001 0 0.00052534 3.3 0.00052526 3.3 0.00052536 0 0.00052528 0 0.00052538 3.3 0.0005253 3.3 0.0005254 0 0.00052532 0 0.00052542 3.3 0.00052534 3.3 0.00052544 0 0.00052536 0 0.00052546 3.3 0.00052538 3.3 0.0005254799999999999 0 0.0005254000000000001 0 0.0005255 3.3 0.0005254200000000001 3.3 0.00052552 0 0.0005254400000000001 0 0.00052554 3.3 0.0005254600000000001 3.3 0.00052556 0 0.00052548 0 0.00052558 3.3 0.0005255 3.3 0.0005256 0 0.00052552 0 0.00052562 3.3 0.00052554 3.3 0.00052564 0 0.00052556 0 0.00052566 3.3 0.00052558 3.3 0.0005256799999999999 0 0.0005256000000000001 0 0.0005257 3.3 0.0005256200000000001 3.3 0.00052572 0 0.0005256400000000001 0 0.00052574 3.3 0.0005256600000000001 3.3 0.00052576 0 0.00052568 0 0.00052578 3.3 0.0005257 3.3 0.0005258 0 0.00052572 0 0.00052582 3.3 0.00052574 3.3 0.00052584 0 0.00052576 0 0.00052586 3.3 0.00052578 3.3 0.0005258799999999999 0 0.0005258 0 0.0005258999999999999 3.3 0.0005258200000000001 3.3 0.00052592 0 0.0005258400000000001 0 0.00052594 3.3 0.0005258600000000001 3.3 0.00052596 0 0.00052588 0 0.00052598 3.3 0.0005259 3.3 0.000526 0 0.00052592 0 0.00052602 3.3 0.00052594 3.3 0.00052604 0 0.00052596 0 0.00052606 3.3 0.00052598 3.3 0.00052608 0 0.000526 0 0.0005260999999999999 3.3 0.0005260200000000001 3.3 0.00052612 0 0.0005260400000000001 0 0.00052614 3.3 0.0005260600000000001 3.3 0.00052616 0 0.0005260800000000001 0 0.00052618 3.3 0.0005261 3.3 0.0005262 0 0.00052612 0 0.00052622 3.3 0.00052614 3.3 0.00052624 0 0.00052616 0 0.00052626 3.3 0.00052618 3.3 0.00052628 0 0.0005262 0 0.0005262999999999999 3.3 0.0005262200000000001 3.3 0.00052632 0 0.0005262400000000001 0 0.00052634 3.3 0.0005262600000000001 3.3 0.00052636 0 0.0005262800000000001 0 0.00052638 3.3 0.0005263 3.3 0.0005264 0 0.00052632 0 0.00052642 3.3 0.00052634 3.3 0.00052644 0 0.00052636 0 0.00052646 3.3 0.00052638 3.3 0.00052648 0 0.0005264 0 0.0005265 3.3 0.00052642 3.3 0.0005265199999999999 0 0.0005264400000000001 0 0.00052654 3.3 0.0005264600000000001 3.3 0.00052656 0 0.0005264800000000001 0 0.00052658 3.3 0.0005265000000000001 3.3 0.0005266 0 0.00052652 0 0.00052662 3.3 0.00052654 3.3 0.00052664 0 0.00052656 0 0.00052666 3.3 0.00052658 3.3 0.00052668 0 0.0005266 0 0.0005267 3.3 0.00052662 3.3 0.0005267199999999999 0 0.0005266400000000001 0 0.00052674 3.3 0.0005266600000000001 3.3 0.00052676 0 0.0005266800000000001 0 0.00052678 3.3 0.0005267000000000001 3.3 0.0005268 0 0.00052672 0 0.00052682 3.3 0.00052674 3.3 0.00052684 0 0.00052676 0 0.00052686 3.3 0.00052678 3.3 0.00052688 0 0.0005268 0 0.0005269 3.3 0.00052682 3.3 0.00052692 0 0.00052684 0 0.0005269399999999999 3.3 0.0005268600000000001 3.3 0.00052696 0 0.0005268800000000001 0 0.00052698 3.3 0.0005269000000000001 3.3 0.000527 0 0.0005269200000000001 0 0.00052702 3.3 0.00052694 3.3 0.00052704 0 0.00052696 0 0.00052706 3.3 0.00052698 3.3 0.00052708 0 0.000527 0 0.0005271 3.3 0.00052702 3.3 0.00052712 0 0.00052704 0 0.0005271399999999999 3.3 0.0005270600000000001 3.3 0.00052716 0 0.0005270800000000001 0 0.00052718 3.3 0.0005271000000000001 3.3 0.0005272 0 0.0005271200000000001 0 0.00052722 3.3 0.00052714 3.3 0.00052724 0 0.00052716 0 0.00052726 3.3 0.00052718 3.3 0.00052728 0 0.0005272 0 0.0005273 3.3 0.00052722 3.3 0.00052732 0 0.00052724 0 0.00052734 3.3 0.00052726 3.3 0.0005273599999999999 0 0.0005272800000000001 0 0.00052738 3.3 0.0005273000000000001 3.3 0.0005274 0 0.0005273200000000001 0 0.00052742 3.3 0.0005273400000000001 3.3 0.00052744 0 0.00052736 0 0.00052746 3.3 0.00052738 3.3 0.00052748 0 0.0005274 0 0.0005275 3.3 0.00052742 3.3 0.00052752 0 0.00052744 0 0.00052754 3.3 0.00052746 3.3 0.0005275599999999999 0 0.0005274800000000001 0 0.00052758 3.3 0.0005275000000000001 3.3 0.0005276 0 0.0005275200000000001 0 0.00052762 3.3 0.0005275400000000001 3.3 0.00052764 0 0.00052756 0 0.00052766 3.3 0.00052758 3.3 0.00052768 0 0.0005276 0 0.0005277 3.3 0.00052762 3.3 0.00052772 0 0.00052764 0 0.00052774 3.3 0.00052766 3.3 0.00052776 0 0.00052768 0 0.0005277799999999999 3.3 0.0005277000000000001 3.3 0.0005278 0 0.0005277200000000001 0 0.00052782 3.3 0.0005277400000000001 3.3 0.00052784 0 0.0005277600000000001 0 0.00052786 3.3 0.00052778 3.3 0.00052788 0 0.0005278 0 0.0005279 3.3 0.00052782 3.3 0.00052792 0 0.00052784 0 0.00052794 3.3 0.00052786 3.3 0.00052796 0 0.00052788 0 0.0005279799999999999 3.3 0.0005279000000000001 3.3 0.000528 0 0.0005279200000000001 0 0.00052802 3.3 0.0005279400000000001 3.3 0.00052804 0 0.0005279600000000001 0 0.00052806 3.3 0.00052798 3.3 0.00052808 0 0.000528 0 0.0005281 3.3 0.00052802 3.3 0.00052812 0 0.00052804 0 0.00052814 3.3 0.00052806 3.3 0.00052816 0 0.00052808 0 0.00052818 3.3 0.0005281 3.3 0.0005281999999999999 0 0.0005281200000000001 0 0.00052822 3.3 0.0005281400000000001 3.3 0.00052824 0 0.0005281600000000001 0 0.00052826 3.3 0.0005281800000000001 3.3 0.00052828 0 0.0005282 0 0.0005283 3.3 0.00052822 3.3 0.00052832 0 0.00052824 0 0.00052834 3.3 0.00052826 3.3 0.00052836 0 0.00052828 0 0.00052838 3.3 0.0005283 3.3 0.0005283999999999999 0 0.0005283200000000001 0 0.00052842 3.3 0.0005283400000000001 3.3 0.00052844 0 0.0005283600000000001 0 0.00052846 3.3 0.0005283800000000001 3.3 0.00052848 0 0.0005284 0 0.0005285 3.3 0.00052842 3.3 0.00052852 0 0.00052844 0 0.00052854 3.3 0.00052846 3.3 0.00052856 0 0.00052848 0 0.00052858 3.3 0.0005285 3.3 0.0005286 0 0.00052852 0 0.0005286199999999999 3.3 0.0005285400000000001 3.3 0.00052864 0 0.0005285600000000001 0 0.00052866 3.3 0.0005285800000000001 3.3 0.00052868 0 0.0005286000000000001 0 0.0005287 3.3 0.00052862 3.3 0.00052872 0 0.00052864 0 0.00052874 3.3 0.00052866 3.3 0.00052876 0 0.00052868 0 0.00052878 3.3 0.0005287 3.3 0.0005288 0 0.00052872 0 0.0005288199999999999 3.3 0.0005287400000000001 3.3 0.00052884 0 0.0005287600000000001 0 0.00052886 3.3 0.0005287800000000001 3.3 0.00052888 0 0.0005288000000000001 0 0.0005289 3.3 0.00052882 3.3 0.00052892 0 0.00052884 0 0.00052894 3.3 0.00052886 3.3 0.00052896 0 0.00052888 0 0.00052898 3.3 0.0005289 3.3 0.000529 0 0.00052892 0 0.00052902 3.3 0.00052894 3.3 0.0005290399999999999 0 0.0005289600000000001 0 0.00052906 3.3 0.0005289800000000001 3.3 0.00052908 0 0.0005290000000000001 0 0.0005291 3.3 0.0005290200000000001 3.3 0.00052912 0 0.00052904 0 0.00052914 3.3 0.00052906 3.3 0.00052916 0 0.00052908 0 0.00052918 3.3 0.0005291 3.3 0.0005292 0 0.00052912 0 0.00052922 3.3 0.00052914 3.3 0.0005292399999999999 0 0.0005291600000000001 0 0.00052926 3.3 0.0005291800000000001 3.3 0.00052928 0 0.0005292000000000001 0 0.0005293 3.3 0.0005292200000000001 3.3 0.00052932 0 0.00052924 0 0.00052934 3.3 0.00052926 3.3 0.00052936 0 0.00052928 0 0.00052938 3.3 0.0005293 3.3 0.0005294 0 0.00052932 0 0.00052942 3.3 0.00052934 3.3 0.0005294399999999999 0 0.0005293600000000001 0 0.00052946 3.3 0.0005293800000000001 3.3 0.00052948 0 0.0005294000000000001 0 0.0005295 3.3 0.0005294200000000001 3.3 0.00052952 0 0.00052944 0 0.00052954 3.3 0.00052946 3.3 0.00052956 0 0.00052948 0 0.00052958 3.3 0.0005295 3.3 0.0005296 0 0.00052952 0 0.00052962 3.3 0.00052954 3.3 0.00052964 0 0.00052956 0 0.0005296599999999999 3.3 0.0005295800000000001 3.3 0.00052968 0 0.0005296000000000001 0 0.0005297 3.3 0.0005296200000000001 3.3 0.00052972 0 0.0005296400000000001 0 0.00052974 3.3 0.00052966 3.3 0.00052976 0 0.00052968 0 0.00052978 3.3 0.0005297 3.3 0.0005298 0 0.00052972 0 0.00052982 3.3 0.00052974 3.3 0.00052984 0 0.00052976 0 0.0005298599999999999 3.3 0.0005297800000000001 3.3 0.00052988 0 0.0005298000000000001 0 0.0005299 3.3 0.0005298200000000001 3.3 0.00052992 0 0.0005298400000000001 0 0.00052994 3.3 0.00052986 3.3 0.00052996 0 0.00052988 0 0.00052998 3.3 0.0005299 3.3 0.00053 0 0.00052992 0 0.00053002 3.3 0.00052994 3.3 0.00053004 0 0.00052996 0 0.00053006 3.3 0.00052998 3.3 0.0005300799999999999 0 0.0005300000000000001 0 0.0005301 3.3 0.0005300200000000001 3.3 0.00053012 0 0.0005300400000000001 0 0.00053014 3.3 0.0005300600000000001 3.3 0.00053016 0 0.00053008 0 0.00053018 3.3 0.0005301 3.3 0.0005302 0 0.00053012 0 0.00053022 3.3 0.00053014 3.3 0.00053024 0 0.00053016 0 0.00053026 3.3 0.00053018 3.3 0.0005302799999999999 0 0.0005302000000000001 0 0.0005303 3.3 0.0005302200000000001 3.3 0.00053032 0 0.0005302400000000001 0 0.00053034 3.3 0.0005302600000000001 3.3 0.00053036 0 0.00053028 0 0.00053038 3.3 0.0005303 3.3 0.0005304 0 0.00053032 0 0.00053042 3.3 0.00053034 3.3 0.00053044 0 0.00053036 0 0.00053046 3.3 0.00053038 3.3 0.00053048 0 0.0005304 0 0.0005304999999999999 3.3 0.0005304200000000001 3.3 0.00053052 0 0.0005304400000000001 0 0.00053054 3.3 0.0005304600000000001 3.3 0.00053056 0 0.0005304800000000001 0 0.00053058 3.3 0.0005305 3.3 0.0005306 0 0.00053052 0 0.00053062 3.3 0.00053054 3.3 0.00053064 0 0.00053056 0 0.00053066 3.3 0.00053058 3.3 0.00053068 0 0.0005306 0 0.0005306999999999999 3.3 0.0005306200000000001 3.3 0.00053072 0 0.0005306400000000001 0 0.00053074 3.3 0.0005306600000000001 3.3 0.00053076 0 0.0005306800000000001 0 0.00053078 3.3 0.0005307 3.3 0.0005308 0 0.00053072 0 0.00053082 3.3 0.00053074 3.3 0.00053084 0 0.00053076 0 0.00053086 3.3 0.00053078 3.3 0.00053088 0 0.0005308 0 0.0005309 3.3 0.00053082 3.3 0.0005309199999999999 0 0.0005308400000000001 0 0.00053094 3.3 0.0005308600000000001 3.3 0.00053096 0 0.0005308800000000001 0 0.00053098 3.3 0.0005309000000000001 3.3 0.000531 0 0.00053092 0 0.00053102 3.3 0.00053094 3.3 0.00053104 0 0.00053096 0 0.00053106 3.3 0.00053098 3.3 0.00053108 0 0.000531 0 0.0005311 3.3 0.00053102 3.3 0.0005311199999999999 0 0.0005310400000000001 0 0.00053114 3.3 0.0005310600000000001 3.3 0.00053116 0 0.0005310800000000001 0 0.00053118 3.3 0.0005311000000000001 3.3 0.0005312 0 0.00053112 0 0.00053122 3.3 0.00053114 3.3 0.00053124 0 0.00053116 0 0.00053126 3.3 0.00053118 3.3 0.00053128 0 0.0005312 0 0.0005313 3.3 0.00053122 3.3 0.00053132 0 0.00053124 0 0.0005313399999999999 3.3 0.0005312600000000001 3.3 0.00053136 0 0.0005312800000000001 0 0.00053138 3.3 0.0005313000000000001 3.3 0.0005314 0 0.0005313200000000001 0 0.00053142 3.3 0.00053134 3.3 0.00053144 0 0.00053136 0 0.00053146 3.3 0.00053138 3.3 0.00053148 0 0.0005314 0 0.0005315 3.3 0.00053142 3.3 0.00053152 0 0.00053144 0 0.0005315399999999999 3.3 0.0005314600000000001 3.3 0.00053156 0 0.0005314800000000001 0 0.00053158 3.3 0.0005315000000000001 3.3 0.0005316 0 0.0005315200000000001 0 0.00053162 3.3 0.00053154 3.3 0.00053164 0 0.00053156 0 0.00053166 3.3 0.00053158 3.3 0.00053168 0 0.0005316 0 0.0005317 3.3 0.00053162 3.3 0.00053172 0 0.00053164 0 0.00053174 3.3 0.00053166 3.3 0.0005317599999999999 0 0.0005316800000000001 0 0.00053178 3.3 0.0005317000000000001 3.3 0.0005318 0 0.0005317200000000001 0 0.00053182 3.3 0.0005317400000000001 3.3 0.00053184 0 0.00053176 0 0.00053186 3.3 0.00053178 3.3 0.00053188 0 0.0005318 0 0.0005319 3.3 0.00053182 3.3 0.00053192 0 0.00053184 0 0.00053194 3.3 0.00053186 3.3 0.0005319599999999999 0 0.0005318800000000001 0 0.00053198 3.3 0.0005319000000000001 3.3 0.000532 0 0.0005319200000000001 0 0.00053202 3.3 0.0005319400000000001 3.3 0.00053204 0 0.00053196 0 0.00053206 3.3 0.00053198 3.3 0.00053208 0 0.000532 0 0.0005321 3.3 0.00053202 3.3 0.00053212 0 0.00053204 0 0.00053214 3.3 0.00053206 3.3 0.00053216 0 0.00053208 0 0.0005321799999999999 3.3 0.0005321000000000001 3.3 0.0005322 0 0.0005321200000000001 0 0.00053222 3.3 0.0005321400000000001 3.3 0.00053224 0 0.0005321600000000001 0 0.00053226 3.3 0.00053218 3.3 0.00053228 0 0.0005322 0 0.0005323 3.3 0.00053222 3.3 0.00053232 0 0.00053224 0 0.00053234 3.3 0.00053226 3.3 0.00053236 0 0.00053228 0 0.0005323799999999999 3.3 0.0005323000000000001 3.3 0.0005324 0 0.0005323200000000001 0 0.00053242 3.3 0.0005323400000000001 3.3 0.00053244 0 0.0005323600000000001 0 0.00053246 3.3 0.00053238 3.3 0.00053248 0 0.0005324 0 0.0005325 3.3 0.00053242 3.3 0.00053252 0 0.00053244 0 0.00053254 3.3 0.00053246 3.3 0.00053256 0 0.00053248 0 0.00053258 3.3 0.0005325 3.3 0.0005325999999999999 0 0.0005325200000000001 0 0.00053262 3.3 0.0005325400000000001 3.3 0.00053264 0 0.0005325600000000001 0 0.00053266 3.3 0.0005325800000000001 3.3 0.00053268 0 0.0005326 0 0.0005327 3.3 0.00053262 3.3 0.00053272 0 0.00053264 0 0.00053274 3.3 0.00053266 3.3 0.00053276 0 0.00053268 0 0.00053278 3.3 0.0005327 3.3 0.0005327999999999999 0 0.0005327200000000001 0 0.00053282 3.3 0.0005327400000000001 3.3 0.00053284 0 0.0005327600000000001 0 0.00053286 3.3 0.0005327800000000001 3.3 0.00053288 0 0.0005328 0 0.0005329 3.3 0.00053282 3.3 0.00053292 0 0.00053284 0 0.00053294 3.3 0.00053286 3.3 0.00053296 0 0.00053288 0 0.00053298 3.3 0.0005329 3.3 0.0005329999999999999 0 0.0005329200000000001 0 0.00053302 3.3 0.0005329400000000001 3.3 0.00053304 0 0.0005329600000000001 0 0.00053306 3.3 0.0005329800000000001 3.3 0.00053308 0 0.000533 0 0.0005331 3.3 0.00053302 3.3 0.00053312 0 0.00053304 0 0.00053314 3.3 0.00053306 3.3 0.00053316 0 0.00053308 0 0.00053318 3.3 0.0005331 3.3 0.0005332 0 0.00053312 0 0.0005332199999999999 3.3 0.0005331400000000001 3.3 0.00053324 0 0.0005331600000000001 0 0.00053326 3.3 0.0005331800000000001 3.3 0.00053328 0 0.0005332000000000001 0 0.0005333 3.3 0.00053322 3.3 0.00053332 0 0.00053324 0 0.00053334 3.3 0.00053326 3.3 0.00053336 0 0.00053328 0 0.00053338 3.3 0.0005333 3.3 0.0005334 0 0.00053332 0 0.0005334199999999999 3.3 0.0005333400000000001 3.3 0.00053344 0 0.0005333600000000001 0 0.00053346 3.3 0.0005333800000000001 3.3 0.00053348 0 0.0005334000000000001 0 0.0005335 3.3 0.00053342 3.3 0.00053352 0 0.00053344 0 0.00053354 3.3 0.00053346 3.3 0.00053356 0 0.00053348 0 0.00053358 3.3 0.0005335 3.3 0.0005336 0 0.00053352 0 0.00053362 3.3 0.00053354 3.3 0.0005336399999999999 0 0.0005335600000000001 0 0.00053366 3.3 0.0005335800000000001 3.3 0.00053368 0 0.0005336000000000001 0 0.0005337 3.3 0.0005336200000000001 3.3 0.00053372 0 0.00053364 0 0.00053374 3.3 0.00053366 3.3 0.00053376 0 0.00053368 0 0.00053378 3.3 0.0005337 3.3 0.0005338 0 0.00053372 0 0.00053382 3.3 0.00053374 3.3 0.0005338399999999999 0 0.0005337600000000001 0 0.00053386 3.3 0.0005337800000000001 3.3 0.00053388 0 0.0005338000000000001 0 0.0005339 3.3 0.0005338200000000001 3.3 0.00053392 0 0.00053384 0 0.00053394 3.3 0.00053386 3.3 0.00053396 0 0.00053388 0 0.00053398 3.3 0.0005339 3.3 0.000534 0 0.00053392 0 0.00053402 3.3 0.00053394 3.3 0.00053404 0 0.00053396 0 0.0005340599999999999 3.3 0.0005339800000000001 3.3 0.00053408 0 0.0005340000000000001 0 0.0005341 3.3 0.0005340200000000001 3.3 0.00053412 0 0.0005340400000000001 0 0.00053414 3.3 0.00053406 3.3 0.00053416 0 0.00053408 0 0.00053418 3.3 0.0005341 3.3 0.0005342 0 0.00053412 0 0.00053422 3.3 0.00053414 3.3 0.00053424 0 0.00053416 0 0.0005342599999999999 3.3 0.0005341800000000001 3.3 0.00053428 0 0.0005342000000000001 0 0.0005343 3.3 0.0005342200000000001 3.3 0.00053432 0 0.0005342400000000001 0 0.00053434 3.3 0.00053426 3.3 0.00053436 0 0.00053428 0 0.00053438 3.3 0.0005343 3.3 0.0005344 0 0.00053432 0 0.00053442 3.3 0.00053434 3.3 0.00053444 0 0.00053436 0 0.00053446 3.3 0.00053438 3.3 0.0005344799999999999 0 0.0005344000000000001 0 0.0005345 3.3 0.0005344200000000001 3.3 0.00053452 0 0.0005344400000000001 0 0.00053454 3.3 0.0005344600000000001 3.3 0.00053456 0 0.00053448 0 0.00053458 3.3 0.0005345 3.3 0.0005346 0 0.00053452 0 0.00053462 3.3 0.00053454 3.3 0.00053464 0 0.00053456 0 0.00053466 3.3 0.00053458 3.3 0.0005346799999999999 0 0.0005346000000000001 0 0.0005347 3.3 0.0005346200000000001 3.3 0.00053472 0 0.0005346400000000001 0 0.00053474 3.3 0.0005346600000000001 3.3 0.00053476 0 0.00053468 0 0.00053478 3.3 0.0005347 3.3 0.0005348 0 0.00053472 0 0.00053482 3.3 0.00053474 3.3 0.00053484 0 0.00053476 0 0.00053486 3.3 0.00053478 3.3 0.00053488 0 0.0005348 0 0.0005348999999999999 3.3 0.0005348200000000001 3.3 0.00053492 0 0.0005348400000000001 0 0.00053494 3.3 0.0005348600000000001 3.3 0.00053496 0 0.0005348800000000001 0 0.00053498 3.3 0.0005349 3.3 0.000535 0 0.00053492 0 0.00053502 3.3 0.00053494 3.3 0.00053504 0 0.00053496 0 0.00053506 3.3 0.00053498 3.3 0.00053508 0 0.000535 0 0.0005350999999999999 3.3 0.0005350200000000001 3.3 0.00053512 0 0.0005350400000000001 0 0.00053514 3.3 0.0005350600000000001 3.3 0.00053516 0 0.0005350800000000001 0 0.00053518 3.3 0.0005351 3.3 0.0005352 0 0.00053512 0 0.00053522 3.3 0.00053514 3.3 0.00053524 0 0.00053516 0 0.00053526 3.3 0.00053518 3.3 0.00053528 0 0.0005352 0 0.0005353 3.3 0.00053522 3.3 0.0005353199999999999 0 0.0005352400000000001 0 0.00053534 3.3 0.0005352600000000001 3.3 0.00053536 0 0.0005352800000000001 0 0.00053538 3.3 0.0005353000000000001 3.3 0.0005354 0 0.00053532 0 0.00053542 3.3 0.00053534 3.3 0.00053544 0 0.00053536 0 0.00053546 3.3 0.00053538 3.3 0.00053548 0 0.0005354 0 0.0005355 3.3 0.00053542 3.3 0.0005355199999999999 0 0.0005354400000000001 0 0.00053554 3.3 0.0005354600000000001 3.3 0.00053556 0 0.0005354800000000001 0 0.00053558 3.3 0.0005355000000000001 3.3 0.0005356 0 0.00053552 0 0.00053562 3.3 0.00053554 3.3 0.00053564 0 0.00053556 0 0.00053566 3.3 0.00053558 3.3 0.00053568 0 0.0005356 0 0.0005357 3.3 0.00053562 3.3 0.00053572 0 0.00053564 0 0.0005357399999999999 3.3 0.0005356600000000001 3.3 0.00053576 0 0.0005356800000000001 0 0.00053578 3.3 0.0005357000000000001 3.3 0.0005358 0 0.0005357200000000001 0 0.00053582 3.3 0.00053574 3.3 0.00053584 0 0.00053576 0 0.00053586 3.3 0.00053578 3.3 0.00053588 0 0.0005358 0 0.0005359 3.3 0.00053582 3.3 0.00053592 0 0.00053584 0 0.0005359399999999999 3.3 0.0005358600000000001 3.3 0.00053596 0 0.0005358800000000001 0 0.00053598 3.3 0.0005359000000000001 3.3 0.000536 0 0.0005359200000000001 0 0.00053602 3.3 0.00053594 3.3 0.00053604 0 0.00053596 0 0.00053606 3.3 0.00053598 3.3 0.00053608 0 0.000536 0 0.0005361 3.3 0.00053602 3.3 0.00053612 0 0.00053604 0 0.0005361399999999999 3.3 0.00053606 3.3 0.0005361599999999999 0 0.0005360800000000001 0 0.00053618 3.3 0.0005361000000000001 3.3 0.0005362 0 0.0005361200000000001 0 0.00053622 3.3 0.00053614 3.3 0.00053624 0 0.00053616 0 0.00053626 3.3 0.00053618 3.3 0.00053628 0 0.0005362 0 0.0005363 3.3 0.00053622 3.3 0.00053632 0 0.00053624 0 0.00053634 3.3 0.00053626 3.3 0.0005363599999999999 0 0.0005362800000000001 0 0.00053638 3.3 0.0005363000000000001 3.3 0.0005364 0 0.0005363200000000001 0 0.00053642 3.3 0.0005363400000000001 3.3 0.00053644 0 0.00053636 0 0.00053646 3.3 0.00053638 3.3 0.00053648 0 0.0005364 0 0.0005365 3.3 0.00053642 3.3 0.00053652 0 0.00053644 0 0.00053654 3.3 0.00053646 3.3 0.0005365599999999999 0 0.0005364800000000001 0 0.00053658 3.3 0.0005365000000000001 3.3 0.0005366 0 0.0005365200000000001 0 0.00053662 3.3 0.0005365400000000001 3.3 0.00053664 0 0.00053656 0 0.00053666 3.3 0.00053658 3.3 0.00053668 0 0.0005366 0 0.0005367 3.3 0.00053662 3.3 0.00053672 0 0.00053664 0 0.00053674 3.3 0.00053666 3.3 0.00053676 0 0.00053668 0 0.0005367799999999999 3.3 0.0005367000000000001 3.3 0.0005368 0 0.0005367200000000001 0 0.00053682 3.3 0.0005367400000000001 3.3 0.00053684 0 0.0005367600000000001 0 0.00053686 3.3 0.00053678 3.3 0.00053688 0 0.0005368 0 0.0005369 3.3 0.00053682 3.3 0.00053692 0 0.00053684 0 0.00053694 3.3 0.00053686 3.3 0.00053696 0 0.00053688 0 0.0005369799999999999 3.3 0.0005369000000000001 3.3 0.000537 0 0.0005369200000000001 0 0.00053702 3.3 0.0005369400000000001 3.3 0.00053704 0 0.0005369600000000001 0 0.00053706 3.3 0.00053698 3.3 0.00053708 0 0.000537 0 0.0005371 3.3 0.00053702 3.3 0.00053712 0 0.00053704 0 0.00053714 3.3 0.00053706 3.3 0.00053716 0 0.00053708 0 0.00053718 3.3 0.0005371 3.3 0.0005371999999999999 0 0.0005371200000000001 0 0.00053722 3.3 0.0005371400000000001 3.3 0.00053724 0 0.0005371600000000001 0 0.00053726 3.3 0.0005371800000000001 3.3 0.00053728 0 0.0005372 0 0.0005373 3.3 0.00053722 3.3 0.00053732 0 0.00053724 0 0.00053734 3.3 0.00053726 3.3 0.00053736 0 0.00053728 0 0.00053738 3.3 0.0005373 3.3 0.0005373999999999999 0 0.0005373200000000001 0 0.00053742 3.3 0.0005373400000000001 3.3 0.00053744 0 0.0005373600000000001 0 0.00053746 3.3 0.0005373800000000001 3.3 0.00053748 0 0.0005374 0 0.0005375 3.3 0.00053742 3.3 0.00053752 0 0.00053744 0 0.00053754 3.3 0.00053746 3.3 0.00053756 0 0.00053748 0 0.00053758 3.3 0.0005375 3.3 0.0005376 0 0.00053752 0 0.0005376199999999999 3.3 0.0005375400000000001 3.3 0.00053764 0 0.0005375600000000001 0 0.00053766 3.3 0.0005375800000000001 3.3 0.00053768 0 0.0005376000000000001 0 0.0005377 3.3 0.00053762 3.3 0.00053772 0 0.00053764 0 0.00053774 3.3 0.00053766 3.3 0.00053776 0 0.00053768 0 0.00053778 3.3 0.0005377 3.3 0.0005378 0 0.00053772 0 0.0005378199999999999 3.3 0.0005377400000000001 3.3 0.00053784 0 0.0005377600000000001 0 0.00053786 3.3 0.0005377800000000001 3.3 0.00053788 0 0.0005378000000000001 0 0.0005379 3.3 0.00053782 3.3 0.00053792 0 0.00053784 0 0.00053794 3.3 0.00053786 3.3 0.00053796 0 0.00053788 0 0.00053798 3.3 0.0005379 3.3 0.000538 0 0.00053792 0 0.00053802 3.3 0.00053794 3.3 0.0005380399999999999 0 0.0005379600000000001 0 0.00053806 3.3 0.0005379800000000001 3.3 0.00053808 0 0.0005380000000000001 0 0.0005381 3.3 0.0005380200000000001 3.3 0.00053812 0 0.00053804 0 0.00053814 3.3 0.00053806 3.3 0.00053816 0 0.00053808 0 0.00053818 3.3 0.0005381 3.3 0.0005382 0 0.00053812 0 0.00053822 3.3 0.00053814 3.3 0.0005382399999999999 0 0.0005381600000000001 0 0.00053826 3.3 0.0005381800000000001 3.3 0.00053828 0 0.0005382000000000001 0 0.0005383 3.3 0.0005382200000000001 3.3 0.00053832 0 0.00053824 0 0.00053834 3.3 0.00053826 3.3 0.00053836 0 0.00053828 0 0.00053838 3.3 0.0005383 3.3 0.0005384 0 0.00053832 0 0.00053842 3.3 0.00053834 3.3 0.00053844 0 0.00053836 0 0.0005384599999999999 3.3 0.0005383800000000001 3.3 0.00053848 0 0.0005384000000000001 0 0.0005385 3.3 0.0005384200000000001 3.3 0.00053852 0 0.0005384400000000001 0 0.00053854 3.3 0.00053846 3.3 0.00053856 0 0.00053848 0 0.00053858 3.3 0.0005385 3.3 0.0005386 0 0.00053852 0 0.00053862 3.3 0.00053854 3.3 0.00053864 0 0.00053856 0 0.0005386599999999999 3.3 0.0005385800000000001 3.3 0.00053868 0 0.0005386000000000001 0 0.0005387 3.3 0.0005386200000000001 3.3 0.00053872 0 0.0005386400000000001 0 0.00053874 3.3 0.00053866 3.3 0.00053876 0 0.00053868 0 0.00053878 3.3 0.0005387 3.3 0.0005388 0 0.00053872 0 0.00053882 3.3 0.00053874 3.3 0.00053884 0 0.00053876 0 0.00053886 3.3 0.00053878 3.3 0.0005388799999999999 0 0.0005388000000000001 0 0.0005389 3.3 0.0005388200000000001 3.3 0.00053892 0 0.0005388400000000001 0 0.00053894 3.3 0.0005388600000000001 3.3 0.00053896 0 0.00053888 0 0.00053898 3.3 0.0005389 3.3 0.000539 0 0.00053892 0 0.00053902 3.3 0.00053894 3.3 0.00053904 0 0.00053896 0 0.00053906 3.3 0.00053898 3.3 0.0005390799999999999 0 0.0005390000000000001 0 0.0005391 3.3 0.0005390200000000001 3.3 0.00053912 0 0.0005390400000000001 0 0.00053914 3.3 0.0005390600000000001 3.3 0.00053916 0 0.00053908 0 0.00053918 3.3 0.0005391 3.3 0.0005392 0 0.00053912 0 0.00053922 3.3 0.00053914 3.3 0.00053924 0 0.00053916 0 0.00053926 3.3 0.00053918 3.3 0.00053928 0 0.0005392 0 0.0005392999999999999 3.3 0.0005392200000000001 3.3 0.00053932 0 0.0005392400000000001 0 0.00053934 3.3 0.0005392600000000001 3.3 0.00053936 0 0.0005392800000000001 0 0.00053938 3.3 0.0005393 3.3 0.0005394 0 0.00053932 0 0.00053942 3.3 0.00053934 3.3 0.00053944 0 0.00053936 0 0.00053946 3.3 0.00053938 3.3 0.00053948 0 0.0005394 0 0.0005394999999999999 3.3 0.0005394200000000001 3.3 0.00053952 0 0.0005394400000000001 0 0.00053954 3.3 0.0005394600000000001 3.3 0.00053956 0 0.0005394800000000001 0 0.00053958 3.3 0.0005395 3.3 0.0005396 0 0.00053952 0 0.00053962 3.3 0.00053954 3.3 0.00053964 0 0.00053956 0 0.00053966 3.3 0.00053958 3.3 0.00053968 0 0.0005396 0 0.0005396999999999999 3.3 0.00053962 3.3 0.0005397199999999999 0 0.0005396400000000001 0 0.00053974 3.3 0.0005396600000000001 3.3 0.00053976 0 0.0005396800000000001 0 0.00053978 3.3 0.0005397 3.3 0.0005398 0 0.00053972 0 0.00053982 3.3 0.00053974 3.3 0.00053984 0 0.00053976 0 0.00053986 3.3 0.00053978 3.3 0.00053988 0 0.0005398 0 0.0005399 3.3 0.00053982 3.3 0.0005399199999999999 0 0.0005398400000000001 0 0.00053994 3.3 0.0005398600000000001 3.3 0.00053996 0 0.0005398800000000001 0 0.00053998 3.3 0.0005399000000000001 3.3 0.00054 0 0.00053992 0 0.00054002 3.3 0.00053994 3.3 0.00054004 0 0.00053996 0 0.00054006 3.3 0.00053998 3.3 0.00054008 0 0.00054 0 0.0005401 3.3 0.00054002 3.3 0.0005401199999999999 0 0.0005400400000000001 0 0.00054014 3.3 0.0005400600000000001 3.3 0.00054016 0 0.0005400800000000001 0 0.00054018 3.3 0.0005401000000000001 3.3 0.0005402 0 0.00054012 0 0.00054022 3.3 0.00054014 3.3 0.00054024 0 0.00054016 0 0.00054026 3.3 0.00054018 3.3 0.00054028 0 0.0005402 0 0.0005403 3.3 0.00054022 3.3 0.00054032 0 0.00054024 0 0.0005403399999999999 3.3 0.0005402600000000001 3.3 0.00054036 0 0.0005402800000000001 0 0.00054038 3.3 0.0005403000000000001 3.3 0.0005404 0 0.0005403200000000001 0 0.00054042 3.3 0.00054034 3.3 0.00054044 0 0.00054036 0 0.00054046 3.3 0.00054038 3.3 0.00054048 0 0.0005404 0 0.0005405 3.3 0.00054042 3.3 0.00054052 0 0.00054044 0 0.0005405399999999999 3.3 0.0005404600000000001 3.3 0.00054056 0 0.0005404800000000001 0 0.00054058 3.3 0.0005405000000000001 3.3 0.0005406 0 0.0005405200000000001 0 0.00054062 3.3 0.00054054 3.3 0.00054064 0 0.00054056 0 0.00054066 3.3 0.00054058 3.3 0.00054068 0 0.0005406 0 0.0005407 3.3 0.00054062 3.3 0.00054072 0 0.00054064 0 0.00054074 3.3 0.00054066 3.3 0.0005407599999999999 0 0.0005406800000000001 0 0.00054078 3.3 0.0005407000000000001 3.3 0.0005408 0 0.0005407200000000001 0 0.00054082 3.3 0.0005407400000000001 3.3 0.00054084 0 0.00054076 0 0.00054086 3.3 0.00054078 3.3 0.00054088 0 0.0005408 0 0.0005409 3.3 0.00054082 3.3 0.00054092 0 0.00054084 0 0.00054094 3.3 0.00054086 3.3 0.0005409599999999999 0 0.0005408800000000001 0 0.00054098 3.3 0.0005409000000000001 3.3 0.000541 0 0.0005409200000000001 0 0.00054102 3.3 0.0005409400000000001 3.3 0.00054104 0 0.00054096 0 0.00054106 3.3 0.00054098 3.3 0.00054108 0 0.000541 0 0.0005411 3.3 0.00054102 3.3 0.00054112 0 0.00054104 0 0.00054114 3.3 0.00054106 3.3 0.00054116 0 0.00054108 0 0.0005411799999999999 3.3 0.0005411000000000001 3.3 0.0005412 0 0.0005411200000000001 0 0.00054122 3.3 0.0005411400000000001 3.3 0.00054124 0 0.0005411600000000001 0 0.00054126 3.3 0.00054118 3.3 0.00054128 0 0.0005412 0 0.0005413 3.3 0.00054122 3.3 0.00054132 0 0.00054124 0 0.00054134 3.3 0.00054126 3.3 0.00054136 0 0.00054128 0 0.0005413799999999999 3.3 0.0005413000000000001 3.3 0.0005414 0 0.0005413200000000001 0 0.00054142 3.3 0.0005413400000000001 3.3 0.00054144 0 0.0005413600000000001 0 0.00054146 3.3 0.00054138 3.3 0.00054148 0 0.0005414 0 0.0005415 3.3 0.00054142 3.3 0.00054152 0 0.00054144 0 0.00054154 3.3 0.00054146 3.3 0.00054156 0 0.00054148 0 0.00054158 3.3 0.0005415 3.3 0.0005415999999999999 0 0.0005415200000000001 0 0.00054162 3.3 0.0005415400000000001 3.3 0.00054164 0 0.0005415600000000001 0 0.00054166 3.3 0.0005415800000000001 3.3 0.00054168 0 0.0005416 0 0.0005417 3.3 0.00054162 3.3 0.00054172 0 0.00054164 0 0.00054174 3.3 0.00054166 3.3 0.00054176 0 0.00054168 0 0.00054178 3.3 0.0005417 3.3 0.0005417999999999999 0 0.0005417200000000001 0 0.00054182 3.3 0.0005417400000000001 3.3 0.00054184 0 0.0005417600000000001 0 0.00054186 3.3 0.0005417800000000001 3.3 0.00054188 0 0.0005418 0 0.0005419 3.3 0.00054182 3.3 0.00054192 0 0.00054184 0 0.00054194 3.3 0.00054186 3.3 0.00054196 0 0.00054188 0 0.00054198 3.3 0.0005419 3.3 0.000542 0 0.00054192 0 0.0005420199999999999 3.3 0.0005419400000000001 3.3 0.00054204 0 0.0005419600000000001 0 0.00054206 3.3 0.0005419800000000001 3.3 0.00054208 0 0.0005420000000000001 0 0.0005421 3.3 0.00054202 3.3 0.00054212 0 0.00054204 0 0.00054214 3.3 0.00054206 3.3 0.00054216 0 0.00054208 0 0.00054218 3.3 0.0005421 3.3 0.0005422 0 0.00054212 0 0.0005422199999999999 3.3 0.0005421400000000001 3.3 0.00054224 0 0.0005421600000000001 0 0.00054226 3.3 0.0005421800000000001 3.3 0.00054228 0 0.0005422000000000001 0 0.0005423 3.3 0.00054222 3.3 0.00054232 0 0.00054224 0 0.00054234 3.3 0.00054226 3.3 0.00054236 0 0.00054228 0 0.00054238 3.3 0.0005423 3.3 0.0005424 0 0.00054232 0 0.00054242 3.3 0.00054234 3.3 0.0005424399999999999 0 0.0005423600000000001 0 0.00054246 3.3 0.0005423800000000001 3.3 0.00054248 0 0.0005424000000000001 0 0.0005425 3.3 0.0005424200000000001 3.3 0.00054252 0 0.00054244 0 0.00054254 3.3 0.00054246 3.3 0.00054256 0 0.00054248 0 0.00054258 3.3 0.0005425 3.3 0.0005426 0 0.00054252 0 0.00054262 3.3 0.00054254 3.3 0.0005426399999999999 0 0.0005425600000000001 0 0.00054266 3.3 0.0005425800000000001 3.3 0.00054268 0 0.0005426000000000001 0 0.0005427 3.3 0.0005426200000000001 3.3 0.00054272 0 0.00054264 0 0.00054274 3.3 0.00054266 3.3 0.00054276 0 0.00054268 0 0.00054278 3.3 0.0005427 3.3 0.0005428 0 0.00054272 0 0.00054282 3.3 0.00054274 3.3 0.00054284 0 0.00054276 0 0.0005428599999999999 3.3 0.0005427800000000001 3.3 0.00054288 0 0.0005428000000000001 0 0.0005429 3.3 0.0005428200000000001 3.3 0.00054292 0 0.0005428400000000001 0 0.00054294 3.3 0.00054286 3.3 0.00054296 0 0.00054288 0 0.00054298 3.3 0.0005429 3.3 0.000543 0 0.00054292 0 0.00054302 3.3 0.00054294 3.3 0.00054304 0 0.00054296 0 0.0005430599999999999 3.3 0.0005429800000000001 3.3 0.00054308 0 0.0005430000000000001 0 0.0005431 3.3 0.0005430200000000001 3.3 0.00054312 0 0.0005430400000000001 0 0.00054314 3.3 0.00054306 3.3 0.00054316 0 0.00054308 0 0.00054318 3.3 0.0005431 3.3 0.0005432 0 0.00054312 0 0.00054322 3.3 0.00054314 3.3 0.00054324 0 0.00054316 0 0.0005432599999999999 3.3 0.0005431800000000001 3.3 0.00054328 0 0.0005432000000000001 0 0.0005433 3.3 0.0005432200000000001 3.3 0.00054332 0 0.0005432400000000001 0 0.00054334 3.3 0.00054326 3.3 0.00054336 0 0.00054328 0 0.00054338 3.3 0.0005433 3.3 0.0005434 0 0.00054332 0 0.00054342 3.3 0.00054334 3.3 0.00054344 0 0.00054336 0 0.00054346 3.3 0.00054338 3.3 0.0005434799999999999 0 0.0005434000000000001 0 0.0005435 3.3 0.0005434200000000001 3.3 0.00054352 0 0.0005434400000000001 0 0.00054354 3.3 0.0005434600000000001 3.3 0.00054356 0 0.00054348 0 0.00054358 3.3 0.0005435 3.3 0.0005436 0 0.00054352 0 0.00054362 3.3 0.00054354 3.3 0.00054364 0 0.00054356 0 0.00054366 3.3 0.00054358 3.3 0.0005436799999999999 0 0.0005436000000000001 0 0.0005437 3.3 0.0005436200000000001 3.3 0.00054372 0 0.0005436400000000001 0 0.00054374 3.3 0.0005436600000000001 3.3 0.00054376 0 0.00054368 0 0.00054378 3.3 0.0005437 3.3 0.0005438 0 0.00054372 0 0.00054382 3.3 0.00054374 3.3 0.00054384 0 0.00054376 0 0.00054386 3.3 0.00054378 3.3 0.00054388 0 0.0005438 0 0.0005438999999999999 3.3 0.0005438200000000001 3.3 0.00054392 0 0.0005438400000000001 0 0.00054394 3.3 0.0005438600000000001 3.3 0.00054396 0 0.0005438800000000001 0 0.00054398 3.3 0.0005439 3.3 0.000544 0 0.00054392 0 0.00054402 3.3 0.00054394 3.3 0.00054404 0 0.00054396 0 0.00054406 3.3 0.00054398 3.3 0.00054408 0 0.000544 0 0.0005440999999999999 3.3 0.0005440200000000001 3.3 0.00054412 0 0.0005440400000000001 0 0.00054414 3.3 0.0005440600000000001 3.3 0.00054416 0 0.0005440800000000001 0 0.00054418 3.3 0.0005441 3.3 0.0005442 0 0.00054412 0 0.00054422 3.3 0.00054414 3.3 0.00054424 0 0.00054416 0 0.00054426 3.3 0.00054418 3.3 0.00054428 0 0.0005442 0 0.0005443 3.3 0.00054422 3.3 0.0005443199999999999 0 0.0005442400000000001 0 0.00054434 3.3 0.0005442600000000001 3.3 0.00054436 0 0.0005442800000000001 0 0.00054438 3.3 0.0005443000000000001 3.3 0.0005444 0 0.00054432 0 0.00054442 3.3 0.00054434 3.3 0.00054444 0 0.00054436 0 0.00054446 3.3 0.00054438 3.3 0.00054448 0 0.0005444 0 0.0005445 3.3 0.00054442 3.3 0.0005445199999999999 0 0.0005444400000000001 0 0.00054454 3.3 0.0005444600000000001 3.3 0.00054456 0 0.0005444800000000001 0 0.00054458 3.3 0.0005445000000000001 3.3 0.0005446 0 0.00054452 0 0.00054462 3.3 0.00054454 3.3 0.00054464 0 0.00054456 0 0.00054466 3.3 0.00054458 3.3 0.00054468 0 0.0005446 0 0.0005447 3.3 0.00054462 3.3 0.00054472 0 0.00054464 0 0.0005447399999999999 3.3 0.0005446600000000001 3.3 0.00054476 0 0.0005446800000000001 0 0.00054478 3.3 0.0005447000000000001 3.3 0.0005448 0 0.0005447200000000001 0 0.00054482 3.3 0.00054474 3.3 0.00054484 0 0.00054476 0 0.00054486 3.3 0.00054478 3.3 0.00054488 0 0.0005448 0 0.0005449 3.3 0.00054482 3.3 0.00054492 0 0.00054484 0 0.0005449399999999999 3.3 0.0005448600000000001 3.3 0.00054496 0 0.0005448800000000001 0 0.00054498 3.3 0.0005449000000000001 3.3 0.000545 0 0.0005449200000000001 0 0.00054502 3.3 0.00054494 3.3 0.00054504 0 0.00054496 0 0.00054506 3.3 0.00054498 3.3 0.00054508 0 0.000545 0 0.0005451 3.3 0.00054502 3.3 0.00054512 0 0.00054504 0 0.00054514 3.3 0.00054506 3.3 0.0005451599999999999 0 0.0005450800000000001 0 0.00054518 3.3 0.0005451000000000001 3.3 0.0005452 0 0.0005451200000000001 0 0.00054522 3.3 0.0005451400000000001 3.3 0.00054524 0 0.00054516 0 0.00054526 3.3 0.00054518 3.3 0.00054528 0 0.0005452 0 0.0005453 3.3 0.00054522 3.3 0.00054532 0 0.00054524 0 0.00054534 3.3 0.00054526 3.3 0.0005453599999999999 0 0.0005452800000000001 0 0.00054538 3.3 0.0005453000000000001 3.3 0.0005454 0 0.0005453200000000001 0 0.00054542 3.3 0.0005453400000000001 3.3 0.00054544 0 0.00054536 0 0.00054546 3.3 0.00054538 3.3 0.00054548 0 0.0005454 0 0.0005455 3.3 0.00054542 3.3 0.00054552 0 0.00054544 0 0.00054554 3.3 0.00054546 3.3 0.00054556 0 0.00054548 0 0.0005455799999999999 3.3 0.0005455000000000001 3.3 0.0005456 0 0.0005455200000000001 0 0.00054562 3.3 0.0005455400000000001 3.3 0.00054564 0 0.0005455600000000001 0 0.00054566 3.3 0.00054558 3.3 0.00054568 0 0.0005456 0 0.0005457 3.3 0.00054562 3.3 0.00054572 0 0.00054564 0 0.00054574 3.3 0.00054566 3.3 0.00054576 0 0.00054568 0 0.0005457799999999999 3.3 0.0005457000000000001 3.3 0.0005458 0 0.0005457200000000001 0 0.00054582 3.3 0.0005457400000000001 3.3 0.00054584 0 0.0005457600000000001 0 0.00054586 3.3 0.00054578 3.3 0.00054588 0 0.0005458 0 0.0005459 3.3 0.00054582 3.3 0.00054592 0 0.00054584 0 0.00054594 3.3 0.00054586 3.3 0.00054596 0 0.00054588 0 0.00054598 3.3 0.0005459 3.3 0.0005459999999999999 0 0.0005459200000000001 0 0.00054602 3.3 0.0005459400000000001 3.3 0.00054604 0 0.0005459600000000001 0 0.00054606 3.3 0.0005459800000000001 3.3 0.00054608 0 0.000546 0 0.0005461 3.3 0.00054602 3.3 0.00054612 0 0.00054604 0 0.00054614 3.3 0.00054606 3.3 0.00054616 0 0.00054608 0 0.00054618 3.3 0.0005461 3.3 0.0005461999999999999 0 0.0005461200000000001 0 0.00054622 3.3 0.0005461400000000001 3.3 0.00054624 0 0.0005461600000000001 0 0.00054626 3.3 0.0005461800000000001 3.3 0.00054628 0 0.0005462 0 0.0005463 3.3 0.00054622 3.3 0.00054632 0 0.00054624 0 0.00054634 3.3 0.00054626 3.3 0.00054636 0 0.00054628 0 0.00054638 3.3 0.0005463 3.3 0.0005463999999999999 0 0.00054632 0 0.0005464199999999999 3.3 0.0005463400000000001 3.3 0.00054644 0 0.0005463600000000001 0 0.00054646 3.3 0.0005463800000000001 3.3 0.00054648 0 0.0005464 0 0.0005465 3.3 0.00054642 3.3 0.00054652 0 0.00054644 0 0.00054654 3.3 0.00054646 3.3 0.00054656 0 0.00054648 0 0.00054658 3.3 0.0005465 3.3 0.0005466 0 0.00054652 0 0.0005466199999999999 3.3 0.0005465400000000001 3.3 0.00054664 0 0.0005465600000000001 0 0.00054666 3.3 0.0005465800000000001 3.3 0.00054668 0 0.0005466000000000001 0 0.0005467 3.3 0.00054662 3.3 0.00054672 0 0.00054664 0 0.00054674 3.3 0.00054666 3.3 0.00054676 0 0.00054668 0 0.00054678 3.3 0.0005467 3.3 0.0005468 0 0.00054672 0 0.0005468199999999999 3.3 0.0005467400000000001 3.3 0.00054684 0 0.0005467600000000001 0 0.00054686 3.3 0.0005467800000000001 3.3 0.00054688 0 0.0005468000000000001 0 0.0005469 3.3 0.00054682 3.3 0.00054692 0 0.00054684 0 0.00054694 3.3 0.00054686 3.3 0.00054696 0 0.00054688 0 0.00054698 3.3 0.0005469 3.3 0.000547 0 0.00054692 0 0.00054702 3.3 0.00054694 3.3 0.0005470399999999999 0 0.0005469600000000001 0 0.00054706 3.3 0.0005469800000000001 3.3 0.00054708 0 0.0005470000000000001 0 0.0005471 3.3 0.0005470200000000001 3.3 0.00054712 0 0.00054704 0 0.00054714 3.3 0.00054706 3.3 0.00054716 0 0.00054708 0 0.00054718 3.3 0.0005471 3.3 0.0005472 0 0.00054712 0 0.00054722 3.3 0.00054714 3.3 0.0005472399999999999 0 0.0005471600000000001 0 0.00054726 3.3 0.0005471800000000001 3.3 0.00054728 0 0.0005472000000000001 0 0.0005473 3.3 0.0005472200000000001 3.3 0.00054732 0 0.00054724 0 0.00054734 3.3 0.00054726 3.3 0.00054736 0 0.00054728 0 0.00054738 3.3 0.0005473 3.3 0.0005474 0 0.00054732 0 0.00054742 3.3 0.00054734 3.3 0.00054744 0 0.00054736 0 0.0005474599999999999 3.3 0.0005473800000000001 3.3 0.00054748 0 0.0005474000000000001 0 0.0005475 3.3 0.0005474200000000001 3.3 0.00054752 0 0.0005474400000000001 0 0.00054754 3.3 0.00054746 3.3 0.00054756 0 0.00054748 0 0.00054758 3.3 0.0005475 3.3 0.0005476 0 0.00054752 0 0.00054762 3.3 0.00054754 3.3 0.00054764 0 0.00054756 0 0.0005476599999999999 3.3 0.0005475800000000001 3.3 0.00054768 0 0.0005476000000000001 0 0.0005477 3.3 0.0005476200000000001 3.3 0.00054772 0 0.0005476400000000001 0 0.00054774 3.3 0.00054766 3.3 0.00054776 0 0.00054768 0 0.00054778 3.3 0.0005477 3.3 0.0005478 0 0.00054772 0 0.00054782 3.3 0.00054774 3.3 0.00054784 0 0.00054776 0 0.00054786 3.3 0.00054778 3.3 0.0005478799999999999 0 0.0005478000000000001 0 0.0005479 3.3 0.0005478200000000001 3.3 0.00054792 0 0.0005478400000000001 0 0.00054794 3.3 0.0005478600000000001 3.3 0.00054796 0 0.00054788 0 0.00054798 3.3 0.0005479 3.3 0.000548 0 0.00054792 0 0.00054802 3.3 0.00054794 3.3 0.00054804 0 0.00054796 0 0.00054806 3.3 0.00054798 3.3 0.0005480799999999999 0 0.0005480000000000001 0 0.0005481 3.3 0.0005480200000000001 3.3 0.00054812 0 0.0005480400000000001 0 0.00054814 3.3 0.0005480600000000001 3.3 0.00054816 0 0.00054808 0 0.00054818 3.3 0.0005481 3.3 0.0005482 0 0.00054812 0 0.00054822 3.3 0.00054814 3.3 0.00054824 0 0.00054816 0 0.00054826 3.3 0.00054818 3.3 0.00054828 0 0.0005482 0 0.0005482999999999999 3.3 0.0005482200000000001 3.3 0.00054832 0 0.0005482400000000001 0 0.00054834 3.3 0.0005482600000000001 3.3 0.00054836 0 0.0005482800000000001 0 0.00054838 3.3 0.0005483 3.3 0.0005484 0 0.00054832 0 0.00054842 3.3 0.00054834 3.3 0.00054844 0 0.00054836 0 0.00054846 3.3 0.00054838 3.3 0.00054848 0 0.0005484 0 0.0005484999999999999 3.3 0.0005484200000000001 3.3 0.00054852 0 0.0005484400000000001 0 0.00054854 3.3 0.0005484600000000001 3.3 0.00054856 0 0.0005484800000000001 0 0.00054858 3.3 0.0005485 3.3 0.0005486 0 0.00054852 0 0.00054862 3.3 0.00054854 3.3 0.00054864 0 0.00054856 0 0.00054866 3.3 0.00054858 3.3 0.00054868 0 0.0005486 0 0.0005487 3.3 0.00054862 3.3 0.0005487199999999999 0 0.0005486400000000001 0 0.00054874 3.3 0.0005486600000000001 3.3 0.00054876 0 0.0005486800000000001 0 0.00054878 3.3 0.0005487000000000001 3.3 0.0005488 0 0.00054872 0 0.00054882 3.3 0.00054874 3.3 0.00054884 0 0.00054876 0 0.00054886 3.3 0.00054878 3.3 0.00054888 0 0.0005488 0 0.0005489 3.3 0.00054882 3.3 0.0005489199999999999 0 0.0005488400000000001 0 0.00054894 3.3 0.0005488600000000001 3.3 0.00054896 0 0.0005488800000000001 0 0.00054898 3.3 0.0005489000000000001 3.3 0.000549 0 0.00054892 0 0.00054902 3.3 0.00054894 3.3 0.00054904 0 0.00054896 0 0.00054906 3.3 0.00054898 3.3 0.00054908 0 0.000549 0 0.0005491 3.3 0.00054902 3.3 0.00054912 0 0.00054904 0 0.0005491399999999999 3.3 0.0005490600000000001 3.3 0.00054916 0 0.0005490800000000001 0 0.00054918 3.3 0.0005491000000000001 3.3 0.0005492 0 0.0005491200000000001 0 0.00054922 3.3 0.00054914 3.3 0.00054924 0 0.00054916 0 0.00054926 3.3 0.00054918 3.3 0.00054928 0 0.0005492 0 0.0005493 3.3 0.00054922 3.3 0.00054932 0 0.00054924 0 0.0005493399999999999 3.3 0.0005492600000000001 3.3 0.00054936 0 0.0005492800000000001 0 0.00054938 3.3 0.0005493000000000001 3.3 0.0005494 0 0.0005493200000000001 0 0.00054942 3.3 0.00054934 3.3 0.00054944 0 0.00054936 0 0.00054946 3.3 0.00054938 3.3 0.00054948 0 0.0005494 0 0.0005495 3.3 0.00054942 3.3 0.00054952 0 0.00054944 0 0.00054954 3.3 0.00054946 3.3 0.0005495599999999999 0 0.0005494800000000001 0 0.00054958 3.3 0.0005495000000000001 3.3 0.0005496 0 0.0005495200000000001 0 0.00054962 3.3 0.0005495400000000001 3.3 0.00054964 0 0.00054956 0 0.00054966 3.3 0.00054958 3.3 0.00054968 0 0.0005496 0 0.0005497 3.3 0.00054962 3.3 0.00054972 0 0.00054964 0 0.00054974 3.3 0.00054966 3.3 0.0005497599999999999 0 0.0005496800000000001 0 0.00054978 3.3 0.0005497000000000001 3.3 0.0005498 0 0.0005497200000000001 0 0.00054982 3.3 0.0005497400000000001 3.3 0.00054984 0 0.00054976 0 0.00054986 3.3 0.00054978 3.3 0.00054988 0 0.0005498 0 0.0005499 3.3 0.00054982 3.3 0.00054992 0 0.00054984 0 0.00054994 3.3 0.00054986 3.3 0.0005499599999999999 0 0.00054988 0 0.0005499799999999999 3.3 0.0005499000000000001 3.3 0.00055 0 0.0005499200000000001 0 0.00055002 3.3 0.0005499400000000001 3.3 0.00055004 0 0.00054996 0 0.00055006 3.3 0.00054998 3.3 0.00055008 0 0.00055 0 0.0005501 3.3 0.00055002 3.3 0.00055012 0 0.00055004 0 0.00055014 3.3 0.00055006 3.3 0.00055016 0 0.00055008 0 0.0005501799999999999 3.3 0.0005501000000000001 3.3 0.0005502 0 0.0005501200000000001 0 0.00055022 3.3 0.0005501400000000001 3.3 0.00055024 0 0.0005501600000000001 0 0.00055026 3.3 0.00055018 3.3 0.00055028 0 0.0005502 0 0.0005503 3.3 0.00055022 3.3 0.00055032 0 0.00055024 0 0.00055034 3.3 0.00055026 3.3 0.00055036 0 0.00055028 0 0.0005503799999999999 3.3 0.0005503000000000001 3.3 0.0005504 0 0.0005503200000000001 0 0.00055042 3.3 0.0005503400000000001 3.3 0.00055044 0 0.0005503600000000001 0 0.00055046 3.3 0.00055038 3.3 0.00055048 0 0.0005504 0 0.0005505 3.3 0.00055042 3.3 0.00055052 0 0.00055044 0 0.00055054 3.3 0.00055046 3.3 0.00055056 0 0.00055048 0 0.00055058 3.3 0.0005505 3.3 0.0005505999999999999 0 0.0005505200000000001 0 0.00055062 3.3 0.0005505400000000001 3.3 0.00055064 0 0.0005505600000000001 0 0.00055066 3.3 0.0005505800000000001 3.3 0.00055068 0 0.0005506 0 0.0005507 3.3 0.00055062 3.3 0.00055072 0 0.00055064 0 0.00055074 3.3 0.00055066 3.3 0.00055076 0 0.00055068 0 0.00055078 3.3 0.0005507 3.3 0.0005507999999999999 0 0.0005507200000000001 0 0.00055082 3.3 0.0005507400000000001 3.3 0.00055084 0 0.0005507600000000001 0 0.00055086 3.3 0.0005507800000000001 3.3 0.00055088 0 0.0005508 0 0.0005509 3.3 0.00055082 3.3 0.00055092 0 0.00055084 0 0.00055094 3.3 0.00055086 3.3 0.00055096 0 0.00055088 0 0.00055098 3.3 0.0005509 3.3 0.000551 0 0.00055092 0 0.0005510199999999999 3.3 0.0005509400000000001 3.3 0.00055104 0 0.0005509600000000001 0 0.00055106 3.3 0.0005509800000000001 3.3 0.00055108 0 0.0005510000000000001 0 0.0005511 3.3 0.00055102 3.3 0.00055112 0 0.00055104 0 0.00055114 3.3 0.00055106 3.3 0.00055116 0 0.00055108 0 0.00055118 3.3 0.0005511 3.3 0.0005512 0 0.00055112 0 0.0005512199999999999 3.3 0.0005511400000000001 3.3 0.00055124 0 0.0005511600000000001 0 0.00055126 3.3 0.0005511800000000001 3.3 0.00055128 0 0.0005512000000000001 0 0.0005513 3.3 0.00055122 3.3 0.00055132 0 0.00055124 0 0.00055134 3.3 0.00055126 3.3 0.00055136 0 0.00055128 0 0.00055138 3.3 0.0005513 3.3 0.0005514 0 0.00055132 0 0.00055142 3.3 0.00055134 3.3 0.0005514399999999999 0 0.0005513600000000001 0 0.00055146 3.3 0.0005513800000000001 3.3 0.00055148 0 0.0005514000000000001 0 0.0005515 3.3 0.0005514200000000001 3.3 0.00055152 0 0.00055144 0 0.00055154 3.3 0.00055146 3.3 0.00055156 0 0.00055148 0 0.00055158 3.3 0.0005515 3.3 0.0005516 0 0.00055152 0 0.00055162 3.3 0.00055154 3.3 0.0005516399999999999 0 0.0005515600000000001 0 0.00055166 3.3 0.0005515800000000001 3.3 0.00055168 0 0.0005516000000000001 0 0.0005517 3.3 0.0005516200000000001 3.3 0.00055172 0 0.00055164 0 0.00055174 3.3 0.00055166 3.3 0.00055176 0 0.00055168 0 0.00055178 3.3 0.0005517 3.3 0.0005518 0 0.00055172 0 0.00055182 3.3 0.00055174 3.3 0.00055184 0 0.00055176 0 0.0005518599999999999 3.3 0.0005517800000000001 3.3 0.00055188 0 0.0005518000000000001 0 0.0005519 3.3 0.0005518200000000001 3.3 0.00055192 0 0.0005518400000000001 0 0.00055194 3.3 0.00055186 3.3 0.00055196 0 0.00055188 0 0.00055198 3.3 0.0005519 3.3 0.000552 0 0.00055192 0 0.00055202 3.3 0.00055194 3.3 0.00055204 0 0.00055196 0 0.0005520599999999999 3.3 0.0005519800000000001 3.3 0.00055208 0 0.0005520000000000001 0 0.0005521 3.3 0.0005520200000000001 3.3 0.00055212 0 0.0005520400000000001 0 0.00055214 3.3 0.00055206 3.3 0.00055216 0 0.00055208 0 0.00055218 3.3 0.0005521 3.3 0.0005522 0 0.00055212 0 0.00055222 3.3 0.00055214 3.3 0.00055224 0 0.00055216 0 0.00055226 3.3 0.00055218 3.3 0.0005522799999999999 0 0.0005522000000000001 0 0.0005523 3.3 0.0005522200000000001 3.3 0.00055232 0 0.0005522400000000001 0 0.00055234 3.3 0.0005522600000000001 3.3 0.00055236 0 0.00055228 0 0.00055238 3.3 0.0005523 3.3 0.0005524 0 0.00055232 0 0.00055242 3.3 0.00055234 3.3 0.00055244 0 0.00055236 0 0.00055246 3.3 0.00055238 3.3 0.0005524799999999999 0 0.0005524000000000001 0 0.0005525 3.3 0.0005524200000000001 3.3 0.00055252 0 0.0005524400000000001 0 0.00055254 3.3 0.0005524600000000001 3.3 0.00055256 0 0.00055248 0 0.00055258 3.3 0.0005525 3.3 0.0005526 0 0.00055252 0 0.00055262 3.3 0.00055254 3.3 0.00055264 0 0.00055256 0 0.00055266 3.3 0.00055258 3.3 0.00055268 0 0.0005526 0 0.0005526999999999999 3.3 0.0005526200000000001 3.3 0.00055272 0 0.0005526400000000001 0 0.00055274 3.3 0.0005526600000000001 3.3 0.00055276 0 0.0005526800000000001 0 0.00055278 3.3 0.0005527 3.3 0.0005528 0 0.00055272 0 0.00055282 3.3 0.00055274 3.3 0.00055284 0 0.00055276 0 0.00055286 3.3 0.00055278 3.3 0.00055288 0 0.0005528 0 0.0005528999999999999 3.3 0.0005528200000000001 3.3 0.00055292 0 0.0005528400000000001 0 0.00055294 3.3 0.0005528600000000001 3.3 0.00055296 0 0.0005528800000000001 0 0.00055298 3.3 0.0005529 3.3 0.000553 0 0.00055292 0 0.00055302 3.3 0.00055294 3.3 0.00055304 0 0.00055296 0 0.00055306 3.3 0.00055298 3.3 0.00055308 0 0.000553 0 0.0005531 3.3 0.00055302 3.3 0.0005531199999999999 0 0.0005530400000000001 0 0.00055314 3.3 0.0005530600000000001 3.3 0.00055316 0 0.0005530800000000001 0 0.00055318 3.3 0.0005531000000000001 3.3 0.0005532 0 0.00055312 0 0.00055322 3.3 0.00055314 3.3 0.00055324 0 0.00055316 0 0.00055326 3.3 0.00055318 3.3 0.00055328 0 0.0005532 0 0.0005533 3.3 0.00055322 3.3 0.0005533199999999999 0 0.0005532400000000001 0 0.00055334 3.3 0.0005532600000000001 3.3 0.00055336 0 0.0005532800000000001 0 0.00055338 3.3 0.0005533000000000001 3.3 0.0005534 0 0.00055332 0 0.00055342 3.3 0.00055334 3.3 0.00055344 0 0.00055336 0 0.00055346 3.3 0.00055338 3.3 0.00055348 0 0.0005534 0 0.0005535 3.3 0.00055342 3.3 0.0005535199999999999 0 0.00055344 0 0.0005535399999999999 3.3 0.0005534600000000001 3.3 0.00055356 0 0.0005534800000000001 0 0.00055358 3.3 0.0005535000000000001 3.3 0.0005536 0 0.00055352 0 0.00055362 3.3 0.00055354 3.3 0.00055364 0 0.00055356 0 0.00055366 3.3 0.00055358 3.3 0.00055368 0 0.0005536 0 0.0005537 3.3 0.00055362 3.3 0.00055372 0 0.00055364 0 0.0005537399999999999 3.3 0.0005536600000000001 3.3 0.00055376 0 0.0005536800000000001 0 0.00055378 3.3 0.0005537000000000001 3.3 0.0005538 0 0.0005537200000000001 0 0.00055382 3.3 0.00055374 3.3 0.00055384 0 0.00055376 0 0.00055386 3.3 0.00055378 3.3 0.00055388 0 0.0005538 0 0.0005539 3.3 0.00055382 3.3 0.00055392 0 0.00055384 0 0.0005539399999999999 3.3 0.0005538600000000001 3.3 0.00055396 0 0.0005538800000000001 0 0.00055398 3.3 0.0005539000000000001 3.3 0.000554 0 0.0005539200000000001 0 0.00055402 3.3 0.00055394 3.3 0.00055404 0 0.00055396 0 0.00055406 3.3 0.00055398 3.3 0.00055408 0 0.000554 0 0.0005541 3.3 0.00055402 3.3 0.00055412 0 0.00055404 0 0.00055414 3.3 0.00055406 3.3 0.0005541599999999999 0 0.0005540800000000001 0 0.00055418 3.3 0.0005541000000000001 3.3 0.0005542 0 0.0005541200000000001 0 0.00055422 3.3 0.0005541400000000001 3.3 0.00055424 0 0.00055416 0 0.00055426 3.3 0.00055418 3.3 0.00055428 0 0.0005542 0 0.0005543 3.3 0.00055422 3.3 0.00055432 0 0.00055424 0 0.00055434 3.3 0.00055426 3.3 0.0005543599999999999 0 0.0005542800000000001 0 0.00055438 3.3 0.0005543000000000001 3.3 0.0005544 0 0.0005543200000000001 0 0.00055442 3.3 0.0005543400000000001 3.3 0.00055444 0 0.00055436 0 0.00055446 3.3 0.00055438 3.3 0.00055448 0 0.0005544 0 0.0005545 3.3 0.00055442 3.3 0.00055452 0 0.00055444 0 0.00055454 3.3 0.00055446 3.3 0.00055456 0 0.00055448 0 0.0005545799999999999 3.3 0.0005545000000000001 3.3 0.0005546 0 0.0005545200000000001 0 0.00055462 3.3 0.0005545400000000001 3.3 0.00055464 0 0.0005545600000000001 0 0.00055466 3.3 0.00055458 3.3 0.00055468 0 0.0005546 0 0.0005547 3.3 0.00055462 3.3 0.00055472 0 0.00055464 0 0.00055474 3.3 0.00055466 3.3 0.00055476 0 0.00055468 0 0.0005547799999999999 3.3 0.0005547000000000001 3.3 0.0005548 0 0.0005547200000000001 0 0.00055482 3.3 0.0005547400000000001 3.3 0.00055484 0 0.0005547600000000001 0 0.00055486 3.3 0.00055478 3.3 0.00055488 0 0.0005548 0 0.0005549 3.3 0.00055482 3.3 0.00055492 0 0.00055484 0 0.00055494 3.3 0.00055486 3.3 0.00055496 0 0.00055488 0 0.00055498 3.3 0.0005549 3.3 0.0005549999999999999 0 0.0005549200000000001 0 0.00055502 3.3 0.0005549400000000001 3.3 0.00055504 0 0.0005549600000000001 0 0.00055506 3.3 0.0005549800000000001 3.3 0.00055508 0 0.000555 0 0.0005551 3.3 0.00055502 3.3 0.00055512 0 0.00055504 0 0.00055514 3.3 0.00055506 3.3 0.00055516 0 0.00055508 0 0.00055518 3.3 0.0005551 3.3 0.0005551999999999999 0 0.0005551200000000001 0 0.00055522 3.3 0.0005551400000000001 3.3 0.00055524 0 0.0005551600000000001 0 0.00055526 3.3 0.0005551800000000001 3.3 0.00055528 0 0.0005552 0 0.0005553 3.3 0.00055522 3.3 0.00055532 0 0.00055524 0 0.00055534 3.3 0.00055526 3.3 0.00055536 0 0.00055528 0 0.00055538 3.3 0.0005553 3.3 0.0005554 0 0.00055532 0 0.0005554199999999999 3.3 0.0005553400000000001 3.3 0.00055544 0 0.0005553600000000001 0 0.00055546 3.3 0.0005553800000000001 3.3 0.00055548 0 0.0005554000000000001 0 0.0005555 3.3 0.00055542 3.3 0.00055552 0 0.00055544 0 0.00055554 3.3 0.00055546 3.3 0.00055556 0 0.00055548 0 0.00055558 3.3 0.0005555 3.3 0.0005556 0 0.00055552 0 0.0005556199999999999 3.3 0.0005555400000000001 3.3 0.00055564 0 0.0005555600000000001 0 0.00055566 3.3 0.0005555800000000001 3.3 0.00055568 0 0.0005556000000000001 0 0.0005557 3.3 0.00055562 3.3 0.00055572 0 0.00055564 0 0.00055574 3.3 0.00055566 3.3 0.00055576 0 0.00055568 0 0.00055578 3.3 0.0005557 3.3 0.0005558 0 0.00055572 0 0.00055582 3.3 0.00055574 3.3 0.0005558399999999999 0 0.0005557600000000001 0 0.00055586 3.3 0.0005557800000000001 3.3 0.00055588 0 0.0005558000000000001 0 0.0005559 3.3 0.0005558200000000001 3.3 0.00055592 0 0.00055584 0 0.00055594 3.3 0.00055586 3.3 0.00055596 0 0.00055588 0 0.00055598 3.3 0.0005559 3.3 0.000556 0 0.00055592 0 0.00055602 3.3 0.00055594 3.3 0.0005560399999999999 0 0.0005559600000000001 0 0.00055606 3.3 0.0005559800000000001 3.3 0.00055608 0 0.0005560000000000001 0 0.0005561 3.3 0.0005560200000000001 3.3 0.00055612 0 0.00055604 0 0.00055614 3.3 0.00055606 3.3 0.00055616 0 0.00055608 0 0.00055618 3.3 0.0005561 3.3 0.0005562 0 0.00055612 0 0.00055622 3.3 0.00055614 3.3 0.00055624 0 0.00055616 0 0.0005562599999999999 3.3 0.0005561800000000001 3.3 0.00055628 0 0.0005562000000000001 0 0.0005563 3.3 0.0005562200000000001 3.3 0.00055632 0 0.0005562400000000001 0 0.00055634 3.3 0.00055626 3.3 0.00055636 0 0.00055628 0 0.00055638 3.3 0.0005563 3.3 0.0005564 0 0.00055632 0 0.00055642 3.3 0.00055634 3.3 0.00055644 0 0.00055636 0 0.0005564599999999999 3.3 0.0005563800000000001 3.3 0.00055648 0 0.0005564000000000001 0 0.0005565 3.3 0.0005564200000000001 3.3 0.00055652 0 0.0005564400000000001 0 0.00055654 3.3 0.00055646 3.3 0.00055656 0 0.00055648 0 0.00055658 3.3 0.0005565 3.3 0.0005566 0 0.00055652 0 0.00055662 3.3 0.00055654 3.3 0.00055664 0 0.00055656 0 0.0005566599999999999 3.3 0.00055658 3.3 0.0005566799999999999 0 0.0005566000000000001 0 0.0005567 3.3 0.0005566200000000001 3.3 0.00055672 0 0.0005566400000000001 0 0.00055674 3.3 0.00055666 3.3 0.00055676 0 0.00055668 0 0.00055678 3.3 0.0005567 3.3 0.0005568 0 0.00055672 0 0.00055682 3.3 0.00055674 3.3 0.00055684 0 0.00055676 0 0.00055686 3.3 0.00055678 3.3 0.0005568799999999999 0 0.0005568000000000001 0 0.0005569 3.3 0.0005568200000000001 3.3 0.00055692 0 0.0005568400000000001 0 0.00055694 3.3 0.0005568600000000001 3.3 0.00055696 0 0.00055688 0 0.00055698 3.3 0.0005569 3.3 0.000557 0 0.00055692 0 0.00055702 3.3 0.00055694 3.3 0.00055704 0 0.00055696 0 0.00055706 3.3 0.00055698 3.3 0.0005570799999999999 0 0.000557 0 0.0005570999999999999 3.3 0.0005570200000000001 3.3 0.00055712 0 0.0005570400000000001 0 0.00055714 3.3 0.0005570600000000001 3.3 0.00055716 0 0.00055708 0 0.00055718 3.3 0.0005571 3.3 0.0005572 0 0.00055712 0 0.00055722 3.3 0.00055714 3.3 0.00055724 0 0.00055716 0 0.00055726 3.3 0.00055718 3.3 0.00055728 0 0.0005572 0 0.0005572999999999999 3.3 0.0005572200000000001 3.3 0.00055732 0 0.0005572400000000001 0 0.00055734 3.3 0.0005572600000000001 3.3 0.00055736 0 0.0005572800000000001 0 0.00055738 3.3 0.0005573 3.3 0.0005574 0 0.00055732 0 0.00055742 3.3 0.00055734 3.3 0.00055744 0 0.00055736 0 0.00055746 3.3 0.00055738 3.3 0.00055748 0 0.0005574 0 0.0005574999999999999 3.3 0.0005574200000000001 3.3 0.00055752 0 0.0005574400000000001 0 0.00055754 3.3 0.0005574600000000001 3.3 0.00055756 0 0.0005574800000000001 0 0.00055758 3.3 0.0005575 3.3 0.0005576 0 0.00055752 0 0.00055762 3.3 0.00055754 3.3 0.00055764 0 0.00055756 0 0.00055766 3.3 0.00055758 3.3 0.00055768 0 0.0005576 0 0.0005577 3.3 0.00055762 3.3 0.0005577199999999999 0 0.0005576400000000001 0 0.00055774 3.3 0.0005576600000000001 3.3 0.00055776 0 0.0005576800000000001 0 0.00055778 3.3 0.0005577000000000001 3.3 0.0005578 0 0.00055772 0 0.00055782 3.3 0.00055774 3.3 0.00055784 0 0.00055776 0 0.00055786 3.3 0.00055778 3.3 0.00055788 0 0.0005578 0 0.0005579 3.3 0.00055782 3.3 0.0005579199999999999 0 0.0005578400000000001 0 0.00055794 3.3 0.0005578600000000001 3.3 0.00055796 0 0.0005578800000000001 0 0.00055798 3.3 0.0005579000000000001 3.3 0.000558 0 0.00055792 0 0.00055802 3.3 0.00055794 3.3 0.00055804 0 0.00055796 0 0.00055806 3.3 0.00055798 3.3 0.00055808 0 0.000558 0 0.0005581 3.3 0.00055802 3.3 0.00055812 0 0.00055804 0 0.0005581399999999999 3.3 0.0005580600000000001 3.3 0.00055816 0 0.0005580800000000001 0 0.00055818 3.3 0.0005581000000000001 3.3 0.0005582 0 0.0005581200000000001 0 0.00055822 3.3 0.00055814 3.3 0.00055824 0 0.00055816 0 0.00055826 3.3 0.00055818 3.3 0.00055828 0 0.0005582 0 0.0005583 3.3 0.00055822 3.3 0.00055832 0 0.00055824 0 0.0005583399999999999 3.3 0.0005582600000000001 3.3 0.00055836 0 0.0005582800000000001 0 0.00055838 3.3 0.0005583000000000001 3.3 0.0005584 0 0.0005583200000000001 0 0.00055842 3.3 0.00055834 3.3 0.00055844 0 0.00055836 0 0.00055846 3.3 0.00055838 3.3 0.00055848 0 0.0005584 0 0.0005585 3.3 0.00055842 3.3 0.00055852 0 0.00055844 0 0.00055854 3.3 0.00055846 3.3 0.0005585599999999999 0 0.0005584800000000001 0 0.00055858 3.3 0.0005585000000000001 3.3 0.0005586 0 0.0005585200000000001 0 0.00055862 3.3 0.0005585400000000001 3.3 0.00055864 0 0.00055856 0 0.00055866 3.3 0.00055858 3.3 0.00055868 0 0.0005586 0 0.0005587 3.3 0.00055862 3.3 0.00055872 0 0.00055864 0 0.00055874 3.3 0.00055866 3.3 0.0005587599999999999 0 0.0005586800000000001 0 0.00055878 3.3 0.0005587000000000001 3.3 0.0005588 0 0.0005587200000000001 0 0.00055882 3.3 0.0005587400000000001 3.3 0.00055884 0 0.00055876 0 0.00055886 3.3 0.00055878 3.3 0.00055888 0 0.0005588 0 0.0005589 3.3 0.00055882 3.3 0.00055892 0 0.00055884 0 0.00055894 3.3 0.00055886 3.3 0.00055896 0 0.00055888 0 0.0005589799999999999 3.3 0.0005589000000000001 3.3 0.000559 0 0.0005589200000000001 0 0.00055902 3.3 0.0005589400000000001 3.3 0.00055904 0 0.0005589600000000001 0 0.00055906 3.3 0.00055898 3.3 0.00055908 0 0.000559 0 0.0005591 3.3 0.00055902 3.3 0.00055912 0 0.00055904 0 0.00055914 3.3 0.00055906 3.3 0.00055916 0 0.00055908 0 0.0005591799999999999 3.3 0.0005591000000000001 3.3 0.0005592 0 0.0005591200000000001 0 0.00055922 3.3 0.0005591400000000001 3.3 0.00055924 0 0.0005591600000000001 0 0.00055926 3.3 0.00055918 3.3 0.00055928 0 0.0005592 0 0.0005593 3.3 0.00055922 3.3 0.00055932 0 0.00055924 0 0.00055934 3.3 0.00055926 3.3 0.00055936 0 0.00055928 0 0.00055938 3.3 0.0005593 3.3 0.0005593999999999999 0 0.0005593200000000001 0 0.00055942 3.3 0.0005593400000000001 3.3 0.00055944 0 0.0005593600000000001 0 0.00055946 3.3 0.0005593800000000001 3.3 0.00055948 0 0.0005594 0 0.0005595 3.3 0.00055942 3.3 0.00055952 0 0.00055944 0 0.00055954 3.3 0.00055946 3.3 0.00055956 0 0.00055948 0 0.00055958 3.3 0.0005595 3.3 0.0005595999999999999 0 0.0005595200000000001 0 0.00055962 3.3 0.0005595400000000001 3.3 0.00055964 0 0.0005595600000000001 0 0.00055966 3.3 0.0005595800000000001 3.3 0.00055968 0 0.0005596 0 0.0005597 3.3 0.00055962 3.3 0.00055972 0 0.00055964 0 0.00055974 3.3 0.00055966 3.3 0.00055976 0 0.00055968 0 0.00055978 3.3 0.0005597 3.3 0.0005598 0 0.00055972 0 0.0005598199999999999 3.3 0.0005597400000000001 3.3 0.00055984 0 0.0005597600000000001 0 0.00055986 3.3 0.0005597800000000001 3.3 0.00055988 0 0.0005598000000000001 0 0.0005599 3.3 0.00055982 3.3 0.00055992 0 0.00055984 0 0.00055994 3.3 0.00055986 3.3 0.00055996 0 0.00055988 0 0.00055998 3.3 0.0005599 3.3 0.00056 0 0.00055992 0 0.0005600199999999999 3.3 0.0005599400000000001 3.3 0.00056004 0 0.0005599600000000001 0 0.00056006 3.3 0.0005599800000000001 3.3 0.00056008 0 0.0005600000000000001 0 0.0005601 3.3 0.00056002 3.3 0.00056012 0 0.00056004 0 0.00056014 3.3 0.00056006 3.3 0.00056016 0 0.00056008 0 0.00056018 3.3 0.0005601 3.3 0.0005602 0 0.00056012 0 0.0005602199999999999 3.3 0.00056014 3.3 0.0005602399999999999 0 0.0005601600000000001 0 0.00056026 3.3 0.0005601800000000001 3.3 0.00056028 0 0.0005602000000000001 0 0.0005603 3.3 0.00056022 3.3 0.00056032 0 0.00056024 0 0.00056034 3.3 0.00056026 3.3 0.00056036 0 0.00056028 0 0.00056038 3.3 0.0005603 3.3 0.0005604 0 0.00056032 0 0.00056042 3.3 0.00056034 3.3 0.0005604399999999999 0 0.0005603600000000001 0 0.00056046 3.3 0.0005603800000000001 3.3 0.00056048 0 0.0005604000000000001 0 0.0005605 3.3 0.0005604200000000001 3.3 0.00056052 0 0.00056044 0 0.00056054 3.3 0.00056046 3.3 0.00056056 0 0.00056048 0 0.00056058 3.3 0.0005605 3.3 0.0005606 0 0.00056052 0 0.00056062 3.3 0.00056054 3.3 0.0005606399999999999 0 0.0005605600000000001 0 0.00056066 3.3 0.0005605800000000001 3.3 0.00056068 0 0.0005606000000000001 0 0.0005607 3.3 0.0005606200000000001 3.3 0.00056072 0 0.00056064 0 0.00056074 3.3 0.00056066 3.3 0.00056076 0 0.00056068 0 0.00056078 3.3 0.0005607 3.3 0.0005608 0 0.00056072 0 0.00056082 3.3 0.00056074 3.3 0.00056084 0 0.00056076 0 0.0005608599999999999 3.3 0.0005607800000000001 3.3 0.00056088 0 0.0005608000000000001 0 0.0005609 3.3 0.0005608200000000001 3.3 0.00056092 0 0.0005608400000000001 0 0.00056094 3.3 0.00056086 3.3 0.00056096 0 0.00056088 0 0.00056098 3.3 0.0005609 3.3 0.000561 0 0.00056092 0 0.00056102 3.3 0.00056094 3.3 0.00056104 0 0.00056096 0 0.0005610599999999999 3.3 0.0005609800000000001 3.3 0.00056108 0 0.0005610000000000001 0 0.0005611 3.3 0.0005610200000000001 3.3 0.00056112 0 0.0005610400000000001 0 0.00056114 3.3 0.00056106 3.3 0.00056116 0 0.00056108 0 0.00056118 3.3 0.0005611 3.3 0.0005612 0 0.00056112 0 0.00056122 3.3 0.00056114 3.3 0.00056124 0 0.00056116 0 0.00056126 3.3 0.00056118 3.3 0.0005612799999999999 0 0.0005612000000000001 0 0.0005613 3.3 0.0005612200000000001 3.3 0.00056132 0 0.0005612400000000001 0 0.00056134 3.3 0.0005612600000000001 3.3 0.00056136 0 0.00056128 0 0.00056138 3.3 0.0005613 3.3 0.0005614 0 0.00056132 0 0.00056142 3.3 0.00056134 3.3 0.00056144 0 0.00056136 0 0.00056146 3.3 0.00056138 3.3 0.0005614799999999999 0 0.0005614000000000001 0 0.0005615 3.3 0.0005614200000000001 3.3 0.00056152 0 0.0005614400000000001 0 0.00056154 3.3 0.0005614600000000001 3.3 0.00056156 0 0.00056148 0 0.00056158 3.3 0.0005615 3.3 0.0005616 0 0.00056152 0 0.00056162 3.3 0.00056154 3.3 0.00056164 0 0.00056156 0 0.00056166 3.3 0.00056158 3.3 0.00056168 0 0.0005616 0 0.0005616999999999999 3.3 0.0005616200000000001 3.3 0.00056172 0 0.0005616400000000001 0 0.00056174 3.3 0.0005616600000000001 3.3 0.00056176 0 0.0005616800000000001 0 0.00056178 3.3 0.0005617 3.3 0.0005618 0 0.00056172 0 0.00056182 3.3 0.00056174 3.3 0.00056184 0 0.00056176 0 0.00056186 3.3 0.00056178 3.3 0.00056188 0 0.0005618 0 0.0005618999999999999 3.3 0.0005618200000000001 3.3 0.00056192 0 0.0005618400000000001 0 0.00056194 3.3 0.0005618600000000001 3.3 0.00056196 0 0.0005618800000000001 0 0.00056198 3.3 0.0005619 3.3 0.000562 0 0.00056192 0 0.00056202 3.3 0.00056194 3.3 0.00056204 0 0.00056196 0 0.00056206 3.3 0.00056198 3.3 0.00056208 0 0.000562 0 0.0005621 3.3 0.00056202 3.3 0.0005621199999999999 0 0.0005620400000000001 0 0.00056214 3.3 0.0005620600000000001 3.3 0.00056216 0 0.0005620800000000001 0 0.00056218 3.3 0.0005621000000000001 3.3 0.0005622 0 0.00056212 0 0.00056222 3.3 0.00056214 3.3 0.00056224 0 0.00056216 0 0.00056226 3.3 0.00056218 3.3 0.00056228 0 0.0005622 0 0.0005623 3.3 0.00056222 3.3 0.0005623199999999999 0 0.0005622400000000001 0 0.00056234 3.3 0.0005622600000000001 3.3 0.00056236 0 0.0005622800000000001 0 0.00056238 3.3 0.0005623000000000001 3.3 0.0005624 0 0.00056232 0 0.00056242 3.3 0.00056234 3.3 0.00056244 0 0.00056236 0 0.00056246 3.3 0.00056238 3.3 0.00056248 0 0.0005624 0 0.0005625 3.3 0.00056242 3.3 0.00056252 0 0.00056244 0 0.0005625399999999999 3.3 0.0005624600000000001 3.3 0.00056256 0 0.0005624800000000001 0 0.00056258 3.3 0.0005625000000000001 3.3 0.0005626 0 0.0005625200000000001 0 0.00056262 3.3 0.00056254 3.3 0.00056264 0 0.00056256 0 0.00056266 3.3 0.00056258 3.3 0.00056268 0 0.0005626 0 0.0005627 3.3 0.00056262 3.3 0.00056272 0 0.00056264 0 0.0005627399999999999 3.3 0.0005626600000000001 3.3 0.00056276 0 0.0005626800000000001 0 0.00056278 3.3 0.0005627000000000001 3.3 0.0005628 0 0.0005627200000000001 0 0.00056282 3.3 0.00056274 3.3 0.00056284 0 0.00056276 0 0.00056286 3.3 0.00056278 3.3 0.00056288 0 0.0005628 0 0.0005629 3.3 0.00056282 3.3 0.00056292 0 0.00056284 0 0.00056294 3.3 0.00056286 3.3 0.0005629599999999999 0 0.0005628800000000001 0 0.00056298 3.3 0.0005629000000000001 3.3 0.000563 0 0.0005629200000000001 0 0.00056302 3.3 0.0005629400000000001 3.3 0.00056304 0 0.00056296 0 0.00056306 3.3 0.00056298 3.3 0.00056308 0 0.000563 0 0.0005631 3.3 0.00056302 3.3 0.00056312 0 0.00056304 0 0.00056314 3.3 0.00056306 3.3 0.0005631599999999999 0 0.0005630800000000001 0 0.00056318 3.3 0.0005631000000000001 3.3 0.0005632 0 0.0005631200000000001 0 0.00056322 3.3 0.0005631400000000001 3.3 0.00056324 0 0.00056316 0 0.00056326 3.3 0.00056318 3.3 0.00056328 0 0.0005632 0 0.0005633 3.3 0.00056322 3.3 0.00056332 0 0.00056324 0 0.00056334 3.3 0.00056326 3.3 0.00056336 0 0.00056328 0 0.0005633799999999999 3.3 0.0005633000000000001 3.3 0.0005634 0 0.0005633200000000001 0 0.00056342 3.3 0.0005633400000000001 3.3 0.00056344 0 0.0005633600000000001 0 0.00056346 3.3 0.00056338 3.3 0.00056348 0 0.0005634 0 0.0005635 3.3 0.00056342 3.3 0.00056352 0 0.00056344 0 0.00056354 3.3 0.00056346 3.3 0.00056356 0 0.00056348 0 0.0005635799999999999 3.3 0.0005635000000000001 3.3 0.0005636 0 0.0005635200000000001 0 0.00056362 3.3 0.0005635400000000001 3.3 0.00056364 0 0.0005635600000000001 0 0.00056366 3.3 0.00056358 3.3 0.00056368 0 0.0005636 0 0.0005637 3.3 0.00056362 3.3 0.00056372 0 0.00056364 0 0.00056374 3.3 0.00056366 3.3 0.00056376 0 0.00056368 0 0.0005637799999999999 3.3 0.0005637 3.3 0.0005637999999999999 0 0.0005637200000000001 0 0.00056382 3.3 0.0005637400000000001 3.3 0.00056384 0 0.0005637600000000001 0 0.00056386 3.3 0.00056378 3.3 0.00056388 0 0.0005638 0 0.0005639 3.3 0.00056382 3.3 0.00056392 0 0.00056384 0 0.00056394 3.3 0.00056386 3.3 0.00056396 0 0.00056388 0 0.00056398 3.3 0.0005639 3.3 0.0005639999999999999 0 0.0005639200000000001 0 0.00056402 3.3 0.0005639400000000001 3.3 0.00056404 0 0.0005639600000000001 0 0.00056406 3.3 0.0005639800000000001 3.3 0.00056408 0 0.000564 0 0.0005641 3.3 0.00056402 3.3 0.00056412 0 0.00056404 0 0.00056414 3.3 0.00056406 3.3 0.00056416 0 0.00056408 0 0.00056418 3.3 0.0005641 3.3 0.0005641999999999999 0 0.0005641200000000001 0 0.00056422 3.3 0.0005641400000000001 3.3 0.00056424 0 0.0005641600000000001 0 0.00056426 3.3 0.0005641800000000001 3.3 0.00056428 0 0.0005642 0 0.0005643 3.3 0.00056422 3.3 0.00056432 0 0.00056424 0 0.00056434 3.3 0.00056426 3.3 0.00056436 0 0.00056428 0 0.00056438 3.3 0.0005643 3.3 0.0005644 0 0.00056432 0 0.0005644199999999999 3.3 0.0005643400000000001 3.3 0.00056444 0 0.0005643600000000001 0 0.00056446 3.3 0.0005643800000000001 3.3 0.00056448 0 0.0005644000000000001 0 0.0005645 3.3 0.00056442 3.3 0.00056452 0 0.00056444 0 0.00056454 3.3 0.00056446 3.3 0.00056456 0 0.00056448 0 0.00056458 3.3 0.0005645 3.3 0.0005646 0 0.00056452 0 0.0005646199999999999 3.3 0.0005645400000000001 3.3 0.00056464 0 0.0005645600000000001 0 0.00056466 3.3 0.0005645800000000001 3.3 0.00056468 0 0.0005646000000000001 0 0.0005647 3.3 0.00056462 3.3 0.00056472 0 0.00056464 0 0.00056474 3.3 0.00056466 3.3 0.00056476 0 0.00056468 0 0.00056478 3.3 0.0005647 3.3 0.0005648 0 0.00056472 0 0.00056482 3.3 0.00056474 3.3 0.0005648399999999999 0 0.0005647600000000001 0 0.00056486 3.3 0.0005647800000000001 3.3 0.00056488 0 0.0005648000000000001 0 0.0005649 3.3 0.0005648200000000001 3.3 0.00056492 0 0.00056484 0 0.00056494 3.3 0.00056486 3.3 0.00056496 0 0.00056488 0 0.00056498 3.3 0.0005649 3.3 0.000565 0 0.00056492 0 0.00056502 3.3 0.00056494 3.3 0.0005650399999999999 0 0.0005649600000000001 0 0.00056506 3.3 0.0005649800000000001 3.3 0.00056508 0 0.0005650000000000001 0 0.0005651 3.3 0.0005650200000000001 3.3 0.00056512 0 0.00056504 0 0.00056514 3.3 0.00056506 3.3 0.00056516 0 0.00056508 0 0.00056518 3.3 0.0005651 3.3 0.0005652 0 0.00056512 0 0.00056522 3.3 0.00056514 3.3 0.00056524 0 0.00056516 0 0.0005652599999999999 3.3 0.0005651800000000001 3.3 0.00056528 0 0.0005652000000000001 0 0.0005653 3.3 0.0005652200000000001 3.3 0.00056532 0 0.0005652400000000001 0 0.00056534 3.3 0.00056526 3.3 0.00056536 0 0.00056528 0 0.00056538 3.3 0.0005653 3.3 0.0005654 0 0.00056532 0 0.00056542 3.3 0.00056534 3.3 0.00056544 0 0.00056536 0 0.0005654599999999999 3.3 0.0005653800000000001 3.3 0.00056548 0 0.0005654000000000001 0 0.0005655 3.3 0.0005654200000000001 3.3 0.00056552 0 0.0005654400000000001 0 0.00056554 3.3 0.00056546 3.3 0.00056556 0 0.00056548 0 0.00056558 3.3 0.0005655 3.3 0.0005656 0 0.00056552 0 0.00056562 3.3 0.00056554 3.3 0.00056564 0 0.00056556 0 0.00056566 3.3 0.00056558 3.3 0.0005656799999999999 0 0.0005656000000000001 0 0.0005657 3.3 0.0005656200000000001 3.3 0.00056572 0 0.0005656400000000001 0 0.00056574 3.3 0.0005656600000000001 3.3 0.00056576 0 0.00056568 0 0.00056578 3.3 0.0005657 3.3 0.0005658 0 0.00056572 0 0.00056582 3.3 0.00056574 3.3 0.00056584 0 0.00056576 0 0.00056586 3.3 0.00056578 3.3 0.0005658799999999999 0 0.0005658000000000001 0 0.0005659 3.3 0.0005658200000000001 3.3 0.00056592 0 0.0005658400000000001 0 0.00056594 3.3 0.0005658600000000001 3.3 0.00056596 0 0.00056588 0 0.00056598 3.3 0.0005659 3.3 0.000566 0 0.00056592 0 0.00056602 3.3 0.00056594 3.3 0.00056604 0 0.00056596 0 0.00056606 3.3 0.00056598 3.3 0.00056608 0 0.000566 0 0.0005660999999999999 3.3 0.0005660200000000001 3.3 0.00056612 0 0.0005660400000000001 0 0.00056614 3.3 0.0005660600000000001 3.3 0.00056616 0 0.0005660800000000001 0 0.00056618 3.3 0.0005661 3.3 0.0005662 0 0.00056612 0 0.00056622 3.3 0.00056614 3.3 0.00056624 0 0.00056616 0 0.00056626 3.3 0.00056618 3.3 0.00056628 0 0.0005662 0 0.0005662999999999999 3.3 0.0005662200000000001 3.3 0.00056632 0 0.0005662400000000001 0 0.00056634 3.3 0.0005662600000000001 3.3 0.00056636 0 0.0005662800000000001 0 0.00056638 3.3 0.0005663 3.3 0.0005664 0 0.00056632 0 0.00056642 3.3 0.00056634 3.3 0.00056644 0 0.00056636 0 0.00056646 3.3 0.00056638 3.3 0.00056648 0 0.0005664 0 0.0005665 3.3 0.00056642 3.3 0.0005665199999999999 0 0.0005664400000000001 0 0.00056654 3.3 0.0005664600000000001 3.3 0.00056656 0 0.0005664800000000001 0 0.00056658 3.3 0.0005665000000000001 3.3 0.0005666 0 0.00056652 0 0.00056662 3.3 0.00056654 3.3 0.00056664 0 0.00056656 0 0.00056666 3.3 0.00056658 3.3 0.00056668 0 0.0005666 0 0.0005667 3.3 0.00056662 3.3 0.0005667199999999999 0 0.0005666400000000001 0 0.00056674 3.3 0.0005666600000000001 3.3 0.00056676 0 0.0005666800000000001 0 0.00056678 3.3 0.0005667000000000001 3.3 0.0005668 0 0.00056672 0 0.00056682 3.3 0.00056674 3.3 0.00056684 0 0.00056676 0 0.00056686 3.3 0.00056678 3.3 0.00056688 0 0.0005668 0 0.0005669 3.3 0.00056682 3.3 0.0005669199999999999 0 0.00056684 0 0.0005669399999999999 3.3 0.0005668600000000001 3.3 0.00056696 0 0.0005668800000000001 0 0.00056698 3.3 0.0005669000000000001 3.3 0.000567 0 0.00056692 0 0.00056702 3.3 0.00056694 3.3 0.00056704 0 0.00056696 0 0.00056706 3.3 0.00056698 3.3 0.00056708 0 0.000567 0 0.0005671 3.3 0.00056702 3.3 0.00056712 0 0.00056704 0 0.0005671399999999999 3.3 0.0005670600000000001 3.3 0.00056716 0 0.0005670800000000001 0 0.00056718 3.3 0.0005671000000000001 3.3 0.0005672 0 0.0005671200000000001 0 0.00056722 3.3 0.00056714 3.3 0.00056724 0 0.00056716 0 0.00056726 3.3 0.00056718 3.3 0.00056728 0 0.0005672 0 0.0005673 3.3 0.00056722 3.3 0.00056732 0 0.00056724 0 0.0005673399999999999 3.3 0.00056726 3.3 0.0005673599999999999 0 0.0005672800000000001 0 0.00056738 3.3 0.0005673000000000001 3.3 0.0005674 0 0.0005673200000000001 0 0.00056742 3.3 0.00056734 3.3 0.00056744 0 0.00056736 0 0.00056746 3.3 0.00056738 3.3 0.00056748 0 0.0005674 0 0.0005675 3.3 0.00056742 3.3 0.00056752 0 0.00056744 0 0.00056754 3.3 0.00056746 3.3 0.0005675599999999999 0 0.0005674800000000001 0 0.00056758 3.3 0.0005675000000000001 3.3 0.0005676 0 0.0005675200000000001 0 0.00056762 3.3 0.0005675400000000001 3.3 0.00056764 0 0.00056756 0 0.00056766 3.3 0.00056758 3.3 0.00056768 0 0.0005676 0 0.0005677 3.3 0.00056762 3.3 0.00056772 0 0.00056764 0 0.00056774 3.3 0.00056766 3.3 0.0005677599999999999 0 0.0005676800000000001 0 0.00056778 3.3 0.0005677000000000001 3.3 0.0005678 0 0.0005677200000000001 0 0.00056782 3.3 0.0005677400000000001 3.3 0.00056784 0 0.00056776 0 0.00056786 3.3 0.00056778 3.3 0.00056788 0 0.0005678 0 0.0005679 3.3 0.00056782 3.3 0.00056792 0 0.00056784 0 0.00056794 3.3 0.00056786 3.3 0.00056796 0 0.00056788 0 0.0005679799999999999 3.3 0.0005679000000000001 3.3 0.000568 0 0.0005679200000000001 0 0.00056802 3.3 0.0005679400000000001 3.3 0.00056804 0 0.0005679600000000001 0 0.00056806 3.3 0.00056798 3.3 0.00056808 0 0.000568 0 0.0005681 3.3 0.00056802 3.3 0.00056812 0 0.00056804 0 0.00056814 3.3 0.00056806 3.3 0.00056816 0 0.00056808 0 0.0005681799999999999 3.3 0.0005681000000000001 3.3 0.0005682 0 0.0005681200000000001 0 0.00056822 3.3 0.0005681400000000001 3.3 0.00056824 0 0.0005681600000000001 0 0.00056826 3.3 0.00056818 3.3 0.00056828 0 0.0005682 0 0.0005683 3.3 0.00056822 3.3 0.00056832 0 0.00056824 0 0.00056834 3.3 0.00056826 3.3 0.00056836 0 0.00056828 0 0.00056838 3.3 0.0005683 3.3 0.0005683999999999999 0 0.0005683200000000001 0 0.00056842 3.3 0.0005683400000000001 3.3 0.00056844 0 0.0005683600000000001 0 0.00056846 3.3 0.0005683800000000001 3.3 0.00056848 0 0.0005684 0 0.0005685 3.3 0.00056842 3.3 0.00056852 0 0.00056844 0 0.00056854 3.3 0.00056846 3.3 0.00056856 0 0.00056848 0 0.00056858 3.3 0.0005685 3.3 0.0005685999999999999 0 0.0005685200000000001 0 0.00056862 3.3 0.0005685400000000001 3.3 0.00056864 0 0.0005685600000000001 0 0.00056866 3.3 0.0005685800000000001 3.3 0.00056868 0 0.0005686 0 0.0005687 3.3 0.00056862 3.3 0.00056872 0 0.00056864 0 0.00056874 3.3 0.00056866 3.3 0.00056876 0 0.00056868 0 0.00056878 3.3 0.0005687 3.3 0.0005688 0 0.00056872 0 0.0005688199999999999 3.3 0.0005687400000000001 3.3 0.00056884 0 0.0005687600000000001 0 0.00056886 3.3 0.0005687800000000001 3.3 0.00056888 0 0.0005688000000000001 0 0.0005689 3.3 0.00056882 3.3 0.00056892 0 0.00056884 0 0.00056894 3.3 0.00056886 3.3 0.00056896 0 0.00056888 0 0.00056898 3.3 0.0005689 3.3 0.000569 0 0.00056892 0 0.0005690199999999999 3.3 0.0005689400000000001 3.3 0.00056904 0 0.0005689600000000001 0 0.00056906 3.3 0.0005689800000000001 3.3 0.00056908 0 0.0005690000000000001 0 0.0005691 3.3 0.00056902 3.3 0.00056912 0 0.00056904 0 0.00056914 3.3 0.00056906 3.3 0.00056916 0 0.00056908 0 0.00056918 3.3 0.0005691 3.3 0.0005692 0 0.00056912 0 0.00056922 3.3 0.00056914 3.3 0.0005692399999999999 0 0.0005691600000000001 0 0.00056926 3.3 0.0005691800000000001 3.3 0.00056928 0 0.0005692000000000001 0 0.0005693 3.3 0.0005692200000000001 3.3 0.00056932 0 0.00056924 0 0.00056934 3.3 0.00056926 3.3 0.00056936 0 0.00056928 0 0.00056938 3.3 0.0005693 3.3 0.0005694 0 0.00056932 0 0.00056942 3.3 0.00056934 3.3 0.0005694399999999999 0 0.0005693600000000001 0 0.00056946 3.3 0.0005693800000000001 3.3 0.00056948 0 0.0005694000000000001 0 0.0005695 3.3 0.0005694200000000001 3.3 0.00056952 0 0.00056944 0 0.00056954 3.3 0.00056946 3.3 0.00056956 0 0.00056948 0 0.00056958 3.3 0.0005695 3.3 0.0005696 0 0.00056952 0 0.00056962 3.3 0.00056954 3.3 0.00056964 0 0.00056956 0 0.0005696599999999999 3.3 0.0005695800000000001 3.3 0.00056968 0 0.0005696000000000001 0 0.0005697 3.3 0.0005696200000000001 3.3 0.00056972 0 0.0005696400000000001 0 0.00056974 3.3 0.00056966 3.3 0.00056976 0 0.00056968 0 0.00056978 3.3 0.0005697 3.3 0.0005698 0 0.00056972 0 0.00056982 3.3 0.00056974 3.3 0.00056984 0 0.00056976 0 0.0005698599999999999 3.3 0.0005697800000000001 3.3 0.00056988 0 0.0005698000000000001 0 0.0005699 3.3 0.0005698200000000001 3.3 0.00056992 0 0.0005698400000000001 0 0.00056994 3.3 0.00056986 3.3 0.00056996 0 0.00056988 0 0.00056998 3.3 0.0005699 3.3 0.00057 0 0.00056992 0 0.00057002 3.3 0.00056994 3.3 0.00057004 0 0.00056996 0 0.00057006 3.3 0.00056998 3.3 0.0005700799999999999 0 0.0005700000000000001 0 0.0005701 3.3 0.0005700200000000001 3.3 0.00057012 0 0.0005700400000000001 0 0.00057014 3.3 0.0005700600000000001 3.3 0.00057016 0 0.00057008 0 0.00057018 3.3 0.0005701 3.3 0.0005702 0 0.00057012 0 0.00057022 3.3 0.00057014 3.3 0.00057024 0 0.00057016 0 0.00057026 3.3 0.00057018 3.3 0.0005702799999999999 0 0.0005702000000000001 0 0.0005703 3.3 0.0005702200000000001 3.3 0.00057032 0 0.0005702400000000001 0 0.00057034 3.3 0.0005702600000000001 3.3 0.00057036 0 0.00057028 0 0.00057038 3.3 0.0005703 3.3 0.0005704 0 0.00057032 0 0.00057042 3.3 0.00057034 3.3 0.00057044 0 0.00057036 0 0.00057046 3.3 0.00057038 3.3 0.0005704799999999999 0 0.0005704 0 0.0005704999999999999 3.3 0.0005704200000000001 3.3 0.00057052 0 0.0005704400000000001 0 0.00057054 3.3 0.0005704600000000001 3.3 0.00057056 0 0.00057048 0 0.00057058 3.3 0.0005705 3.3 0.0005706 0 0.00057052 0 0.00057062 3.3 0.00057054 3.3 0.00057064 0 0.00057056 0 0.00057066 3.3 0.00057058 3.3 0.00057068 0 0.0005706 0 0.0005706999999999999 3.3 0.0005706200000000001 3.3 0.00057072 0 0.0005706400000000001 0 0.00057074 3.3 0.0005706600000000001 3.3 0.00057076 0 0.0005706800000000001 0 0.00057078 3.3 0.0005707 3.3 0.0005708 0 0.00057072 0 0.00057082 3.3 0.00057074 3.3 0.00057084 0 0.00057076 0 0.00057086 3.3 0.00057078 3.3 0.00057088 0 0.0005708 0 0.0005708999999999999 3.3 0.00057082 3.3 0.0005709199999999999 0 0.0005708400000000001 0 0.00057094 3.3 0.0005708600000000001 3.3 0.00057096 0 0.0005708800000000001 0 0.00057098 3.3 0.0005709 3.3 0.000571 0 0.00057092 0 0.00057102 3.3 0.00057094 3.3 0.00057104 0 0.00057096 0 0.00057106 3.3 0.00057098 3.3 0.00057108 0 0.000571 0 0.0005711 3.3 0.00057102 3.3 0.0005711199999999999 0 0.0005710400000000001 0 0.00057114 3.3 0.0005710600000000001 3.3 0.00057116 0 0.0005710800000000001 0 0.00057118 3.3 0.0005711000000000001 3.3 0.0005712 0 0.00057112 0 0.00057122 3.3 0.00057114 3.3 0.00057124 0 0.00057116 0 0.00057126 3.3 0.00057118 3.3 0.00057128 0 0.0005712 0 0.0005713 3.3 0.00057122 3.3 0.0005713199999999999 0 0.0005712400000000001 0 0.00057134 3.3 0.0005712600000000001 3.3 0.00057136 0 0.0005712800000000001 0 0.00057138 3.3 0.0005713000000000001 3.3 0.0005714 0 0.00057132 0 0.00057142 3.3 0.00057134 3.3 0.00057144 0 0.00057136 0 0.00057146 3.3 0.00057138 3.3 0.00057148 0 0.0005714 0 0.0005715 3.3 0.00057142 3.3 0.00057152 0 0.00057144 0 0.0005715399999999999 3.3 0.0005714600000000001 3.3 0.00057156 0 0.0005714800000000001 0 0.00057158 3.3 0.0005715000000000001 3.3 0.0005716 0 0.0005715200000000001 0 0.00057162 3.3 0.00057154 3.3 0.00057164 0 0.00057156 0 0.00057166 3.3 0.00057158 3.3 0.00057168 0 0.0005716 0 0.0005717 3.3 0.00057162 3.3 0.00057172 0 0.00057164 0 0.0005717399999999999 3.3 0.0005716600000000001 3.3 0.00057176 0 0.0005716800000000001 0 0.00057178 3.3 0.0005717000000000001 3.3 0.0005718 0 0.0005717200000000001 0 0.00057182 3.3 0.00057174 3.3 0.00057184 0 0.00057176 0 0.00057186 3.3 0.00057178 3.3 0.00057188 0 0.0005718 0 0.0005719 3.3 0.00057182 3.3 0.00057192 0 0.00057184 0 0.00057194 3.3 0.00057186 3.3 0.0005719599999999999 0 0.0005718800000000001 0 0.00057198 3.3 0.0005719000000000001 3.3 0.000572 0 0.0005719200000000001 0 0.00057202 3.3 0.0005719400000000001 3.3 0.00057204 0 0.00057196 0 0.00057206 3.3 0.00057198 3.3 0.00057208 0 0.000572 0 0.0005721 3.3 0.00057202 3.3 0.00057212 0 0.00057204 0 0.00057214 3.3 0.00057206 3.3 0.0005721599999999999 0 0.0005720800000000001 0 0.00057218 3.3 0.0005721000000000001 3.3 0.0005722 0 0.0005721200000000001 0 0.00057222 3.3 0.0005721400000000001 3.3 0.00057224 0 0.00057216 0 0.00057226 3.3 0.00057218 3.3 0.00057228 0 0.0005722 0 0.0005723 3.3 0.00057222 3.3 0.00057232 0 0.00057224 0 0.00057234 3.3 0.00057226 3.3 0.00057236 0 0.00057228 0 0.0005723799999999999 3.3 0.0005723000000000001 3.3 0.0005724 0 0.0005723200000000001 0 0.00057242 3.3 0.0005723400000000001 3.3 0.00057244 0 0.0005723600000000001 0 0.00057246 3.3 0.00057238 3.3 0.00057248 0 0.0005724 0 0.0005725 3.3 0.00057242 3.3 0.00057252 0 0.00057244 0 0.00057254 3.3 0.00057246 3.3 0.00057256 0 0.00057248 0 0.0005725799999999999 3.3 0.0005725000000000001 3.3 0.0005726 0 0.0005725200000000001 0 0.00057262 3.3 0.0005725400000000001 3.3 0.00057264 0 0.0005725600000000001 0 0.00057266 3.3 0.00057258 3.3 0.00057268 0 0.0005726 0 0.0005727 3.3 0.00057262 3.3 0.00057272 0 0.00057264 0 0.00057274 3.3 0.00057266 3.3 0.00057276 0 0.00057268 0 0.00057278 3.3 0.0005727 3.3 0.0005727999999999999 0 0.0005727200000000001 0 0.00057282 3.3 0.0005727400000000001 3.3 0.00057284 0 0.0005727600000000001 0 0.00057286 3.3 0.0005727800000000001 3.3 0.00057288 0 0.0005728 0 0.0005729 3.3 0.00057282 3.3 0.00057292 0 0.00057284 0 0.00057294 3.3 0.00057286 3.3 0.00057296 0 0.00057288 0 0.00057298 3.3 0.0005729 3.3 0.0005729999999999999 0 0.0005729200000000001 0 0.00057302 3.3 0.0005729400000000001 3.3 0.00057304 0 0.0005729600000000001 0 0.00057306 3.3 0.0005729800000000001 3.3 0.00057308 0 0.000573 0 0.0005731 3.3 0.00057302 3.3 0.00057312 0 0.00057304 0 0.00057314 3.3 0.00057306 3.3 0.00057316 0 0.00057308 0 0.00057318 3.3 0.0005731 3.3 0.0005732 0 0.00057312 0 0.0005732199999999999 3.3 0.0005731400000000001 3.3 0.00057324 0 0.0005731600000000001 0 0.00057326 3.3 0.0005731800000000001 3.3 0.00057328 0 0.0005732000000000001 0 0.0005733 3.3 0.00057322 3.3 0.00057332 0 0.00057324 0 0.00057334 3.3 0.00057326 3.3 0.00057336 0 0.00057328 0 0.00057338 3.3 0.0005733 3.3 0.0005734 0 0.00057332 0 0.0005734199999999999 3.3 0.0005733400000000001 3.3 0.00057344 0 0.0005733600000000001 0 0.00057346 3.3 0.0005733800000000001 3.3 0.00057348 0 0.0005734000000000001 0 0.0005735 3.3 0.00057342 3.3 0.00057352 0 0.00057344 0 0.00057354 3.3 0.00057346 3.3 0.00057356 0 0.00057348 0 0.00057358 3.3 0.0005735 3.3 0.0005736 0 0.00057352 0 0.00057362 3.3 0.00057354 3.3 0.0005736399999999999 0 0.0005735600000000001 0 0.00057366 3.3 0.0005735800000000001 3.3 0.00057368 0 0.0005736000000000001 0 0.0005737 3.3 0.0005736200000000001 3.3 0.00057372 0 0.00057364 0 0.00057374 3.3 0.00057366 3.3 0.00057376 0 0.00057368 0 0.00057378 3.3 0.0005737 3.3 0.0005738 0 0.00057372 0 0.00057382 3.3 0.00057374 3.3 0.0005738399999999999 0 0.0005737600000000001 0 0.00057386 3.3 0.0005737800000000001 3.3 0.00057388 0 0.0005738000000000001 0 0.0005739 3.3 0.0005738200000000001 3.3 0.00057392 0 0.00057384 0 0.00057394 3.3 0.00057386 3.3 0.00057396 0 0.00057388 0 0.00057398 3.3 0.0005739 3.3 0.000574 0 0.00057392 0 0.00057402 3.3 0.00057394 3.3 0.0005740399999999999 0 0.00057396 0 0.0005740599999999999 3.3 0.0005739800000000001 3.3 0.00057408 0 0.0005740000000000001 0 0.0005741 3.3 0.0005740200000000001 3.3 0.00057412 0 0.00057404 0 0.00057414 3.3 0.00057406 3.3 0.00057416 0 0.00057408 0 0.00057418 3.3 0.0005741 3.3 0.0005742 0 0.00057412 0 0.00057422 3.3 0.00057414 3.3 0.00057424 0 0.00057416 0 0.0005742599999999999 3.3 0.0005741800000000001 3.3 0.00057428 0 0.0005742000000000001 0 0.0005743 3.3 0.0005742200000000001 3.3 0.00057432 0 0.0005742400000000001 0 0.00057434 3.3 0.00057426 3.3 0.00057436 0 0.00057428 0 0.00057438 3.3 0.0005743 3.3 0.0005744 0 0.00057432 0 0.00057442 3.3 0.00057434 3.3 0.00057444 0 0.00057436 0 0.0005744599999999999 3.3 0.00057438 3.3 0.0005744799999999999 0 0.0005744000000000001 0 0.0005745 3.3 0.0005744200000000001 3.3 0.00057452 0 0.0005744400000000001 0 0.00057454 3.3 0.00057446 3.3 0.00057456 0 0.00057448 0 0.00057458 3.3 0.0005745 3.3 0.0005746 0 0.00057452 0 0.00057462 3.3 0.00057454 3.3 0.00057464 0 0.00057456 0 0.00057466 3.3 0.00057458 3.3 0.0005746799999999999 0 0.0005746000000000001 0 0.0005747 3.3 0.0005746200000000001 3.3 0.00057472 0 0.0005746400000000001 0 0.00057474 3.3 0.0005746600000000001 3.3 0.00057476 0 0.00057468 0 0.00057478 3.3 0.0005747 3.3 0.0005748 0 0.00057472 0 0.00057482 3.3 0.00057474 3.3 0.00057484 0 0.00057476 0 0.00057486 3.3 0.00057478 3.3 0.0005748799999999999 0 0.0005748000000000001 0 0.0005749 3.3 0.0005748200000000001 3.3 0.00057492 0 0.0005748400000000001 0 0.00057494 3.3 0.0005748600000000001 3.3 0.00057496 0 0.00057488 0 0.00057498 3.3 0.0005749 3.3 0.000575 0 0.00057492 0 0.00057502 3.3 0.00057494 3.3 0.00057504 0 0.00057496 0 0.00057506 3.3 0.00057498 3.3 0.00057508 0 0.000575 0 0.0005750999999999999 3.3 0.0005750200000000001 3.3 0.00057512 0 0.0005750400000000001 0 0.00057514 3.3 0.0005750600000000001 3.3 0.00057516 0 0.0005750800000000001 0 0.00057518 3.3 0.0005751 3.3 0.0005752 0 0.00057512 0 0.00057522 3.3 0.00057514 3.3 0.00057524 0 0.00057516 0 0.00057526 3.3 0.00057518 3.3 0.00057528 0 0.0005752 0 0.0005752999999999999 3.3 0.0005752200000000001 3.3 0.00057532 0 0.0005752400000000001 0 0.00057534 3.3 0.0005752600000000001 3.3 0.00057536 0 0.0005752800000000001 0 0.00057538 3.3 0.0005753 3.3 0.0005754 0 0.00057532 0 0.00057542 3.3 0.00057534 3.3 0.00057544 0 0.00057536 0 0.00057546 3.3 0.00057538 3.3 0.00057548 0 0.0005754 0 0.0005755 3.3 0.00057542 3.3 0.0005755199999999999 0 0.0005754400000000001 0 0.00057554 3.3 0.0005754600000000001 3.3 0.00057556 0 0.0005754800000000001 0 0.00057558 3.3 0.0005755000000000001 3.3 0.0005756 0 0.00057552 0 0.00057562 3.3 0.00057554 3.3 0.00057564 0 0.00057556 0 0.00057566 3.3 0.00057558 3.3 0.00057568 0 0.0005756 0 0.0005757 3.3 0.00057562 3.3 0.0005757199999999999 0 0.0005756400000000001 0 0.00057574 3.3 0.0005756600000000001 3.3 0.00057576 0 0.0005756800000000001 0 0.00057578 3.3 0.0005757000000000001 3.3 0.0005758 0 0.00057572 0 0.00057582 3.3 0.00057574 3.3 0.00057584 0 0.00057576 0 0.00057586 3.3 0.00057578 3.3 0.00057588 0 0.0005758 0 0.0005759 3.3 0.00057582 3.3 0.00057592 0 0.00057584 0 0.0005759399999999999 3.3 0.0005758600000000001 3.3 0.00057596 0 0.0005758800000000001 0 0.00057598 3.3 0.0005759000000000001 3.3 0.000576 0 0.0005759200000000001 0 0.00057602 3.3 0.00057594 3.3 0.00057604 0 0.00057596 0 0.00057606 3.3 0.00057598 3.3 0.00057608 0 0.000576 0 0.0005761 3.3 0.00057602 3.3 0.00057612 0 0.00057604 0 0.0005761399999999999 3.3 0.0005760600000000001 3.3 0.00057616 0 0.0005760800000000001 0 0.00057618 3.3 0.0005761000000000001 3.3 0.0005762 0 0.0005761200000000001 0 0.00057622 3.3 0.00057614 3.3 0.00057624 0 0.00057616 0 0.00057626 3.3 0.00057618 3.3 0.00057628 0 0.0005762 0 0.0005763 3.3 0.00057622 3.3 0.00057632 0 0.00057624 0 0.00057634 3.3 0.00057626 3.3 0.0005763599999999999 0 0.0005762800000000001 0 0.00057638 3.3 0.0005763000000000001 3.3 0.0005764 0 0.0005763200000000001 0 0.00057642 3.3 0.0005763400000000001 3.3 0.00057644 0 0.00057636 0 0.00057646 3.3 0.00057638 3.3 0.00057648 0 0.0005764 0 0.0005765 3.3 0.00057642 3.3 0.00057652 0 0.00057644 0 0.00057654 3.3 0.00057646 3.3 0.0005765599999999999 0 0.0005764800000000001 0 0.00057658 3.3 0.0005765000000000001 3.3 0.0005766 0 0.0005765200000000001 0 0.00057662 3.3 0.0005765400000000001 3.3 0.00057664 0 0.00057656 0 0.00057666 3.3 0.00057658 3.3 0.00057668 0 0.0005766 0 0.0005767 3.3 0.00057662 3.3 0.00057672 0 0.00057664 0 0.00057674 3.3 0.00057666 3.3 0.00057676 0 0.00057668 0 0.0005767799999999999 3.3 0.0005767000000000001 3.3 0.0005768 0 0.0005767200000000001 0 0.00057682 3.3 0.0005767400000000001 3.3 0.00057684 0 0.0005767600000000001 0 0.00057686 3.3 0.00057678 3.3 0.00057688 0 0.0005768 0 0.0005769 3.3 0.00057682 3.3 0.00057692 0 0.00057684 0 0.00057694 3.3 0.00057686 3.3 0.00057696 0 0.00057688 0 0.0005769799999999999 3.3 0.0005769000000000001 3.3 0.000577 0 0.0005769200000000001 0 0.00057702 3.3 0.0005769400000000001 3.3 0.00057704 0 0.0005769600000000001 0 0.00057706 3.3 0.00057698 3.3 0.00057708 0 0.000577 0 0.0005771 3.3 0.00057702 3.3 0.00057712 0 0.00057704 0 0.00057714 3.3 0.00057706 3.3 0.00057716 0 0.00057708 0 0.0005771799999999999 3.3 0.0005771 3.3 0.0005771999999999999 0 0.0005771200000000001 0 0.00057722 3.3 0.0005771400000000001 3.3 0.00057724 0 0.0005771600000000001 0 0.00057726 3.3 0.00057718 3.3 0.00057728 0 0.0005772 0 0.0005773 3.3 0.00057722 3.3 0.00057732 0 0.00057724 0 0.00057734 3.3 0.00057726 3.3 0.00057736 0 0.00057728 0 0.00057738 3.3 0.0005773 3.3 0.0005773999999999999 0 0.0005773200000000001 0 0.00057742 3.3 0.0005773400000000001 3.3 0.00057744 0 0.0005773600000000001 0 0.00057746 3.3 0.0005773800000000001 3.3 0.00057748 0 0.0005774 0 0.0005775 3.3 0.00057742 3.3 0.00057752 0 0.00057744 0 0.00057754 3.3 0.00057746 3.3 0.00057756 0 0.00057748 0 0.00057758 3.3 0.0005775 3.3 0.0005775999999999999 0 0.00057752 0 0.0005776199999999999 3.3 0.0005775400000000001 3.3 0.00057764 0 0.0005775600000000001 0 0.00057766 3.3 0.0005775800000000001 3.3 0.00057768 0 0.0005776 0 0.0005777 3.3 0.00057762 3.3 0.00057772 0 0.00057764 0 0.00057774 3.3 0.00057766 3.3 0.00057776 0 0.00057768 0 0.00057778 3.3 0.0005777 3.3 0.0005778 0 0.00057772 0 0.0005778199999999999 3.3 0.0005777400000000001 3.3 0.00057784 0 0.0005777600000000001 0 0.00057786 3.3 0.0005777800000000001 3.3 0.00057788 0 0.0005778000000000001 0 0.0005779 3.3 0.00057782 3.3 0.00057792 0 0.00057784 0 0.00057794 3.3 0.00057786 3.3 0.00057796 0 0.00057788 0 0.00057798 3.3 0.0005779 3.3 0.000578 0 0.00057792 0 0.0005780199999999999 3.3 0.0005779400000000001 3.3 0.00057804 0 0.0005779600000000001 0 0.00057806 3.3 0.0005779800000000001 3.3 0.00057808 0 0.0005780000000000001 0 0.0005781 3.3 0.00057802 3.3 0.00057812 0 0.00057804 0 0.00057814 3.3 0.00057806 3.3 0.00057816 0 0.00057808 0 0.00057818 3.3 0.0005781 3.3 0.0005782 0 0.00057812 0 0.00057822 3.3 0.00057814 3.3 0.0005782399999999999 0 0.0005781600000000001 0 0.00057826 3.3 0.0005781800000000001 3.3 0.00057828 0 0.0005782000000000001 0 0.0005783 3.3 0.0005782200000000001 3.3 0.00057832 0 0.00057824 0 0.00057834 3.3 0.00057826 3.3 0.00057836 0 0.00057828 0 0.00057838 3.3 0.0005783 3.3 0.0005784 0 0.00057832 0 0.00057842 3.3 0.00057834 3.3 0.0005784399999999999 0 0.0005783600000000001 0 0.00057846 3.3 0.0005783800000000001 3.3 0.00057848 0 0.0005784000000000001 0 0.0005785 3.3 0.0005784200000000001 3.3 0.00057852 0 0.00057844 0 0.00057854 3.3 0.00057846 3.3 0.00057856 0 0.00057848 0 0.00057858 3.3 0.0005785 3.3 0.0005786 0 0.00057852 0 0.00057862 3.3 0.00057854 3.3 0.00057864 0 0.00057856 0 0.0005786599999999999 3.3 0.0005785800000000001 3.3 0.00057868 0 0.0005786000000000001 0 0.0005787 3.3 0.0005786200000000001 3.3 0.00057872 0 0.0005786400000000001 0 0.00057874 3.3 0.00057866 3.3 0.00057876 0 0.00057868 0 0.00057878 3.3 0.0005787 3.3 0.0005788 0 0.00057872 0 0.00057882 3.3 0.00057874 3.3 0.00057884 0 0.00057876 0 0.0005788599999999999 3.3 0.0005787800000000001 3.3 0.00057888 0 0.0005788000000000001 0 0.0005789 3.3 0.0005788200000000001 3.3 0.00057892 0 0.0005788400000000001 0 0.00057894 3.3 0.00057886 3.3 0.00057896 0 0.00057888 0 0.00057898 3.3 0.0005789 3.3 0.000579 0 0.00057892 0 0.00057902 3.3 0.00057894 3.3 0.00057904 0 0.00057896 0 0.00057906 3.3 0.00057898 3.3 0.0005790799999999999 0 0.0005790000000000001 0 0.0005791 3.3 0.0005790200000000001 3.3 0.00057912 0 0.0005790400000000001 0 0.00057914 3.3 0.0005790600000000001 3.3 0.00057916 0 0.00057908 0 0.00057918 3.3 0.0005791 3.3 0.0005792 0 0.00057912 0 0.00057922 3.3 0.00057914 3.3 0.00057924 0 0.00057916 0 0.00057926 3.3 0.00057918 3.3 0.0005792799999999999 0 0.0005792000000000001 0 0.0005793 3.3 0.0005792200000000001 3.3 0.00057932 0 0.0005792400000000001 0 0.00057934 3.3 0.0005792600000000001 3.3 0.00057936 0 0.00057928 0 0.00057938 3.3 0.0005793 3.3 0.0005794 0 0.00057932 0 0.00057942 3.3 0.00057934 3.3 0.00057944 0 0.00057936 0 0.00057946 3.3 0.00057938 3.3 0.00057948 0 0.0005794 0 0.0005794999999999999 3.3 0.0005794200000000001 3.3 0.00057952 0 0.0005794400000000001 0 0.00057954 3.3 0.0005794600000000001 3.3 0.00057956 0 0.0005794800000000001 0 0.00057958 3.3 0.0005795 3.3 0.0005796 0 0.00057952 0 0.00057962 3.3 0.00057954 3.3 0.00057964 0 0.00057956 0 0.00057966 3.3 0.00057958 3.3 0.00057968 0 0.0005796 0 0.0005796999999999999 3.3 0.0005796200000000001 3.3 0.00057972 0 0.0005796400000000001 0 0.00057974 3.3 0.0005796600000000001 3.3 0.00057976 0 0.0005796800000000001 0 0.00057978 3.3 0.0005797 3.3 0.0005798 0 0.00057972 0 0.00057982 3.3 0.00057974 3.3 0.00057984 0 0.00057976 0 0.00057986 3.3 0.00057978 3.3 0.00057988 0 0.0005798 0 0.0005799 3.3 0.00057982 3.3 0.0005799199999999999 0 0.0005798400000000001 0 0.00057994 3.3 0.0005798600000000001 3.3 0.00057996 0 0.0005798800000000001 0 0.00057998 3.3 0.0005799000000000001 3.3 0.00058 0 0.00057992 0 0.00058002 3.3 0.00057994 3.3 0.00058004 0 0.00057996 0 0.00058006 3.3 0.00057998 3.3 0.00058008 0 0.00058 0 0.0005801 3.3 0.00058002 3.3 0.0005801199999999999 0 0.0005800400000000001 0 0.00058014 3.3 0.0005800600000000001 3.3 0.00058016 0 0.0005800800000000001 0 0.00058018 3.3 0.0005801000000000001 3.3 0.0005802 0 0.00058012 0 0.00058022 3.3 0.00058014 3.3 0.00058024 0 0.00058016 0 0.00058026 3.3 0.00058018 3.3 0.00058028 0 0.0005802 0 0.0005803 3.3 0.00058022 3.3 0.00058032 0 0.00058024 0 0.0005803399999999999 3.3 0.0005802600000000001 3.3 0.00058036 0 0.0005802800000000001 0 0.00058038 3.3 0.0005803000000000001 3.3 0.0005804 0 0.0005803200000000001 0 0.00058042 3.3 0.00058034 3.3 0.00058044 0 0.00058036 0 0.00058046 3.3 0.00058038 3.3 0.00058048 0 0.0005804 0 0.0005805 3.3 0.00058042 3.3 0.00058052 0 0.00058044 0 0.0005805399999999999 3.3 0.0005804600000000001 3.3 0.00058056 0 0.0005804800000000001 0 0.00058058 3.3 0.0005805000000000001 3.3 0.0005806 0 0.0005805200000000001 0 0.00058062 3.3 0.00058054 3.3 0.00058064 0 0.00058056 0 0.00058066 3.3 0.00058058 3.3 0.00058068 0 0.0005806 0 0.0005807 3.3 0.00058062 3.3 0.00058072 0 0.00058064 0 0.0005807399999999999 3.3 0.00058066 3.3 0.0005807599999999999 0 0.0005806800000000001 0 0.00058078 3.3 0.0005807000000000001 3.3 0.0005808 0 0.0005807200000000001 0 0.00058082 3.3 0.00058074 3.3 0.00058084 0 0.00058076 0 0.00058086 3.3 0.00058078 3.3 0.00058088 0 0.0005808 0 0.0005809 3.3 0.00058082 3.3 0.00058092 0 0.00058084 0 0.00058094 3.3 0.00058086 3.3 0.0005809599999999999 0 0.0005808800000000001 0 0.00058098 3.3 0.0005809000000000001 3.3 0.000581 0 0.0005809200000000001 0 0.00058102 3.3 0.0005809400000000001 3.3 0.00058104 0 0.00058096 0 0.00058106 3.3 0.00058098 3.3 0.00058108 0 0.000581 0 0.0005811 3.3 0.00058102 3.3 0.00058112 0 0.00058104 0 0.00058114 3.3 0.00058106 3.3 0.0005811599999999999 0 0.00058108 0 0.0005811799999999999 3.3 0.0005811000000000001 3.3 0.0005812 0 0.0005811200000000001 0 0.00058122 3.3 0.0005811400000000001 3.3 0.00058124 0 0.00058116 0 0.00058126 3.3 0.00058118 3.3 0.00058128 0 0.0005812 0 0.0005813 3.3 0.00058122 3.3 0.00058132 0 0.00058124 0 0.00058134 3.3 0.00058126 3.3 0.00058136 0 0.00058128 0 0.0005813799999999999 3.3 0.0005813000000000001 3.3 0.0005814 0 0.0005813200000000001 0 0.00058142 3.3 0.0005813400000000001 3.3 0.00058144 0 0.0005813600000000001 0 0.00058146 3.3 0.00058138 3.3 0.00058148 0 0.0005814 0 0.0005815 3.3 0.00058142 3.3 0.00058152 0 0.00058144 0 0.00058154 3.3 0.00058146 3.3 0.00058156 0 0.00058148 0 0.0005815799999999999 3.3 0.0005815000000000001 3.3 0.0005816 0 0.0005815200000000001 0 0.00058162 3.3 0.0005815400000000001 3.3 0.00058164 0 0.0005815600000000001 0 0.00058166 3.3 0.00058158 3.3 0.00058168 0 0.0005816 0 0.0005817 3.3 0.00058162 3.3 0.00058172 0 0.00058164 0 0.00058174 3.3 0.00058166 3.3 0.00058176 0 0.00058168 0 0.00058178 3.3 0.0005817 3.3 0.0005817999999999999 0 0.0005817200000000001 0 0.00058182 3.3 0.0005817400000000001 3.3 0.00058184 0 0.0005817600000000001 0 0.00058186 3.3 0.0005817800000000001 3.3 0.00058188 0 0.0005818 0 0.0005819 3.3 0.00058182 3.3 0.00058192 0 0.00058184 0 0.00058194 3.3 0.00058186 3.3 0.00058196 0 0.00058188 0 0.00058198 3.3 0.0005819 3.3 0.0005819999999999999 0 0.0005819200000000001 0 0.00058202 3.3 0.0005819400000000001 3.3 0.00058204 0 0.0005819600000000001 0 0.00058206 3.3 0.0005819800000000001 3.3 0.00058208 0 0.000582 0 0.0005821 3.3 0.00058202 3.3 0.00058212 0 0.00058204 0 0.00058214 3.3 0.00058206 3.3 0.00058216 0 0.00058208 0 0.00058218 3.3 0.0005821 3.3 0.0005822 0 0.00058212 0 0.0005822199999999999 3.3 0.0005821400000000001 3.3 0.00058224 0 0.0005821600000000001 0 0.00058226 3.3 0.0005821800000000001 3.3 0.00058228 0 0.0005822000000000001 0 0.0005823 3.3 0.00058222 3.3 0.00058232 0 0.00058224 0 0.00058234 3.3 0.00058226 3.3 0.00058236 0 0.00058228 0 0.00058238 3.3 0.0005823 3.3 0.0005824 0 0.00058232 0 0.0005824199999999999 3.3 0.0005823400000000001 3.3 0.00058244 0 0.0005823600000000001 0 0.00058246 3.3 0.0005823800000000001 3.3 0.00058248 0 0.0005824000000000001 0 0.0005825 3.3 0.00058242 3.3 0.00058252 0 0.00058244 0 0.00058254 3.3 0.00058246 3.3 0.00058256 0 0.00058248 0 0.00058258 3.3 0.0005825 3.3 0.0005826 0 0.00058252 0 0.00058262 3.3 0.00058254 3.3 0.0005826399999999999 0 0.0005825600000000001 0 0.00058266 3.3 0.0005825800000000001 3.3 0.00058268 0 0.0005826000000000001 0 0.0005827 3.3 0.0005826200000000001 3.3 0.00058272 0 0.00058264 0 0.00058274 3.3 0.00058266 3.3 0.00058276 0 0.00058268 0 0.00058278 3.3 0.0005827 3.3 0.0005828 0 0.00058272 0 0.00058282 3.3 0.00058274 3.3 0.0005828399999999999 0 0.0005827600000000001 0 0.00058286 3.3 0.0005827800000000001 3.3 0.00058288 0 0.0005828000000000001 0 0.0005829 3.3 0.0005828200000000001 3.3 0.00058292 0 0.00058284 0 0.00058294 3.3 0.00058286 3.3 0.00058296 0 0.00058288 0 0.00058298 3.3 0.0005829 3.3 0.000583 0 0.00058292 0 0.00058302 3.3 0.00058294 3.3 0.00058304 0 0.00058296 0 0.0005830599999999999 3.3 0.0005829800000000001 3.3 0.00058308 0 0.0005830000000000001 0 0.0005831 3.3 0.0005830200000000001 3.3 0.00058312 0 0.0005830400000000001 0 0.00058314 3.3 0.00058306 3.3 0.00058316 0 0.00058308 0 0.00058318 3.3 0.0005831 3.3 0.0005832 0 0.00058312 0 0.00058322 3.3 0.00058314 3.3 0.00058324 0 0.00058316 0 0.0005832599999999999 3.3 0.0005831800000000001 3.3 0.00058328 0 0.0005832000000000001 0 0.0005833 3.3 0.0005832200000000001 3.3 0.00058332 0 0.0005832400000000001 0 0.00058334 3.3 0.00058326 3.3 0.00058336 0 0.00058328 0 0.00058338 3.3 0.0005833 3.3 0.0005834 0 0.00058332 0 0.00058342 3.3 0.00058334 3.3 0.00058344 0 0.00058336 0 0.00058346 3.3 0.00058338 3.3 0.0005834799999999999 0 0.0005834000000000001 0 0.0005835 3.3 0.0005834200000000001 3.3 0.00058352 0 0.0005834400000000001 0 0.00058354 3.3 0.0005834600000000001 3.3 0.00058356 0 0.00058348 0 0.00058358 3.3 0.0005835 3.3 0.0005836 0 0.00058352 0 0.00058362 3.3 0.00058354 3.3 0.00058364 0 0.00058356 0 0.00058366 3.3 0.00058358 3.3 0.0005836799999999999 0 0.0005836000000000001 0 0.0005837 3.3 0.0005836200000000001 3.3 0.00058372 0 0.0005836400000000001 0 0.00058374 3.3 0.0005836600000000001 3.3 0.00058376 0 0.00058368 0 0.00058378 3.3 0.0005837 3.3 0.0005838 0 0.00058372 0 0.00058382 3.3 0.00058374 3.3 0.00058384 0 0.00058376 0 0.00058386 3.3 0.00058378 3.3 0.00058388 0 0.0005838 0 0.0005838999999999999 3.3 0.0005838200000000001 3.3 0.00058392 0 0.0005838400000000001 0 0.00058394 3.3 0.0005838600000000001 3.3 0.00058396 0 0.0005838800000000001 0 0.00058398 3.3 0.0005839 3.3 0.000584 0 0.00058392 0 0.00058402 3.3 0.00058394 3.3 0.00058404 0 0.00058396 0 0.00058406 3.3 0.00058398 3.3 0.00058408 0 0.000584 0 0.0005840999999999999 3.3 0.0005840200000000001 3.3 0.00058412 0 0.0005840400000000001 0 0.00058414 3.3 0.0005840600000000001 3.3 0.00058416 0 0.0005840800000000001 0 0.00058418 3.3 0.0005841 3.3 0.0005842 0 0.00058412 0 0.00058422 3.3 0.00058414 3.3 0.00058424 0 0.00058416 0 0.00058426 3.3 0.00058418 3.3 0.00058428 0 0.0005842 0 0.0005842999999999999 3.3 0.00058422 3.3 0.0005843199999999999 0 0.0005842400000000001 0 0.00058434 3.3 0.0005842600000000001 3.3 0.00058436 0 0.0005842800000000001 0 0.00058438 3.3 0.0005843 3.3 0.0005844 0 0.00058432 0 0.00058442 3.3 0.00058434 3.3 0.00058444 0 0.00058436 0 0.00058446 3.3 0.00058438 3.3 0.00058448 0 0.0005844 0 0.0005845 3.3 0.00058442 3.3 0.0005845199999999999 0 0.0005844400000000001 0 0.00058454 3.3 0.0005844600000000001 3.3 0.00058456 0 0.0005844800000000001 0 0.00058458 3.3 0.0005845000000000001 3.3 0.0005846 0 0.00058452 0 0.00058462 3.3 0.00058454 3.3 0.00058464 0 0.00058456 0 0.00058466 3.3 0.00058458 3.3 0.00058468 0 0.0005846 0 0.0005847 3.3 0.00058462 3.3 0.0005847199999999999 0 0.00058464 0 0.0005847399999999999 3.3 0.0005846600000000001 3.3 0.00058476 0 0.0005846800000000001 0 0.00058478 3.3 0.0005847000000000001 3.3 0.0005848 0 0.00058472 0 0.00058482 3.3 0.00058474 3.3 0.00058484 0 0.00058476 0 0.00058486 3.3 0.00058478 3.3 0.00058488 0 0.0005848 0 0.0005849 3.3 0.00058482 3.3 0.00058492 0 0.00058484 0 0.0005849399999999999 3.3 0.0005848600000000001 3.3 0.00058496 0 0.0005848800000000001 0 0.00058498 3.3 0.0005849000000000001 3.3 0.000585 0 0.0005849200000000001 0 0.00058502 3.3 0.00058494 3.3 0.00058504 0 0.00058496 0 0.00058506 3.3 0.00058498 3.3 0.00058508 0 0.000585 0 0.0005851 3.3 0.00058502 3.3 0.00058512 0 0.00058504 0 0.0005851399999999999 3.3 0.0005850600000000001 3.3 0.00058516 0 0.0005850800000000001 0 0.00058518 3.3 0.0005851000000000001 3.3 0.0005852 0 0.0005851200000000001 0 0.00058522 3.3 0.00058514 3.3 0.00058524 0 0.00058516 0 0.00058526 3.3 0.00058518 3.3 0.00058528 0 0.0005852 0 0.0005853 3.3 0.00058522 3.3 0.00058532 0 0.00058524 0 0.00058534 3.3 0.00058526 3.3 0.0005853599999999999 0 0.0005852800000000001 0 0.00058538 3.3 0.0005853000000000001 3.3 0.0005854 0 0.0005853200000000001 0 0.00058542 3.3 0.0005853400000000001 3.3 0.00058544 0 0.00058536 0 0.00058546 3.3 0.00058538 3.3 0.00058548 0 0.0005854 0 0.0005855 3.3 0.00058542 3.3 0.00058552 0 0.00058544 0 0.00058554 3.3 0.00058546 3.3 0.0005855599999999999 0 0.0005854800000000001 0 0.00058558 3.3 0.0005855000000000001 3.3 0.0005856 0 0.0005855200000000001 0 0.00058562 3.3 0.0005855400000000001 3.3 0.00058564 0 0.00058556 0 0.00058566 3.3 0.00058558 3.3 0.00058568 0 0.0005856 0 0.0005857 3.3 0.00058562 3.3 0.00058572 0 0.00058564 0 0.00058574 3.3 0.00058566 3.3 0.00058576 0 0.00058568 0 0.0005857799999999999 3.3 0.0005857000000000001 3.3 0.0005858 0 0.0005857200000000001 0 0.00058582 3.3 0.0005857400000000001 3.3 0.00058584 0 0.0005857600000000001 0 0.00058586 3.3 0.00058578 3.3 0.00058588 0 0.0005858 0 0.0005859 3.3 0.00058582 3.3 0.00058592 0 0.00058584 0 0.00058594 3.3 0.00058586 3.3 0.00058596 0 0.00058588 0 0.0005859799999999999 3.3 0.0005859000000000001 3.3 0.000586 0 0.0005859200000000001 0 0.00058602 3.3 0.0005859400000000001 3.3 0.00058604 0 0.0005859600000000001 0 0.00058606 3.3 0.00058598 3.3 0.00058608 0 0.000586 0 0.0005861 3.3 0.00058602 3.3 0.00058612 0 0.00058604 0 0.00058614 3.3 0.00058606 3.3 0.00058616 0 0.00058608 0 0.00058618 3.3 0.0005861 3.3 0.0005861999999999999 0 0.0005861200000000001 0 0.00058622 3.3 0.0005861400000000001 3.3 0.00058624 0 0.0005861600000000001 0 0.00058626 3.3 0.0005861800000000001 3.3 0.00058628 0 0.0005862 0 0.0005863 3.3 0.00058622 3.3 0.00058632 0 0.00058624 0 0.00058634 3.3 0.00058626 3.3 0.00058636 0 0.00058628 0 0.00058638 3.3 0.0005863 3.3 0.0005863999999999999 0 0.0005863200000000001 0 0.00058642 3.3 0.0005863400000000001 3.3 0.00058644 0 0.0005863600000000001 0 0.00058646 3.3 0.0005863800000000001 3.3 0.00058648 0 0.0005864 0 0.0005865 3.3 0.00058642 3.3 0.00058652 0 0.00058644 0 0.00058654 3.3 0.00058646 3.3 0.00058656 0 0.00058648 0 0.00058658 3.3 0.0005865 3.3 0.0005866 0 0.00058652 0 0.0005866199999999999 3.3 0.0005865400000000001 3.3 0.00058664 0 0.0005865600000000001 0 0.00058666 3.3 0.0005865800000000001 3.3 0.00058668 0 0.0005866000000000001 0 0.0005867 3.3 0.00058662 3.3 0.00058672 0 0.00058664 0 0.00058674 3.3 0.00058666 3.3 0.00058676 0 0.00058668 0 0.00058678 3.3 0.0005867 3.3 0.0005868 0 0.00058672 0 0.0005868199999999999 3.3 0.0005867400000000001 3.3 0.00058684 0 0.0005867600000000001 0 0.00058686 3.3 0.0005867800000000001 3.3 0.00058688 0 0.0005868000000000001 0 0.0005869 3.3 0.00058682 3.3 0.00058692 0 0.00058684 0 0.00058694 3.3 0.00058686 3.3 0.00058696 0 0.00058688 0 0.00058698 3.3 0.0005869 3.3 0.000587 0 0.00058692 0 0.00058702 3.3 0.00058694 3.3 0.0005870399999999999 0 0.0005869600000000001 0 0.00058706 3.3 0.0005869800000000001 3.3 0.00058708 0 0.0005870000000000001 0 0.0005871 3.3 0.0005870200000000001 3.3 0.00058712 0 0.00058704 0 0.00058714 3.3 0.00058706 3.3 0.00058716 0 0.00058708 0 0.00058718 3.3 0.0005871 3.3 0.0005872 0 0.00058712 0 0.00058722 3.3 0.00058714 3.3 0.0005872399999999999 0 0.0005871600000000001 0 0.00058726 3.3 0.0005871800000000001 3.3 0.00058728 0 0.0005872000000000001 0 0.0005873 3.3 0.0005872200000000001 3.3 0.00058732 0 0.00058724 0 0.00058734 3.3 0.00058726 3.3 0.00058736 0 0.00058728 0 0.00058738 3.3 0.0005873 3.3 0.0005874 0 0.00058732 0 0.00058742 3.3 0.00058734 3.3 0.0005874399999999999 0 0.00058736 0 0.0005874599999999999 3.3 0.0005873800000000001 3.3 0.00058748 0 0.0005874000000000001 0 0.0005875 3.3 0.0005874200000000001 3.3 0.00058752 0 0.00058744 0 0.00058754 3.3 0.00058746 3.3 0.00058756 0 0.00058748 0 0.00058758 3.3 0.0005875 3.3 0.0005876 0 0.00058752 0 0.00058762 3.3 0.00058754 3.3 0.00058764 0 0.00058756 0 0.0005876599999999999 3.3 0.0005875800000000001 3.3 0.00058768 0 0.0005876000000000001 0 0.0005877 3.3 0.0005876200000000001 3.3 0.00058772 0 0.0005876400000000001 0 0.00058774 3.3 0.00058766 3.3 0.00058776 0 0.00058768 0 0.00058778 3.3 0.0005877 3.3 0.0005878 0 0.00058772 0 0.00058782 3.3 0.00058774 3.3 0.00058784 0 0.00058776 0 0.0005878599999999999 3.3 0.00058778 3.3 0.0005878799999999999 0 0.0005878000000000001 0 0.0005879 3.3 0.0005878200000000001 3.3 0.00058792 0 0.0005878400000000001 0 0.00058794 3.3 0.00058786 3.3 0.00058796 0 0.00058788 0 0.00058798 3.3 0.0005879 3.3 0.000588 0 0.00058792 0 0.00058802 3.3 0.00058794 3.3 0.00058804 0 0.00058796 0 0.00058806 3.3 0.00058798 3.3 0.0005880799999999999 0 0.0005880000000000001 0 0.0005881 3.3 0.0005880200000000001 3.3 0.00058812 0 0.0005880400000000001 0 0.00058814 3.3 0.0005880600000000001 3.3 0.00058816 0 0.00058808 0 0.00058818 3.3 0.0005881 3.3 0.0005882 0 0.00058812 0 0.00058822 3.3 0.00058814 3.3 0.00058824 0 0.00058816 0 0.00058826 3.3 0.00058818 3.3 0.0005882799999999999 0 0.0005882 0 0.0005882999999999999 3.3 0.0005882200000000001 3.3 0.00058832 0 0.0005882400000000001 0 0.00058834 3.3 0.0005882600000000001 3.3 0.00058836 0 0.00058828 0 0.00058838 3.3 0.0005883 3.3 0.0005884 0 0.00058832 0 0.00058842 3.3 0.00058834 3.3 0.00058844 0 0.00058836 0 0.00058846 3.3 0.00058838 3.3 0.00058848 0 0.0005884 0 0.0005884999999999999 3.3 0.0005884200000000001 3.3 0.00058852 0 0.0005884400000000001 0 0.00058854 3.3 0.0005884600000000001 3.3 0.00058856 0 0.0005884800000000001 0 0.00058858 3.3 0.0005885 3.3 0.0005886 0 0.00058852 0 0.00058862 3.3 0.00058854 3.3 0.00058864 0 0.00058856 0 0.00058866 3.3 0.00058858 3.3 0.00058868 0 0.0005886 0 0.0005886999999999999 3.3 0.0005886200000000001 3.3 0.00058872 0 0.0005886400000000001 0 0.00058874 3.3 0.0005886600000000001 3.3 0.00058876 0 0.0005886800000000001 0 0.00058878 3.3 0.0005887 3.3 0.0005888 0 0.00058872 0 0.00058882 3.3 0.00058874 3.3 0.00058884 0 0.00058876 0 0.00058886 3.3 0.00058878 3.3 0.00058888 0 0.0005888 0 0.0005889 3.3 0.00058882 3.3 0.0005889199999999999 0 0.0005888400000000001 0 0.00058894 3.3 0.0005888600000000001 3.3 0.00058896 0 0.0005888800000000001 0 0.00058898 3.3 0.0005889000000000001 3.3 0.000589 0 0.00058892 0 0.00058902 3.3 0.00058894 3.3 0.00058904 0 0.00058896 0 0.00058906 3.3 0.00058898 3.3 0.00058908 0 0.000589 0 0.0005891 3.3 0.00058902 3.3 0.0005891199999999999 0 0.0005890400000000001 0 0.00058914 3.3 0.0005890600000000001 3.3 0.00058916 0 0.0005890800000000001 0 0.00058918 3.3 0.0005891000000000001 3.3 0.0005892 0 0.00058912 0 0.00058922 3.3 0.00058914 3.3 0.00058924 0 0.00058916 0 0.00058926 3.3 0.00058918 3.3 0.00058928 0 0.0005892 0 0.0005893 3.3 0.00058922 3.3 0.00058932 0 0.00058924 0 0.0005893399999999999 3.3 0.0005892600000000001 3.3 0.00058936 0 0.0005892800000000001 0 0.00058938 3.3 0.0005893000000000001 3.3 0.0005894 0 0.0005893200000000001 0 0.00058942 3.3 0.00058934 3.3 0.00058944 0 0.00058936 0 0.00058946 3.3 0.00058938 3.3 0.00058948 0 0.0005894 0 0.0005895 3.3 0.00058942 3.3 0.00058952 0 0.00058944 0 0.0005895399999999999 3.3 0.0005894600000000001 3.3 0.00058956 0 0.0005894800000000001 0 0.00058958 3.3 0.0005895000000000001 3.3 0.0005896 0 0.0005895200000000001 0 0.00058962 3.3 0.00058954 3.3 0.00058964 0 0.00058956 0 0.00058966 3.3 0.00058958 3.3 0.00058968 0 0.0005896 0 0.0005897 3.3 0.00058962 3.3 0.00058972 0 0.00058964 0 0.00058974 3.3 0.00058966 3.3 0.0005897599999999999 0 0.0005896800000000001 0 0.00058978 3.3 0.0005897000000000001 3.3 0.0005898 0 0.0005897200000000001 0 0.00058982 3.3 0.0005897400000000001 3.3 0.00058984 0 0.00058976 0 0.00058986 3.3 0.00058978 3.3 0.00058988 0 0.0005898 0 0.0005899 3.3 0.00058982 3.3 0.00058992 0 0.00058984 0 0.00058994 3.3 0.00058986 3.3 0.0005899599999999999 0 0.0005898800000000001 0 0.00058998 3.3 0.0005899000000000001 3.3 0.00059 0 0.0005899200000000001 0 0.00059002 3.3 0.0005899400000000001 3.3 0.00059004 0 0.00058996 0 0.00059006 3.3 0.00058998 3.3 0.00059008 0 0.00059 0 0.0005901 3.3 0.00059002 3.3 0.00059012 0 0.00059004 0 0.00059014 3.3 0.00059006 3.3 0.00059016 0 0.00059008 0 0.0005901799999999999 3.3 0.0005901000000000001 3.3 0.0005902 0 0.0005901200000000001 0 0.00059022 3.3 0.0005901400000000001 3.3 0.00059024 0 0.0005901600000000001 0 0.00059026 3.3 0.00059018 3.3 0.00059028 0 0.0005902 0 0.0005903 3.3 0.00059022 3.3 0.00059032 0 0.00059024 0 0.00059034 3.3 0.00059026 3.3 0.00059036 0 0.00059028 0 0.0005903799999999999 3.3 0.0005903000000000001 3.3 0.0005904 0 0.0005903200000000001 0 0.00059042 3.3 0.0005903400000000001 3.3 0.00059044 0 0.0005903600000000001 0 0.00059046 3.3 0.00059038 3.3 0.00059048 0 0.0005904 0 0.0005905 3.3 0.00059042 3.3 0.00059052 0 0.00059044 0 0.00059054 3.3 0.00059046 3.3 0.00059056 0 0.00059048 0 0.00059058 3.3 0.0005905 3.3 0.0005905999999999999 0 0.0005905200000000001 0 0.00059062 3.3 0.0005905400000000001 3.3 0.00059064 0 0.0005905600000000001 0 0.00059066 3.3 0.0005905800000000001 3.3 0.00059068 0 0.0005906 0 0.0005907 3.3 0.00059062 3.3 0.00059072 0 0.00059064 0 0.00059074 3.3 0.00059066 3.3 0.00059076 0 0.00059068 0 0.00059078 3.3 0.0005907 3.3 0.0005907999999999999 0 0.0005907200000000001 0 0.00059082 3.3 0.0005907400000000001 3.3 0.00059084 0 0.0005907600000000001 0 0.00059086 3.3 0.0005907800000000001 3.3 0.00059088 0 0.0005908 0 0.0005909 3.3 0.00059082 3.3 0.00059092 0 0.00059084 0 0.00059094 3.3 0.00059086 3.3 0.00059096 0 0.00059088 0 0.00059098 3.3 0.0005909 3.3 0.0005909999999999999 0 0.00059092 0 0.0005910199999999999 3.3 0.0005909400000000001 3.3 0.00059104 0 0.0005909600000000001 0 0.00059106 3.3 0.0005909800000000001 3.3 0.00059108 0 0.000591 0 0.0005911 3.3 0.00059102 3.3 0.00059112 0 0.00059104 0 0.00059114 3.3 0.00059106 3.3 0.00059116 0 0.00059108 0 0.00059118 3.3 0.0005911 3.3 0.0005912 0 0.00059112 0 0.0005912199999999999 3.3 0.0005911400000000001 3.3 0.00059124 0 0.0005911600000000001 0 0.00059126 3.3 0.0005911800000000001 3.3 0.00059128 0 0.0005912000000000001 0 0.0005913 3.3 0.00059122 3.3 0.00059132 0 0.00059124 0 0.00059134 3.3 0.00059126 3.3 0.00059136 0 0.00059128 0 0.00059138 3.3 0.0005913 3.3 0.0005914 0 0.00059132 0 0.0005914199999999999 3.3 0.00059134 3.3 0.0005914399999999999 0 0.0005913600000000001 0 0.00059146 3.3 0.0005913800000000001 3.3 0.00059148 0 0.0005914000000000001 0 0.0005915 3.3 0.00059142 3.3 0.00059152 0 0.00059144 0 0.00059154 3.3 0.00059146 3.3 0.00059156 0 0.00059148 0 0.00059158 3.3 0.0005915 3.3 0.0005916 0 0.00059152 0 0.00059162 3.3 0.00059154 3.3 0.0005916399999999999 0 0.0005915600000000001 0 0.00059166 3.3 0.0005915800000000001 3.3 0.00059168 0 0.0005916000000000001 0 0.0005917 3.3 0.0005916200000000001 3.3 0.00059172 0 0.00059164 0 0.00059174 3.3 0.00059166 3.3 0.00059176 0 0.00059168 0 0.00059178 3.3 0.0005917 3.3 0.0005918 0 0.00059172 0 0.00059182 3.3 0.00059174 3.3 0.0005918399999999999 0 0.00059176 0 0.0005918599999999999 3.3 0.0005917800000000001 3.3 0.00059188 0 0.0005918000000000001 0 0.0005919 3.3 0.0005918200000000001 3.3 0.00059192 0 0.00059184 0 0.00059194 3.3 0.00059186 3.3 0.00059196 0 0.00059188 0 0.00059198 3.3 0.0005919 3.3 0.000592 0 0.00059192 0 0.00059202 3.3 0.00059194 3.3 0.00059204 0 0.00059196 0 0.0005920599999999999 3.3 0.0005919800000000001 3.3 0.00059208 0 0.0005920000000000001 0 0.0005921 3.3 0.0005920200000000001 3.3 0.00059212 0 0.0005920400000000001 0 0.00059214 3.3 0.00059206 3.3 0.00059216 0 0.00059208 0 0.00059218 3.3 0.0005921 3.3 0.0005922 0 0.00059212 0 0.00059222 3.3 0.00059214 3.3 0.00059224 0 0.00059216 0 0.0005922599999999999 3.3 0.0005921800000000001 3.3 0.00059228 0 0.0005922000000000001 0 0.0005923 3.3 0.0005922200000000001 3.3 0.00059232 0 0.0005922400000000001 0 0.00059234 3.3 0.00059226 3.3 0.00059236 0 0.00059228 0 0.00059238 3.3 0.0005923 3.3 0.0005924 0 0.00059232 0 0.00059242 3.3 0.00059234 3.3 0.00059244 0 0.00059236 0 0.00059246 3.3 0.00059238 3.3 0.0005924799999999999 0 0.0005924000000000001 0 0.0005925 3.3 0.0005924200000000001 3.3 0.00059252 0 0.0005924400000000001 0 0.00059254 3.3 0.0005924600000000001 3.3 0.00059256 0 0.00059248 0 0.00059258 3.3 0.0005925 3.3 0.0005926 0 0.00059252 0 0.00059262 3.3 0.00059254 3.3 0.00059264 0 0.00059256 0 0.00059266 3.3 0.00059258 3.3 0.0005926799999999999 0 0.0005926000000000001 0 0.0005927 3.3 0.0005926200000000001 3.3 0.00059272 0 0.0005926400000000001 0 0.00059274 3.3 0.0005926600000000001 3.3 0.00059276 0 0.00059268 0 0.00059278 3.3 0.0005927 3.3 0.0005928 0 0.00059272 0 0.00059282 3.3 0.00059274 3.3 0.00059284 0 0.00059276 0 0.00059286 3.3 0.00059278 3.3 0.00059288 0 0.0005928 0 0.0005928999999999999 3.3 0.0005928200000000001 3.3 0.00059292 0 0.0005928400000000001 0 0.00059294 3.3 0.0005928600000000001 3.3 0.00059296 0 0.0005928800000000001 0 0.00059298 3.3 0.0005929 3.3 0.000593 0 0.00059292 0 0.00059302 3.3 0.00059294 3.3 0.00059304 0 0.00059296 0 0.00059306 3.3 0.00059298 3.3 0.00059308 0 0.000593 0 0.0005930999999999999 3.3 0.0005930200000000001 3.3 0.00059312 0 0.0005930400000000001 0 0.00059314 3.3 0.0005930600000000001 3.3 0.00059316 0 0.0005930800000000001 0 0.00059318 3.3 0.0005931 3.3 0.0005932 0 0.00059312 0 0.00059322 3.3 0.00059314 3.3 0.00059324 0 0.00059316 0 0.00059326 3.3 0.00059318 3.3 0.00059328 0 0.0005932 0 0.0005933 3.3 0.00059322 3.3 0.0005933199999999999 0 0.0005932400000000001 0 0.00059334 3.3 0.0005932600000000001 3.3 0.00059336 0 0.0005932800000000001 0 0.00059338 3.3 0.0005933000000000001 3.3 0.0005934 0 0.00059332 0 0.00059342 3.3 0.00059334 3.3 0.00059344 0 0.00059336 0 0.00059346 3.3 0.00059338 3.3 0.00059348 0 0.0005934 0 0.0005935 3.3 0.00059342 3.3 0.0005935199999999999 0 0.0005934400000000001 0 0.00059354 3.3 0.0005934600000000001 3.3 0.00059356 0 0.0005934800000000001 0 0.00059358 3.3 0.0005935000000000001 3.3 0.0005936 0 0.00059352 0 0.00059362 3.3 0.00059354 3.3 0.00059364 0 0.00059356 0 0.00059366 3.3 0.00059358 3.3 0.00059368 0 0.0005936 0 0.0005937 3.3 0.00059362 3.3 0.00059372 0 0.00059364 0 0.0005937399999999999 3.3 0.0005936600000000001 3.3 0.00059376 0 0.0005936800000000001 0 0.00059378 3.3 0.0005937000000000001 3.3 0.0005938 0 0.0005937200000000001 0 0.00059382 3.3 0.00059374 3.3 0.00059384 0 0.00059376 0 0.00059386 3.3 0.00059378 3.3 0.00059388 0 0.0005938 0 0.0005939 3.3 0.00059382 3.3 0.00059392 0 0.00059384 0 0.0005939399999999999 3.3 0.0005938600000000001 3.3 0.00059396 0 0.0005938800000000001 0 0.00059398 3.3 0.0005939000000000001 3.3 0.000594 0 0.0005939200000000001 0 0.00059402 3.3 0.00059394 3.3 0.00059404 0 0.00059396 0 0.00059406 3.3 0.00059398 3.3 0.00059408 0 0.000594 0 0.0005941 3.3 0.00059402 3.3 0.00059412 0 0.00059404 0 0.00059414 3.3 0.00059406 3.3 0.0005941599999999999 0 0.0005940800000000001 0 0.00059418 3.3 0.0005941000000000001 3.3 0.0005942 0 0.0005941200000000001 0 0.00059422 3.3 0.0005941400000000001 3.3 0.00059424 0 0.00059416 0 0.00059426 3.3 0.00059418 3.3 0.00059428 0 0.0005942 0 0.0005943 3.3 0.00059422 3.3 0.00059432 0 0.00059424 0 0.00059434 3.3 0.00059426 3.3 0.0005943599999999999 0 0.0005942800000000001 0 0.00059438 3.3 0.0005943000000000001 3.3 0.0005944 0 0.0005943200000000001 0 0.00059442 3.3 0.0005943400000000001 3.3 0.00059444 0 0.00059436 0 0.00059446 3.3 0.00059438 3.3 0.00059448 0 0.0005944 0 0.0005945 3.3 0.00059442 3.3 0.00059452 0 0.00059444 0 0.00059454 3.3 0.00059446 3.3 0.0005945599999999999 0 0.00059448 0 0.0005945799999999999 3.3 0.0005945000000000001 3.3 0.0005946 0 0.0005945200000000001 0 0.00059462 3.3 0.0005945400000000001 3.3 0.00059464 0 0.00059456 0 0.00059466 3.3 0.00059458 3.3 0.00059468 0 0.0005946 0 0.0005947 3.3 0.00059462 3.3 0.00059472 0 0.00059464 0 0.00059474 3.3 0.00059466 3.3 0.00059476 0 0.00059468 0 0.0005947799999999999 3.3 0.0005947000000000001 3.3 0.0005948 0 0.0005947200000000001 0 0.00059482 3.3 0.0005947400000000001 3.3 0.00059484 0 0.0005947600000000001 0 0.00059486 3.3 0.00059478 3.3 0.00059488 0 0.0005948 0 0.0005949 3.3 0.00059482 3.3 0.00059492 0 0.00059484 0 0.00059494 3.3 0.00059486 3.3 0.00059496 0 0.00059488 0 0.0005949799999999999 3.3 0.0005949 3.3 0.0005949999999999999 0 0.0005949200000000001 0 0.00059502 3.3 0.0005949400000000001 3.3 0.00059504 0 0.0005949600000000001 0 0.00059506 3.3 0.00059498 3.3 0.00059508 0 0.000595 0 0.0005951 3.3 0.00059502 3.3 0.00059512 0 0.00059504 0 0.00059514 3.3 0.00059506 3.3 0.00059516 0 0.00059508 0 0.00059518 3.3 0.0005951 3.3 0.0005951999999999999 0 0.0005951200000000001 0 0.00059522 3.3 0.0005951400000000001 3.3 0.00059524 0 0.0005951600000000001 0 0.00059526 3.3 0.0005951800000000001 3.3 0.00059528 0 0.0005952 0 0.0005953 3.3 0.00059522 3.3 0.00059532 0 0.00059524 0 0.00059534 3.3 0.00059526 3.3 0.00059536 0 0.00059528 0 0.00059538 3.3 0.0005953 3.3 0.0005953999999999999 0 0.0005953200000000001 0 0.00059542 3.3 0.0005953400000000001 3.3 0.00059544 0 0.0005953600000000001 0 0.00059546 3.3 0.0005953800000000001 3.3 0.00059548 0 0.0005954 0 0.0005955 3.3 0.00059542 3.3 0.00059552 0 0.00059544 0 0.00059554 3.3 0.00059546 3.3 0.00059556 0 0.00059548 0 0.00059558 3.3 0.0005955 3.3 0.0005956 0 0.00059552 0 0.0005956199999999999 3.3 0.0005955400000000001 3.3 0.00059564 0 0.0005955600000000001 0 0.00059566 3.3 0.0005955800000000001 3.3 0.00059568 0 0.0005956000000000001 0 0.0005957 3.3 0.00059562 3.3 0.00059572 0 0.00059564 0 0.00059574 3.3 0.00059566 3.3 0.00059576 0 0.00059568 0 0.00059578 3.3 0.0005957 3.3 0.0005958 0 0.00059572 0 0.0005958199999999999 3.3 0.0005957400000000001 3.3 0.00059584 0 0.0005957600000000001 0 0.00059586 3.3 0.0005957800000000001 3.3 0.00059588 0 0.0005958000000000001 0 0.0005959 3.3 0.00059582 3.3 0.00059592 0 0.00059584 0 0.00059594 3.3 0.00059586 3.3 0.00059596 0 0.00059588 0 0.00059598 3.3 0.0005959 3.3 0.000596 0 0.00059592 0 0.00059602 3.3 0.00059594 3.3 0.0005960399999999999 0 0.0005959600000000001 0 0.00059606 3.3 0.0005959800000000001 3.3 0.00059608 0 0.0005960000000000001 0 0.0005961 3.3 0.0005960200000000001 3.3 0.00059612 0 0.00059604 0 0.00059614 3.3 0.00059606 3.3 0.00059616 0 0.00059608 0 0.00059618 3.3 0.0005961 3.3 0.0005962 0 0.00059612 0 0.00059622 3.3 0.00059614 3.3 0.0005962399999999999 0 0.0005961600000000001 0 0.00059626 3.3 0.0005961800000000001 3.3 0.00059628 0 0.0005962000000000001 0 0.0005963 3.3 0.0005962200000000001 3.3 0.00059632 0 0.00059624 0 0.00059634 3.3 0.00059626 3.3 0.00059636 0 0.00059628 0 0.00059638 3.3 0.0005963 3.3 0.0005964 0 0.00059632 0 0.00059642 3.3 0.00059634 3.3 0.00059644 0 0.00059636 0 0.0005964599999999999 3.3 0.0005963800000000001 3.3 0.00059648 0 0.0005964000000000001 0 0.0005965 3.3 0.0005964200000000001 3.3 0.00059652 0 0.0005964400000000001 0 0.00059654 3.3 0.00059646 3.3 0.00059656 0 0.00059648 0 0.00059658 3.3 0.0005965 3.3 0.0005966 0 0.00059652 0 0.00059662 3.3 0.00059654 3.3 0.00059664 0 0.00059656 0 0.0005966599999999999 3.3 0.0005965800000000001 3.3 0.00059668 0 0.0005966000000000001 0 0.0005967 3.3 0.0005966200000000001 3.3 0.00059672 0 0.0005966400000000001 0 0.00059674 3.3 0.00059666 3.3 0.00059676 0 0.00059668 0 0.00059678 3.3 0.0005967 3.3 0.0005968 0 0.00059672 0 0.00059682 3.3 0.00059674 3.3 0.00059684 0 0.00059676 0 0.00059686 3.3 0.00059678 3.3 0.0005968799999999999 0 0.0005968000000000001 0 0.0005969 3.3 0.0005968200000000001 3.3 0.00059692 0 0.0005968400000000001 0 0.00059694 3.3 0.0005968600000000001 3.3 0.00059696 0 0.00059688 0 0.00059698 3.3 0.0005969 3.3 0.000597 0 0.00059692 0 0.00059702 3.3 0.00059694 3.3 0.00059704 0 0.00059696 0 0.00059706 3.3 0.00059698 3.3 0.0005970799999999999 0 0.0005970000000000001 0 0.0005971 3.3 0.0005970200000000001 3.3 0.00059712 0 0.0005970400000000001 0 0.00059714 3.3 0.0005970600000000001 3.3 0.00059716 0 0.00059708 0 0.00059718 3.3 0.0005971 3.3 0.0005972 0 0.00059712 0 0.00059722 3.3 0.00059714 3.3 0.00059724 0 0.00059716 0 0.00059726 3.3 0.00059718 3.3 0.00059728 0 0.0005972 0 0.0005972999999999999 3.3 0.0005972200000000001 3.3 0.00059732 0 0.0005972400000000001 0 0.00059734 3.3 0.0005972600000000001 3.3 0.00059736 0 0.0005972800000000001 0 0.00059738 3.3 0.0005973 3.3 0.0005974 0 0.00059732 0 0.00059742 3.3 0.00059734 3.3 0.00059744 0 0.00059736 0 0.00059746 3.3 0.00059738 3.3 0.00059748 0 0.0005974 0 0.0005974999999999999 3.3 0.0005974200000000001 3.3 0.00059752 0 0.0005974400000000001 0 0.00059754 3.3 0.0005974600000000001 3.3 0.00059756 0 0.0005974800000000001 0 0.00059758 3.3 0.0005975 3.3 0.0005976 0 0.00059752 0 0.00059762 3.3 0.00059754 3.3 0.00059764 0 0.00059756 0 0.00059766 3.3 0.00059758 3.3 0.00059768 0 0.0005976 0 0.0005976999999999999 3.3 0.00059762 3.3 0.0005977199999999999 0 0.0005976400000000001 0 0.00059774 3.3 0.0005976600000000001 3.3 0.00059776 0 0.0005976800000000001 0 0.00059778 3.3 0.0005977 3.3 0.0005978 0 0.00059772 0 0.00059782 3.3 0.00059774 3.3 0.00059784 0 0.00059776 0 0.00059786 3.3 0.00059778 3.3 0.00059788 0 0.0005978 0 0.0005979 3.3 0.00059782 3.3 0.0005979199999999999 0 0.0005978400000000001 0 0.00059794 3.3 0.0005978600000000001 3.3 0.00059796 0 0.0005978800000000001 0 0.00059798 3.3 0.0005979000000000001 3.3 0.000598 0 0.00059792 0 0.00059802 3.3 0.00059794 3.3 0.00059804 0 0.00059796 0 0.00059806 3.3 0.00059798 3.3 0.00059808 0 0.000598 0 0.0005981 3.3 0.00059802 3.3 0.0005981199999999999 0 0.00059804 0 0.0005981399999999999 3.3 0.0005980600000000001 3.3 0.00059816 0 0.0005980800000000001 0 0.00059818 3.3 0.0005981000000000001 3.3 0.0005982 0 0.00059812 0 0.00059822 3.3 0.00059814 3.3 0.00059824 0 0.00059816 0 0.00059826 3.3 0.00059818 3.3 0.00059828 0 0.0005982 0 0.0005983 3.3 0.00059822 3.3 0.00059832 0 0.00059824 0 0.0005983399999999999 3.3 0.0005982600000000001 3.3 0.00059836 0 0.0005982800000000001 0 0.00059838 3.3 0.0005983000000000001 3.3 0.0005984 0 0.0005983200000000001 0 0.00059842 3.3 0.00059834 3.3 0.00059844 0 0.00059836 0 0.00059846 3.3 0.00059838 3.3 0.00059848 0 0.0005984 0 0.0005985 3.3 0.00059842 3.3 0.00059852 0 0.00059844 0 0.0005985399999999999 3.3 0.00059846 3.3 0.0005985599999999999 0 0.0005984800000000001 0 0.00059858 3.3 0.0005985000000000001 3.3 0.0005986 0 0.0005985200000000001 0 0.00059862 3.3 0.00059854 3.3 0.00059864 0 0.00059856 0 0.00059866 3.3 0.00059858 3.3 0.00059868 0 0.0005986 0 0.0005987 3.3 0.00059862 3.3 0.00059872 0 0.00059864 0 0.00059874 3.3 0.00059866 3.3 0.0005987599999999999 0 0.0005986800000000001 0 0.00059878 3.3 0.0005987000000000001 3.3 0.0005988 0 0.0005987200000000001 0 0.00059882 3.3 0.0005987400000000001 3.3 0.00059884 0 0.00059876 0 0.00059886 3.3 0.00059878 3.3 0.00059888 0 0.0005988 0 0.0005989 3.3 0.00059882 3.3 0.00059892 0 0.00059884 0 0.00059894 3.3 0.00059886 3.3 0.0005989599999999999 0 0.0005988800000000001 0 0.00059898 3.3 0.0005989000000000001 3.3 0.000599 0 0.0005989200000000001 0 0.00059902 3.3 0.0005989400000000001 3.3 0.00059904 0 0.00059896 0 0.00059906 3.3 0.00059898 3.3 0.00059908 0 0.000599 0 0.0005991 3.3 0.00059902 3.3 0.00059912 0 0.00059904 0 0.00059914 3.3 0.00059906 3.3 0.00059916 0 0.00059908 0 0.0005991799999999999 3.3 0.0005991000000000001 3.3 0.0005992 0 0.0005991200000000001 0 0.00059922 3.3 0.0005991400000000001 3.3 0.00059924 0 0.0005991600000000001 0 0.00059926 3.3 0.00059918 3.3 0.00059928 0 0.0005992 0 0.0005993 3.3 0.00059922 3.3 0.00059932 0 0.00059924 0 0.00059934 3.3 0.00059926 3.3 0.00059936 0 0.00059928 0 0.0005993799999999999 3.3 0.0005993000000000001 3.3 0.0005994 0 0.0005993200000000001 0 0.00059942 3.3 0.0005993400000000001 3.3 0.00059944 0 0.0005993600000000001 0 0.00059946 3.3 0.00059938 3.3 0.00059948 0 0.0005994 0 0.0005995 3.3 0.00059942 3.3 0.00059952 0 0.00059944 0 0.00059954 3.3 0.00059946 3.3 0.00059956 0 0.00059948 0 0.00059958 3.3 0.0005995 3.3 0.0005995999999999999 0 0.0005995200000000001 0 0.00059962 3.3 0.0005995400000000001 3.3 0.00059964 0 0.0005995600000000001 0 0.00059966 3.3 0.0005995800000000001 3.3 0.00059968 0 0.0005996 0 0.0005997 3.3 0.00059962 3.3 0.00059972 0 0.00059964 0 0.00059974 3.3 0.00059966 3.3 0.00059976 0 0.00059968 0 0.00059978 3.3 0.0005997 3.3 0.0005997999999999999 0 0.0005997200000000001 0 0.00059982 3.3 0.0005997400000000001 3.3 0.00059984 0 0.0005997600000000001 0 0.00059986 3.3 0.0005997800000000001 3.3 0.00059988 0 0.0005998 0 0.0005999 3.3 0.00059982 3.3 0.00059992 0 0.00059984 0 0.00059994 3.3 0.00059986 3.3 0.00059996 0 0.00059988 0 0.00059998 3.3 0.0005999 3.3 0.0006 0 0.00059992 0 0.0006000199999999999 3.3 0.0005999400000000001 3.3 0.00060004 0 0.0005999600000000001 0 0.00060006 3.3 0.0005999800000000001 3.3 0.00060008 0 0.0006000000000000001 0 0.0006001 3.3 0.00060002 3.3 0.00060012 0 0.00060004 0 0.00060014 3.3 0.00060006 3.3 0.00060016 0 0.00060008 0 0.00060018 3.3 0.0006001 3.3 0.0006002 0 0.00060012 0 0.0006002199999999999 3.3 0.0006001400000000001 3.3 0.00060024 0 0.0006001600000000001 0 0.00060026 3.3 0.0006001800000000001 3.3 0.00060028 0 0.0006002000000000001 0 0.0006003 3.3 0.00060022 3.3 0.00060032 0 0.00060024 0 0.00060034 3.3 0.00060026 3.3 0.00060036 0 0.00060028 0 0.00060038 3.3 0.0006003 3.3 0.0006004 0 0.00060032 0 0.00060042 3.3 0.00060034 3.3 0.0006004399999999999 0 0.0006003600000000001 0 0.00060046 3.3 0.0006003800000000001 3.3 0.00060048 0 0.0006004000000000001 0 0.0006005 3.3 0.0006004200000000001 3.3 0.00060052 0 0.00060044 0 0.00060054 3.3 0.00060046 3.3 0.00060056 0 0.00060048 0 0.00060058 3.3 0.0006005 3.3 0.0006006 0 0.00060052 0 0.00060062 3.3 0.00060054 3.3 0.0006006399999999999 0 0.0006005600000000001 0 0.00060066 3.3 0.0006005800000000001 3.3 0.00060068 0 0.0006006000000000001 0 0.0006007 3.3 0.0006006200000000001 3.3 0.00060072 0 0.00060064 0 0.00060074 3.3 0.00060066 3.3 0.00060076 0 0.00060068 0 0.00060078 3.3 0.0006007 3.3 0.0006008 0 0.00060072 0 0.00060082 3.3 0.00060074 3.3 0.00060084 0 0.00060076 0 0.0006008599999999999 3.3 0.0006007800000000001 3.3 0.00060088 0 0.0006008000000000001 0 0.0006009 3.3 0.0006008200000000001 3.3 0.00060092 0 0.0006008400000000001 0 0.00060094 3.3 0.00060086 3.3 0.00060096 0 0.00060088 0 0.00060098 3.3 0.0006009 3.3 0.000601 0 0.00060092 0 0.00060102 3.3 0.00060094 3.3 0.00060104 0 0.00060096 0 0.0006010599999999999 3.3 0.0006009800000000001 3.3 0.00060108 0 0.0006010000000000001 0 0.0006011 3.3 0.0006010200000000001 3.3 0.00060112 0 0.0006010400000000001 0 0.00060114 3.3 0.00060106 3.3 0.00060116 0 0.00060108 0 0.00060118 3.3 0.0006011 3.3 0.0006012 0 0.00060112 0 0.00060122 3.3 0.00060114 3.3 0.00060124 0 0.00060116 0 0.0006012599999999999 3.3 0.00060118 3.3 0.0006012799999999999 0 0.0006012000000000001 0 0.0006013 3.3 0.0006012200000000001 3.3 0.00060132 0 0.0006012400000000001 0 0.00060134 3.3 0.00060126 3.3 0.00060136 0 0.00060128 0 0.00060138 3.3 0.0006013 3.3 0.0006014 0 0.00060132 0 0.00060142 3.3 0.00060134 3.3 0.00060144 0 0.00060136 0 0.00060146 3.3 0.00060138 3.3 0.0006014799999999999 0 0.0006014000000000001 0 0.0006015 3.3 0.0006014200000000001 3.3 0.00060152 0 0.0006014400000000001 0 0.00060154 3.3 0.0006014600000000001 3.3 0.00060156 0 0.00060148 0 0.00060158 3.3 0.0006015 3.3 0.0006016 0 0.00060152 0 0.00060162 3.3 0.00060154 3.3 0.00060164 0 0.00060156 0 0.00060166 3.3 0.00060158 3.3 0.0006016799999999999 0 0.0006016 0 0.0006016999999999999 3.3 0.0006016200000000001 3.3 0.00060172 0 0.0006016400000000001 0 0.00060174 3.3 0.0006016600000000001 3.3 0.00060176 0 0.00060168 0 0.00060178 3.3 0.0006017 3.3 0.0006018 0 0.00060172 0 0.00060182 3.3 0.00060174 3.3 0.00060184 0 0.00060176 0 0.00060186 3.3 0.00060178 3.3 0.00060188 0 0.0006018 0 0.0006018999999999999 3.3 0.0006018200000000001 3.3 0.00060192 0 0.0006018400000000001 0 0.00060194 3.3 0.0006018600000000001 3.3 0.00060196 0 0.0006018800000000001 0 0.00060198 3.3 0.0006019 3.3 0.000602 0 0.00060192 0 0.00060202 3.3 0.00060194 3.3 0.00060204 0 0.00060196 0 0.00060206 3.3 0.00060198 3.3 0.00060208 0 0.000602 0 0.0006020999999999999 3.3 0.00060202 3.3 0.0006021199999999999 0 0.0006020400000000001 0 0.00060214 3.3 0.0006020600000000001 3.3 0.00060216 0 0.0006020800000000001 0 0.00060218 3.3 0.0006021 3.3 0.0006022 0 0.00060212 0 0.00060222 3.3 0.00060214 3.3 0.00060224 0 0.00060216 0 0.00060226 3.3 0.00060218 3.3 0.00060228 0 0.0006022 0 0.0006023 3.3 0.00060222 3.3 0.0006023199999999999 0 0.0006022400000000001 0 0.00060234 3.3 0.0006022600000000001 3.3 0.00060236 0 0.0006022800000000001 0 0.00060238 3.3 0.0006023000000000001 3.3 0.0006024 0 0.00060232 0 0.00060242 3.3 0.00060234 3.3 0.00060244 0 0.00060236 0 0.00060246 3.3 0.00060238 3.3 0.00060248 0 0.0006024 0 0.0006025 3.3 0.00060242 3.3 0.0006025199999999999 0 0.0006024400000000001 0 0.00060254 3.3 0.0006024600000000001 3.3 0.00060256 0 0.0006024800000000001 0 0.00060258 3.3 0.0006025000000000001 3.3 0.0006026 0 0.00060252 0 0.00060262 3.3 0.00060254 3.3 0.00060264 0 0.00060256 0 0.00060266 3.3 0.00060258 3.3 0.00060268 0 0.0006026 0 0.0006027 3.3 0.00060262 3.3 0.00060272 0 0.00060264 0 0.0006027399999999999 3.3 0.0006026600000000001 3.3 0.00060276 0 0.0006026800000000001 0 0.00060278 3.3 0.0006027000000000001 3.3 0.0006028 0 0.0006027200000000001 0 0.00060282 3.3 0.00060274 3.3 0.00060284 0 0.00060276 0 0.00060286 3.3 0.00060278 3.3 0.00060288 0 0.0006028 0 0.0006029 3.3 0.00060282 3.3 0.00060292 0 0.00060284 0 0.0006029399999999999 3.3 0.0006028600000000001 3.3 0.00060296 0 0.0006028800000000001 0 0.00060298 3.3 0.0006029000000000001 3.3 0.000603 0 0.0006029200000000001 0 0.00060302 3.3 0.00060294 3.3 0.00060304 0 0.00060296 0 0.00060306 3.3 0.00060298 3.3 0.00060308 0 0.000603 0 0.0006031 3.3 0.00060302 3.3 0.00060312 0 0.00060304 0 0.00060314 3.3 0.00060306 3.3 0.0006031599999999999 0 0.0006030800000000001 0 0.00060318 3.3 0.0006031000000000001 3.3 0.0006032 0 0.0006031200000000001 0 0.00060322 3.3 0.0006031400000000001 3.3 0.00060324 0 0.00060316 0 0.00060326 3.3 0.00060318 3.3 0.00060328 0 0.0006032 0 0.0006033 3.3 0.00060322 3.3 0.00060332 0 0.00060324 0 0.00060334 3.3 0.00060326 3.3 0.0006033599999999999 0 0.0006032800000000001 0 0.00060338 3.3 0.0006033000000000001 3.3 0.0006034 0 0.0006033200000000001 0 0.00060342 3.3 0.0006033400000000001 3.3 0.00060344 0 0.00060336 0 0.00060346 3.3 0.00060338 3.3 0.00060348 0 0.0006034 0 0.0006035 3.3 0.00060342 3.3 0.00060352 0 0.00060344 0 0.00060354 3.3 0.00060346 3.3 0.00060356 0 0.00060348 0 0.0006035799999999999 3.3 0.0006035000000000001 3.3 0.0006036 0 0.0006035200000000001 0 0.00060362 3.3 0.0006035400000000001 3.3 0.00060364 0 0.0006035600000000001 0 0.00060366 3.3 0.00060358 3.3 0.00060368 0 0.0006036 0 0.0006037 3.3 0.00060362 3.3 0.00060372 0 0.00060364 0 0.00060374 3.3 0.00060366 3.3 0.00060376 0 0.00060368 0 0.0006037799999999999 3.3 0.0006037000000000001 3.3 0.0006038 0 0.0006037200000000001 0 0.00060382 3.3 0.0006037400000000001 3.3 0.00060384 0 0.0006037600000000001 0 0.00060386 3.3 0.00060378 3.3 0.00060388 0 0.0006038 0 0.0006039 3.3 0.00060382 3.3 0.00060392 0 0.00060384 0 0.00060394 3.3 0.00060386 3.3 0.00060396 0 0.00060388 0 0.00060398 3.3 0.0006039 3.3 0.0006039999999999999 0 0.0006039200000000001 0 0.00060402 3.3 0.0006039400000000001 3.3 0.00060404 0 0.0006039600000000001 0 0.00060406 3.3 0.0006039800000000001 3.3 0.00060408 0 0.000604 0 0.0006041 3.3 0.00060402 3.3 0.00060412 0 0.00060404 0 0.00060414 3.3 0.00060406 3.3 0.00060416 0 0.00060408 0 0.00060418 3.3 0.0006041 3.3 0.0006041999999999999 0 0.0006041200000000001 0 0.00060422 3.3 0.0006041400000000001 3.3 0.00060424 0 0.0006041600000000001 0 0.00060426 3.3 0.0006041800000000001 3.3 0.00060428 0 0.0006042 0 0.0006043 3.3 0.00060422 3.3 0.00060432 0 0.00060424 0 0.00060434 3.3 0.00060426 3.3 0.00060436 0 0.00060428 0 0.00060438 3.3 0.0006043 3.3 0.0006044 0 0.00060432 0 0.0006044199999999999 3.3 0.0006043400000000001 3.3 0.00060444 0 0.0006043600000000001 0 0.00060446 3.3 0.0006043800000000001 3.3 0.00060448 0 0.0006044000000000001 0 0.0006045 3.3 0.00060442 3.3 0.00060452 0 0.00060444 0 0.00060454 3.3 0.00060446 3.3 0.00060456 0 0.00060448 0 0.00060458 3.3 0.0006045 3.3 0.0006046 0 0.00060452 0 0.0006046199999999999 3.3 0.0006045400000000001 3.3 0.00060464 0 0.0006045600000000001 0 0.00060466 3.3 0.0006045800000000001 3.3 0.00060468 0 0.0006046000000000001 0 0.0006047 3.3 0.00060462 3.3 0.00060472 0 0.00060464 0 0.00060474 3.3 0.00060466 3.3 0.00060476 0 0.00060468 0 0.00060478 3.3 0.0006047 3.3 0.0006048 0 0.00060472 0 0.0006048199999999999 3.3 0.00060474 3.3 0.0006048399999999999 0 0.0006047600000000001 0 0.00060486 3.3 0.0006047800000000001 3.3 0.00060488 0 0.0006048000000000001 0 0.0006049 3.3 0.00060482 3.3 0.00060492 0 0.00060484 0 0.00060494 3.3 0.00060486 3.3 0.00060496 0 0.00060488 0 0.00060498 3.3 0.0006049 3.3 0.000605 0 0.00060492 0 0.00060502 3.3 0.00060494 3.3 0.0006050399999999999 0 0.0006049600000000001 0 0.00060506 3.3 0.0006049800000000001 3.3 0.00060508 0 0.0006050000000000001 0 0.0006051 3.3 0.0006050200000000001 3.3 0.00060512 0 0.00060504 0 0.00060514 3.3 0.00060506 3.3 0.00060516 0 0.00060508 0 0.00060518 3.3 0.0006051 3.3 0.0006052 0 0.00060512 0 0.00060522 3.3 0.00060514 3.3 0.0006052399999999999 0 0.00060516 0 0.0006052599999999999 3.3 0.0006051800000000001 3.3 0.00060528 0 0.0006052000000000001 0 0.0006053 3.3 0.0006052200000000001 3.3 0.00060532 0 0.00060524 0 0.00060534 3.3 0.00060526 3.3 0.00060536 0 0.00060528 0 0.00060538 3.3 0.0006053 3.3 0.0006054 0 0.00060532 0 0.00060542 3.3 0.00060534 3.3 0.00060544 0 0.00060536 0 0.0006054599999999999 3.3 0.0006053800000000001 3.3 0.00060548 0 0.0006054000000000001 0 0.0006055 3.3 0.0006054200000000001 3.3 0.00060552 0 0.0006054400000000001 0 0.00060554 3.3 0.00060546 3.3 0.00060556 0 0.00060548 0 0.00060558 3.3 0.0006055 3.3 0.0006056 0 0.00060552 0 0.00060562 3.3 0.00060554 3.3 0.00060564 0 0.00060556 0 0.0006056599999999999 3.3 0.00060558 3.3 0.0006056799999999999 0 0.0006056000000000001 0 0.0006057 3.3 0.0006056200000000001 3.3 0.00060572 0 0.0006056400000000001 0 0.00060574 3.3 0.00060566 3.3 0.00060576 0 0.00060568 0 0.00060578 3.3 0.0006057 3.3 0.0006058 0 0.00060572 0 0.00060582 3.3 0.00060574 3.3 0.00060584 0 0.00060576 0 0.00060586 3.3 0.00060578 3.3 0.0006058799999999999 0 0.0006058000000000001 0 0.0006059 3.3 0.0006058200000000001 3.3 0.00060592 0 0.0006058400000000001 0 0.00060594 3.3 0.0006058600000000001 3.3 0.00060596 0 0.00060588 0 0.00060598 3.3 0.0006059 3.3 0.000606 0 0.00060592 0 0.00060602 3.3 0.00060594 3.3 0.00060604 0 0.00060596 0 0.00060606 3.3 0.00060598 3.3 0.0006060799999999999 0 0.0006060000000000001 0 0.0006061 3.3 0.0006060200000000001 3.3 0.00060612 0 0.0006060400000000001 0 0.00060614 3.3 0.0006060600000000001 3.3 0.00060616 0 0.00060608 0 0.00060618 3.3 0.0006061 3.3 0.0006062 0 0.00060612 0 0.00060622 3.3 0.00060614 3.3 0.00060624 0 0.00060616 0 0.00060626 3.3 0.00060618 3.3 0.00060628 0 0.0006062 0 0.0006062999999999999 3.3 0.0006062200000000001 3.3 0.00060632 0 0.0006062400000000001 0 0.00060634 3.3 0.0006062600000000001 3.3 0.00060636 0 0.0006062800000000001 0 0.00060638 3.3 0.0006063 3.3 0.0006064 0 0.00060632 0 0.00060642 3.3 0.00060634 3.3 0.00060644 0 0.00060636 0 0.00060646 3.3 0.00060638 3.3 0.00060648 0 0.0006064 0 0.0006064999999999999 3.3 0.0006064200000000001 3.3 0.00060652 0 0.0006064400000000001 0 0.00060654 3.3 0.0006064600000000001 3.3 0.00060656 0 0.0006064800000000001 0 0.00060658 3.3 0.0006065 3.3 0.0006066 0 0.00060652 0 0.00060662 3.3 0.00060654 3.3 0.00060664 0 0.00060656 0 0.00060666 3.3 0.00060658 3.3 0.00060668 0 0.0006066 0 0.0006067 3.3 0.00060662 3.3 0.0006067199999999999 0 0.0006066400000000001 0 0.00060674 3.3 0.0006066600000000001 3.3 0.00060676 0 0.0006066800000000001 0 0.00060678 3.3 0.0006067000000000001 3.3 0.0006068 0 0.00060672 0 0.00060682 3.3 0.00060674 3.3 0.00060684 0 0.00060676 0 0.00060686 3.3 0.00060678 3.3 0.00060688 0 0.0006068 0 0.0006069 3.3 0.00060682 3.3 0.0006069199999999999 0 0.0006068400000000001 0 0.00060694 3.3 0.0006068600000000001 3.3 0.00060696 0 0.0006068800000000001 0 0.00060698 3.3 0.0006069000000000001 3.3 0.000607 0 0.00060692 0 0.00060702 3.3 0.00060694 3.3 0.00060704 0 0.00060696 0 0.00060706 3.3 0.00060698 3.3 0.00060708 0 0.000607 0 0.0006071 3.3 0.00060702 3.3 0.00060712 0 0.00060704 0 0.0006071399999999999 3.3 0.0006070600000000001 3.3 0.00060716 0 0.0006070800000000001 0 0.00060718 3.3 0.0006071000000000001 3.3 0.0006072 0 0.0006071200000000001 0 0.00060722 3.3 0.00060714 3.3 0.00060724 0 0.00060716 0 0.00060726 3.3 0.00060718 3.3 0.00060728 0 0.0006072 0 0.0006073 3.3 0.00060722 3.3 0.00060732 0 0.00060724 0 0.0006073399999999999 3.3 0.0006072600000000001 3.3 0.00060736 0 0.0006072800000000001 0 0.00060738 3.3 0.0006073000000000001 3.3 0.0006074 0 0.0006073200000000001 0 0.00060742 3.3 0.00060734 3.3 0.00060744 0 0.00060736 0 0.00060746 3.3 0.00060738 3.3 0.00060748 0 0.0006074 0 0.0006075 3.3 0.00060742 3.3 0.00060752 0 0.00060744 0 0.00060754 3.3 0.00060746 3.3 0.0006075599999999999 0 0.0006074800000000001 0 0.00060758 3.3 0.0006075000000000001 3.3 0.0006076 0 0.0006075200000000001 0 0.00060762 3.3 0.0006075400000000001 3.3 0.00060764 0 0.00060756 0 0.00060766 3.3 0.00060758 3.3 0.00060768 0 0.0006076 0 0.0006077 3.3 0.00060762 3.3 0.00060772 0 0.00060764 0 0.00060774 3.3 0.00060766 3.3 0.0006077599999999999 0 0.0006076800000000001 0 0.00060778 3.3 0.0006077000000000001 3.3 0.0006078 0 0.0006077200000000001 0 0.00060782 3.3 0.0006077400000000001 3.3 0.00060784 0 0.00060776 0 0.00060786 3.3 0.00060778 3.3 0.00060788 0 0.0006078 0 0.0006079 3.3 0.00060782 3.3 0.00060792 0 0.00060784 0 0.00060794 3.3 0.00060786 3.3 0.0006079599999999999 0 0.00060788 0 0.0006079799999999999 3.3 0.0006079000000000001 3.3 0.000608 0 0.0006079200000000001 0 0.00060802 3.3 0.0006079400000000001 3.3 0.00060804 0 0.00060796 0 0.00060806 3.3 0.00060798 3.3 0.00060808 0 0.000608 0 0.0006081 3.3 0.00060802 3.3 0.00060812 0 0.00060804 0 0.00060814 3.3 0.00060806 3.3 0.00060816 0 0.00060808 0 0.0006081799999999999 3.3 0.0006081000000000001 3.3 0.0006082 0 0.0006081200000000001 0 0.00060822 3.3 0.0006081400000000001 3.3 0.00060824 0 0.0006081600000000001 0 0.00060826 3.3 0.00060818 3.3 0.00060828 0 0.0006082 0 0.0006083 3.3 0.00060822 3.3 0.00060832 0 0.00060824 0 0.00060834 3.3 0.00060826 3.3 0.00060836 0 0.00060828 0 0.0006083799999999999 3.3 0.0006083 3.3 0.0006083999999999999 0 0.0006083200000000001 0 0.00060842 3.3 0.0006083400000000001 3.3 0.00060844 0 0.0006083600000000001 0 0.00060846 3.3 0.00060838 3.3 0.00060848 0 0.0006084 0 0.0006085 3.3 0.00060842 3.3 0.00060852 0 0.00060844 0 0.00060854 3.3 0.00060846 3.3 0.00060856 0 0.00060848 0 0.00060858 3.3 0.0006085 3.3 0.0006085999999999999 0 0.0006085200000000001 0 0.00060862 3.3 0.0006085400000000001 3.3 0.00060864 0 0.0006085600000000001 0 0.00060866 3.3 0.0006085800000000001 3.3 0.00060868 0 0.0006086 0 0.0006087 3.3 0.00060862 3.3 0.00060872 0 0.00060864 0 0.00060874 3.3 0.00060866 3.3 0.00060876 0 0.00060868 0 0.00060878 3.3 0.0006087 3.3 0.0006087999999999999 0 0.00060872 0 0.0006088199999999999 3.3 0.0006087400000000001 3.3 0.00060884 0 0.0006087600000000001 0 0.00060886 3.3 0.0006087800000000001 3.3 0.00060888 0 0.0006088 0 0.0006089 3.3 0.00060882 3.3 0.00060892 0 0.00060884 0 0.00060894 3.3 0.00060886 3.3 0.00060896 0 0.00060888 0 0.00060898 3.3 0.0006089 3.3 0.000609 0 0.00060892 0 0.0006090199999999999 3.3 0.0006089400000000001 3.3 0.00060904 0 0.0006089600000000001 0 0.00060906 3.3 0.0006089800000000001 3.3 0.00060908 0 0.0006090000000000001 0 0.0006091 3.3 0.00060902 3.3 0.00060912 0 0.00060904 0 0.00060914 3.3 0.00060906 3.3 0.00060916 0 0.00060908 0 0.00060918 3.3 0.0006091 3.3 0.0006092 0 0.00060912 0 0.0006092199999999999 3.3 0.0006091400000000001 3.3 0.00060924 0 0.0006091600000000001 0 0.00060926 3.3 0.0006091800000000001 3.3 0.00060928 0 0.0006092000000000001 0 0.0006093 3.3 0.00060922 3.3 0.00060932 0 0.00060924 0 0.00060934 3.3 0.00060926 3.3 0.00060936 0 0.00060928 0 0.00060938 3.3 0.0006093 3.3 0.0006094 0 0.00060932 0 0.00060942 3.3 0.00060934 3.3 0.0006094399999999999 0 0.0006093600000000001 0 0.00060946 3.3 0.0006093800000000001 3.3 0.00060948 0 0.0006094000000000001 0 0.0006095 3.3 0.0006094200000000001 3.3 0.00060952 0 0.00060944 0 0.00060954 3.3 0.00060946 3.3 0.00060956 0 0.00060948 0 0.00060958 3.3 0.0006095 3.3 0.0006096 0 0.00060952 0 0.00060962 3.3 0.00060954 3.3 0.0006096399999999999 0 0.0006095600000000001 0 0.00060966 3.3 0.0006095800000000001 3.3 0.00060968 0 0.0006096000000000001 0 0.0006097 3.3 0.0006096200000000001 3.3 0.00060972 0 0.00060964 0 0.00060974 3.3 0.00060966 3.3 0.00060976 0 0.00060968 0 0.00060978 3.3 0.0006097 3.3 0.0006098 0 0.00060972 0 0.00060982 3.3 0.00060974 3.3 0.00060984 0 0.00060976 0 0.0006098599999999999 3.3 0.0006097800000000001 3.3 0.00060988 0 0.0006098000000000001 0 0.0006099 3.3 0.0006098200000000001 3.3 0.00060992 0 0.0006098400000000001 0 0.00060994 3.3 0.00060986 3.3 0.00060996 0 0.00060988 0 0.00060998 3.3 0.0006099 3.3 0.00061 0 0.00060992 0 0.00061002 3.3 0.00060994 3.3 0.00061004 0 0.00060996 0 0.0006100599999999999 3.3 0.0006099800000000001 3.3 0.00061008 0 0.0006100000000000001 0 0.0006101 3.3 0.0006100200000000001 3.3 0.00061012 0 0.0006100400000000001 0 0.00061014 3.3 0.00061006 3.3 0.00061016 0 0.00061008 0 0.00061018 3.3 0.0006101 3.3 0.0006102 0 0.00061012 0 0.00061022 3.3 0.00061014 3.3 0.00061024 0 0.00061016 0 0.00061026 3.3 0.00061018 3.3 0.0006102799999999999 0 0.0006102000000000001 0 0.0006103 3.3 0.0006102200000000001 3.3 0.00061032 0 0.0006102400000000001 0 0.00061034 3.3 0.0006102600000000001 3.3 0.00061036 0 0.00061028 0 0.00061038 3.3 0.0006103 3.3 0.0006104 0 0.00061032 0 0.00061042 3.3 0.00061034 3.3 0.00061044 0 0.00061036 0 0.00061046 3.3 0.00061038 3.3 0.0006104799999999999 0 0.0006104000000000001 0 0.0006105 3.3 0.0006104200000000001 3.3 0.00061052 0 0.0006104400000000001 0 0.00061054 3.3 0.0006104600000000001 3.3 0.00061056 0 0.00061048 0 0.00061058 3.3 0.0006105 3.3 0.0006106 0 0.00061052 0 0.00061062 3.3 0.00061054 3.3 0.00061064 0 0.00061056 0 0.00061066 3.3 0.00061058 3.3 0.00061068 0 0.0006106 0 0.0006106999999999999 3.3 0.0006106200000000001 3.3 0.00061072 0 0.0006106400000000001 0 0.00061074 3.3 0.0006106600000000001 3.3 0.00061076 0 0.0006106800000000001 0 0.00061078 3.3 0.0006107 3.3 0.0006108 0 0.00061072 0 0.00061082 3.3 0.00061074 3.3 0.00061084 0 0.00061076 0 0.00061086 3.3 0.00061078 3.3 0.00061088 0 0.0006108 0 0.0006108999999999999 3.3 0.0006108200000000001 3.3 0.00061092 0 0.0006108400000000001 0 0.00061094 3.3 0.0006108600000000001 3.3 0.00061096 0 0.0006108800000000001 0 0.00061098 3.3 0.0006109 3.3 0.000611 0 0.00061092 0 0.00061102 3.3 0.00061094 3.3 0.00061104 0 0.00061096 0 0.00061106 3.3 0.00061098 3.3 0.00061108 0 0.000611 0 0.0006111 3.3 0.00061102 3.3 0.0006111199999999999 0 0.0006110400000000001 0 0.00061114 3.3 0.0006110600000000001 3.3 0.00061116 0 0.0006110800000000001 0 0.00061118 3.3 0.0006111000000000001 3.3 0.0006112 0 0.00061112 0 0.00061122 3.3 0.00061114 3.3 0.00061124 0 0.00061116 0 0.00061126 3.3 0.00061118 3.3 0.00061128 0 0.0006112 0 0.0006113 3.3 0.00061122 3.3 0.0006113199999999999 0 0.0006112400000000001 0 0.00061134 3.3 0.0006112600000000001 3.3 0.00061136 0 0.0006112800000000001 0 0.00061138 3.3 0.0006113000000000001 3.3 0.0006114 0 0.00061132 0 0.00061142 3.3 0.00061134 3.3 0.00061144 0 0.00061136 0 0.00061146 3.3 0.00061138 3.3 0.00061148 0 0.0006114 0 0.0006115 3.3 0.00061142 3.3 0.0006115199999999999 0 0.00061144 0 0.0006115399999999999 3.3 0.0006114600000000001 3.3 0.00061156 0 0.0006114800000000001 0 0.00061158 3.3 0.0006115000000000001 3.3 0.0006116 0 0.00061152 0 0.00061162 3.3 0.00061154 3.3 0.00061164 0 0.00061156 0 0.00061166 3.3 0.00061158 3.3 0.00061168 0 0.0006116 0 0.0006117 3.3 0.00061162 3.3 0.00061172 0 0.00061164 0 0.0006117399999999999 3.3 0.0006116600000000001 3.3 0.00061176 0 0.0006116800000000001 0 0.00061178 3.3 0.0006117000000000001 3.3 0.0006118 0 0.0006117200000000001 0 0.00061182 3.3 0.00061174 3.3 0.00061184 0 0.00061176 0 0.00061186 3.3 0.00061178 3.3 0.00061188 0 0.0006118 0 0.0006119 3.3 0.00061182 3.3 0.00061192 0 0.00061184 0 0.0006119399999999999 3.3 0.00061186 3.3 0.0006119599999999999 0 0.0006118800000000001 0 0.00061198 3.3 0.0006119000000000001 3.3 0.000612 0 0.0006119200000000001 0 0.00061202 3.3 0.00061194 3.3 0.00061204 0 0.00061196 0 0.00061206 3.3 0.00061198 3.3 0.00061208 0 0.000612 0 0.0006121 3.3 0.00061202 3.3 0.00061212 0 0.00061204 0 0.00061214 3.3 0.00061206 3.3 0.0006121599999999999 0 0.0006120800000000001 0 0.00061218 3.3 0.0006121000000000001 3.3 0.0006122 0 0.0006121200000000001 0 0.00061222 3.3 0.0006121400000000001 3.3 0.00061224 0 0.00061216 0 0.00061226 3.3 0.00061218 3.3 0.00061228 0 0.0006122 0 0.0006123 3.3 0.00061222 3.3 0.00061232 0 0.00061224 0 0.00061234 3.3 0.00061226 3.3 0.0006123599999999999 0 0.00061228 0 0.0006123799999999999 3.3 0.0006123000000000001 3.3 0.0006124 0 0.0006123200000000001 0 0.00061242 3.3 0.0006123400000000001 3.3 0.00061244 0 0.00061236 0 0.00061246 3.3 0.00061238 3.3 0.00061248 0 0.0006124 0 0.0006125 3.3 0.00061242 3.3 0.00061252 0 0.00061244 0 0.00061254 3.3 0.00061246 3.3 0.00061256 0 0.00061248 0 0.0006125799999999999 3.3 0.0006125000000000001 3.3 0.0006126 0 0.0006125200000000001 0 0.00061262 3.3 0.0006125400000000001 3.3 0.00061264 0 0.0006125600000000001 0 0.00061266 3.3 0.00061258 3.3 0.00061268 0 0.0006126 0 0.0006127 3.3 0.00061262 3.3 0.00061272 0 0.00061264 0 0.00061274 3.3 0.00061266 3.3 0.00061276 0 0.00061268 0 0.0006127799999999999 3.3 0.0006127000000000001 3.3 0.0006128 0 0.0006127200000000001 0 0.00061282 3.3 0.0006127400000000001 3.3 0.00061284 0 0.0006127600000000001 0 0.00061286 3.3 0.00061278 3.3 0.00061288 0 0.0006128 0 0.0006129 3.3 0.00061282 3.3 0.00061292 0 0.00061284 0 0.00061294 3.3 0.00061286 3.3 0.00061296 0 0.00061288 0 0.00061298 3.3 0.0006129 3.3 0.0006129999999999999 0 0.0006129200000000001 0 0.00061302 3.3 0.0006129400000000001 3.3 0.00061304 0 0.0006129600000000001 0 0.00061306 3.3 0.0006129800000000001 3.3 0.00061308 0 0.000613 0 0.0006131 3.3 0.00061302 3.3 0.00061312 0 0.00061304 0 0.00061314 3.3 0.00061306 3.3 0.00061316 0 0.00061308 0 0.00061318 3.3 0.0006131 3.3 0.0006131999999999999 0 0.0006131200000000001 0 0.00061322 3.3 0.0006131400000000001 3.3 0.00061324 0 0.0006131600000000001 0 0.00061326 3.3 0.0006131800000000001 3.3 0.00061328 0 0.0006132 0 0.0006133 3.3 0.00061322 3.3 0.00061332 0 0.00061324 0 0.00061334 3.3 0.00061326 3.3 0.00061336 0 0.00061328 0 0.00061338 3.3 0.0006133 3.3 0.0006134 0 0.00061332 0 0.0006134199999999999 3.3 0.0006133400000000001 3.3 0.00061344 0 0.0006133600000000001 0 0.00061346 3.3 0.0006133800000000001 3.3 0.00061348 0 0.0006134000000000001 0 0.0006135 3.3 0.00061342 3.3 0.00061352 0 0.00061344 0 0.00061354 3.3 0.00061346 3.3 0.00061356 0 0.00061348 0 0.00061358 3.3 0.0006135 3.3 0.0006136 0 0.00061352 0 0.0006136199999999999 3.3 0.0006135400000000001 3.3 0.00061364 0 0.0006135600000000001 0 0.00061366 3.3 0.0006135800000000001 3.3 0.00061368 0 0.0006136000000000001 0 0.0006137 3.3 0.00061362 3.3 0.00061372 0 0.00061364 0 0.00061374 3.3 0.00061366 3.3 0.00061376 0 0.00061368 0 0.00061378 3.3 0.0006137 3.3 0.0006138 0 0.00061372 0 0.00061382 3.3 0.00061374 3.3 0.0006138399999999999 0 0.0006137600000000001 0 0.00061386 3.3 0.0006137800000000001 3.3 0.00061388 0 0.0006138000000000001 0 0.0006139 3.3 0.0006138200000000001 3.3 0.00061392 0 0.00061384 0 0.00061394 3.3 0.00061386 3.3 0.00061396 0 0.00061388 0 0.00061398 3.3 0.0006139 3.3 0.000614 0 0.00061392 0 0.00061402 3.3 0.00061394 3.3 0.0006140399999999999 0 0.0006139600000000001 0 0.00061406 3.3 0.0006139800000000001 3.3 0.00061408 0 0.0006140000000000001 0 0.0006141 3.3 0.0006140200000000001 3.3 0.00061412 0 0.00061404 0 0.00061414 3.3 0.00061406 3.3 0.00061416 0 0.00061408 0 0.00061418 3.3 0.0006141 3.3 0.0006142 0 0.00061412 0 0.00061422 3.3 0.00061414 3.3 0.00061424 0 0.00061416 0 0.0006142599999999999 3.3 0.0006141800000000001 3.3 0.00061428 0 0.0006142000000000001 0 0.0006143 3.3 0.0006142200000000001 3.3 0.00061432 0 0.0006142400000000001 0 0.00061434 3.3 0.00061426 3.3 0.00061436 0 0.00061428 0 0.00061438 3.3 0.0006143 3.3 0.0006144 0 0.00061432 0 0.00061442 3.3 0.00061434 3.3 0.00061444 0 0.00061436 0 0.0006144599999999999 3.3 0.0006143800000000001 3.3 0.00061448 0 0.0006144000000000001 0 0.0006145 3.3 0.0006144200000000001 3.3 0.00061452 0 0.0006144400000000001 0 0.00061454 3.3 0.00061446 3.3 0.00061456 0 0.00061448 0 0.00061458 3.3 0.0006145 3.3 0.0006146 0 0.00061452 0 0.00061462 3.3 0.00061454 3.3 0.00061464 0 0.00061456 0 0.00061466 3.3 0.00061458 3.3 0.0006146799999999999 0 0.0006146000000000001 0 0.0006147 3.3 0.0006146200000000001 3.3 0.00061472 0 0.0006146400000000001 0 0.00061474 3.3 0.0006146600000000001 3.3 0.00061476 0 0.00061468 0 0.00061478 3.3 0.0006147 3.3 0.0006148 0 0.00061472 0 0.00061482 3.3 0.00061474 3.3 0.00061484 0 0.00061476 0 0.00061486 3.3 0.00061478 3.3 0.0006148799999999999 0 0.0006148000000000001 0 0.0006149 3.3 0.0006148200000000001 3.3 0.00061492 0 0.0006148400000000001 0 0.00061494 3.3 0.0006148600000000001 3.3 0.00061496 0 0.00061488 0 0.00061498 3.3 0.0006149 3.3 0.000615 0 0.00061492 0 0.00061502 3.3 0.00061494 3.3 0.00061504 0 0.00061496 0 0.00061506 3.3 0.00061498 3.3 0.0006150799999999999 0 0.000615 0 0.0006150999999999999 3.3 0.0006150200000000001 3.3 0.00061512 0 0.0006150400000000001 0 0.00061514 3.3 0.0006150600000000001 3.3 0.00061516 0 0.00061508 0 0.00061518 3.3 0.0006151 3.3 0.0006152 0 0.00061512 0 0.00061522 3.3 0.00061514 3.3 0.00061524 0 0.00061516 0 0.00061526 3.3 0.00061518 3.3 0.00061528 0 0.0006152 0 0.0006152999999999999 3.3 0.0006152200000000001 3.3 0.00061532 0 0.0006152400000000001 0 0.00061534 3.3 0.0006152600000000001 3.3 0.00061536 0 0.0006152800000000001 0 0.00061538 3.3 0.0006153 3.3 0.0006154 0 0.00061532 0 0.00061542 3.3 0.00061534 3.3 0.00061544 0 0.00061536 0 0.00061546 3.3 0.00061538 3.3 0.00061548 0 0.0006154 0 0.0006154999999999999 3.3 0.00061542 3.3 0.0006155199999999999 0 0.0006154400000000001 0 0.00061554 3.3 0.0006154600000000001 3.3 0.00061556 0 0.0006154800000000001 0 0.00061558 3.3 0.0006155 3.3 0.0006156 0 0.00061552 0 0.00061562 3.3 0.00061554 3.3 0.00061564 0 0.00061556 0 0.00061566 3.3 0.00061558 3.3 0.00061568 0 0.0006156 0 0.0006157 3.3 0.00061562 3.3 0.0006157199999999999 0 0.0006156400000000001 0 0.00061574 3.3 0.0006156600000000001 3.3 0.00061576 0 0.0006156800000000001 0 0.00061578 3.3 0.0006157000000000001 3.3 0.0006158 0 0.00061572 0 0.00061582 3.3 0.00061574 3.3 0.00061584 0 0.00061576 0 0.00061586 3.3 0.00061578 3.3 0.00061588 0 0.0006158 0 0.0006159 3.3 0.00061582 3.3 0.0006159199999999999 0 0.00061584 0 0.0006159399999999999 3.3 0.0006158600000000001 3.3 0.00061596 0 0.0006158800000000001 0 0.00061598 3.3 0.0006159000000000001 3.3 0.000616 0 0.00061592 0 0.00061602 3.3 0.00061594 3.3 0.00061604 0 0.00061596 0 0.00061606 3.3 0.00061598 3.3 0.00061608 0 0.000616 0 0.0006161 3.3 0.00061602 3.3 0.00061612 0 0.00061604 0 0.0006161399999999999 3.3 0.0006160600000000001 3.3 0.00061616 0 0.0006160800000000001 0 0.00061618 3.3 0.0006161000000000001 3.3 0.0006162 0 0.0006161200000000001 0 0.00061622 3.3 0.00061614 3.3 0.00061624 0 0.00061616 0 0.00061626 3.3 0.00061618 3.3 0.00061628 0 0.0006162 0 0.0006163 3.3 0.00061622 3.3 0.00061632 0 0.00061624 0 0.0006163399999999999 3.3 0.0006162600000000001 3.3 0.00061636 0 0.0006162800000000001 0 0.00061638 3.3 0.0006163000000000001 3.3 0.0006164 0 0.0006163200000000001 0 0.00061642 3.3 0.00061634 3.3 0.00061644 0 0.00061636 0 0.00061646 3.3 0.00061638 3.3 0.00061648 0 0.0006164 0 0.0006165 3.3 0.00061642 3.3 0.00061652 0 0.00061644 0 0.00061654 3.3 0.00061646 3.3 0.0006165599999999999 0 0.0006164800000000001 0 0.00061658 3.3 0.0006165000000000001 3.3 0.0006166 0 0.0006165200000000001 0 0.00061662 3.3 0.0006165400000000001 3.3 0.00061664 0 0.00061656 0 0.00061666 3.3 0.00061658 3.3 0.00061668 0 0.0006166 0 0.0006167 3.3 0.00061662 3.3 0.00061672 0 0.00061664 0 0.00061674 3.3 0.00061666 3.3 0.0006167599999999999 0 0.0006166800000000001 0 0.00061678 3.3 0.0006167000000000001 3.3 0.0006168 0 0.0006167200000000001 0 0.00061682 3.3 0.0006167400000000001 3.3 0.00061684 0 0.00061676 0 0.00061686 3.3 0.00061678 3.3 0.00061688 0 0.0006168 0 0.0006169 3.3 0.00061682 3.3 0.00061692 0 0.00061684 0 0.00061694 3.3 0.00061686 3.3 0.00061696 0 0.00061688 0 0.0006169799999999999 3.3 0.0006169000000000001 3.3 0.000617 0 0.0006169200000000001 0 0.00061702 3.3 0.0006169400000000001 3.3 0.00061704 0 0.0006169600000000001 0 0.00061706 3.3 0.00061698 3.3 0.00061708 0 0.000617 0 0.0006171 3.3 0.00061702 3.3 0.00061712 0 0.00061704 0 0.00061714 3.3 0.00061706 3.3 0.00061716 0 0.00061708 0 0.0006171799999999999 3.3 0.0006171000000000001 3.3 0.0006172 0 0.0006171200000000001 0 0.00061722 3.3 0.0006171400000000001 3.3 0.00061724 0 0.0006171600000000001 0 0.00061726 3.3 0.00061718 3.3 0.00061728 0 0.0006172 0 0.0006173 3.3 0.00061722 3.3 0.00061732 0 0.00061724 0 0.00061734 3.3 0.00061726 3.3 0.00061736 0 0.00061728 0 0.00061738 3.3 0.0006173 3.3 0.0006173999999999999 0 0.0006173200000000001 0 0.00061742 3.3 0.0006173400000000001 3.3 0.00061744 0 0.0006173600000000001 0 0.00061746 3.3 0.0006173800000000001 3.3 0.00061748 0 0.0006174 0 0.0006175 3.3 0.00061742 3.3 0.00061752 0 0.00061744 0 0.00061754 3.3 0.00061746 3.3 0.00061756 0 0.00061748 0 0.00061758 3.3 0.0006175 3.3 0.0006175999999999999 0 0.0006175200000000001 0 0.00061762 3.3 0.0006175400000000001 3.3 0.00061764 0 0.0006175600000000001 0 0.00061766 3.3 0.0006175800000000001 3.3 0.00061768 0 0.0006176 0 0.0006177 3.3 0.00061762 3.3 0.00061772 0 0.00061764 0 0.00061774 3.3 0.00061766 3.3 0.00061776 0 0.00061768 0 0.00061778 3.3 0.0006177 3.3 0.0006178 0 0.00061772 0 0.0006178199999999999 3.3 0.0006177400000000001 3.3 0.00061784 0 0.0006177600000000001 0 0.00061786 3.3 0.0006177800000000001 3.3 0.00061788 0 0.0006178000000000001 0 0.0006179 3.3 0.00061782 3.3 0.00061792 0 0.00061784 0 0.00061794 3.3 0.00061786 3.3 0.00061796 0 0.00061788 0 0.00061798 3.3 0.0006179 3.3 0.000618 0 0.00061792 0 0.0006180199999999999 3.3 0.0006179400000000001 3.3 0.00061804 0 0.0006179600000000001 0 0.00061806 3.3 0.0006179800000000001 3.3 0.00061808 0 0.0006180000000000001 0 0.0006181 3.3 0.00061802 3.3 0.00061812 0 0.00061804 0 0.00061814 3.3 0.00061806 3.3 0.00061816 0 0.00061808 0 0.00061818 3.3 0.0006181 3.3 0.0006182 0 0.00061812 0 0.0006182199999999999 3.3 0.00061814 3.3 0.0006182399999999999 0 0.0006181600000000001 0 0.00061826 3.3 0.0006181800000000001 3.3 0.00061828 0 0.0006182000000000001 0 0.0006183 3.3 0.00061822 3.3 0.00061832 0 0.00061824 0 0.00061834 3.3 0.00061826 3.3 0.00061836 0 0.00061828 0 0.00061838 3.3 0.0006183 3.3 0.0006184 0 0.00061832 0 0.00061842 3.3 0.00061834 3.3 0.0006184399999999999 0 0.0006183600000000001 0 0.00061846 3.3 0.0006183800000000001 3.3 0.00061848 0 0.0006184000000000001 0 0.0006185 3.3 0.0006184200000000001 3.3 0.00061852 0 0.00061844 0 0.00061854 3.3 0.00061846 3.3 0.00061856 0 0.00061848 0 0.00061858 3.3 0.0006185 3.3 0.0006186 0 0.00061852 0 0.00061862 3.3 0.00061854 3.3 0.0006186399999999999 0 0.00061856 0 0.0006186599999999999 3.3 0.0006185800000000001 3.3 0.00061868 0 0.0006186000000000001 0 0.0006187 3.3 0.0006186200000000001 3.3 0.00061872 0 0.00061864 0 0.00061874 3.3 0.00061866 3.3 0.00061876 0 0.00061868 0 0.00061878 3.3 0.0006187 3.3 0.0006188 0 0.00061872 0 0.00061882 3.3 0.00061874 3.3 0.00061884 0 0.00061876 0 0.0006188599999999999 3.3 0.0006187800000000001 3.3 0.00061888 0 0.0006188000000000001 0 0.0006189 3.3 0.0006188200000000001 3.3 0.00061892 0 0.0006188400000000001 0 0.00061894 3.3 0.00061886 3.3 0.00061896 0 0.00061888 0 0.00061898 3.3 0.0006189 3.3 0.000619 0 0.00061892 0 0.00061902 3.3 0.00061894 3.3 0.00061904 0 0.00061896 0 0.0006190599999999999 3.3 0.00061898 3.3 0.0006190799999999999 0 0.0006190000000000001 0 0.0006191 3.3 0.0006190200000000001 3.3 0.00061912 0 0.0006190400000000001 0 0.00061914 3.3 0.00061906 3.3 0.00061916 0 0.00061908 0 0.00061918 3.3 0.0006191 3.3 0.0006192 0 0.00061912 0 0.00061922 3.3 0.00061914 3.3 0.00061924 0 0.00061916 0 0.00061926 3.3 0.00061918 3.3 0.0006192799999999999 0 0.0006192000000000001 0 0.0006193 3.3 0.0006192200000000001 3.3 0.00061932 0 0.0006192400000000001 0 0.00061934 3.3 0.0006192600000000001 3.3 0.00061936 0 0.00061928 0 0.00061938 3.3 0.0006193 3.3 0.0006194 0 0.00061932 0 0.00061942 3.3 0.00061934 3.3 0.00061944 0 0.00061936 0 0.00061946 3.3 0.00061938 3.3 0.0006194799999999999 0 0.0006194 0 0.0006194999999999999 3.3 0.0006194200000000001 3.3 0.00061952 0 0.0006194400000000001 0 0.00061954 3.3 0.0006194600000000001 3.3 0.00061956 0 0.00061948 0 0.00061958 3.3 0.0006195 3.3 0.0006196 0 0.00061952 0 0.00061962 3.3 0.00061954 3.3 0.00061964 0 0.00061956 0 0.00061966 3.3 0.00061958 3.3 0.00061968 0 0.0006196 0 0.0006196999999999999 3.3 0.0006196200000000001 3.3 0.00061972 0 0.0006196400000000001 0 0.00061974 3.3 0.0006196600000000001 3.3 0.00061976 0 0.0006196800000000001 0 0.00061978 3.3 0.0006197 3.3 0.0006198 0 0.00061972 0 0.00061982 3.3 0.00061974 3.3 0.00061984 0 0.00061976 0 0.00061986 3.3 0.00061978 3.3 0.00061988 0 0.0006198 0 0.0006198999999999999 3.3 0.0006198200000000001 3.3 0.00061992 0 0.0006198400000000001 0 0.00061994 3.3 0.0006198600000000001 3.3 0.00061996 0 0.0006198800000000001 0 0.00061998 3.3 0.0006199 3.3 0.00062 0 0.00061992 0 0.00062002 3.3 0.00061994 3.3 0.00062004 0 0.00061996 0 0.00062006 3.3 0.00061998 3.3 0.00062008 0 0.00062 0 0.0006201 3.3 0.00062002 3.3 0.0006201199999999999 0 0.0006200400000000001 0 0.00062014 3.3 0.0006200600000000001 3.3 0.00062016 0 0.0006200800000000001 0 0.00062018 3.3 0.0006201000000000001 3.3 0.0006202 0 0.00062012 0 0.00062022 3.3 0.00062014 3.3 0.00062024 0 0.00062016 0 0.00062026 3.3 0.00062018 3.3 0.00062028 0 0.0006202 0 0.0006203 3.3 0.00062022 3.3 0.0006203199999999999 0 0.0006202400000000001 0 0.00062034 3.3 0.0006202600000000001 3.3 0.00062036 0 0.0006202800000000001 0 0.00062038 3.3 0.0006203000000000001 3.3 0.0006204 0 0.00062032 0 0.00062042 3.3 0.00062034 3.3 0.00062044 0 0.00062036 0 0.00062046 3.3 0.00062038 3.3 0.00062048 0 0.0006204 0 0.0006205 3.3 0.00062042 3.3 0.00062052 0 0.00062044 0 0.0006205399999999999 3.3 0.0006204600000000001 3.3 0.00062056 0 0.0006204800000000001 0 0.00062058 3.3 0.0006205000000000001 3.3 0.0006206 0 0.0006205200000000001 0 0.00062062 3.3 0.00062054 3.3 0.00062064 0 0.00062056 0 0.00062066 3.3 0.00062058 3.3 0.00062068 0 0.0006206 0 0.0006207 3.3 0.00062062 3.3 0.00062072 0 0.00062064 0 0.0006207399999999999 3.3 0.0006206600000000001 3.3 0.00062076 0 0.0006206800000000001 0 0.00062078 3.3 0.0006207000000000001 3.3 0.0006208 0 0.0006207200000000001 0 0.00062082 3.3 0.00062074 3.3 0.00062084 0 0.00062076 0 0.00062086 3.3 0.00062078 3.3 0.00062088 0 0.0006208 0 0.0006209 3.3 0.00062082 3.3 0.00062092 0 0.00062084 0 0.00062094 3.3 0.00062086 3.3 0.0006209599999999999 0 0.0006208800000000001 0 0.00062098 3.3 0.0006209000000000001 3.3 0.000621 0 0.0006209200000000001 0 0.00062102 3.3 0.0006209400000000001 3.3 0.00062104 0 0.00062096 0 0.00062106 3.3 0.00062098 3.3 0.00062108 0 0.000621 0 0.0006211 3.3 0.00062102 3.3 0.00062112 0 0.00062104 0 0.00062114 3.3 0.00062106 3.3 0.0006211599999999999 0 0.0006210800000000001 0 0.00062118 3.3 0.0006211000000000001 3.3 0.0006212 0 0.0006211200000000001 0 0.00062122 3.3 0.0006211400000000001 3.3 0.00062124 0 0.00062116 0 0.00062126 3.3 0.00062118 3.3 0.00062128 0 0.0006212 0 0.0006213 3.3 0.00062122 3.3 0.00062132 0 0.00062124 0 0.00062134 3.3 0.00062126 3.3 0.00062136 0 0.00062128 0 0.0006213799999999999 3.3 0.0006213000000000001 3.3 0.0006214 0 0.0006213200000000001 0 0.00062142 3.3 0.0006213400000000001 3.3 0.00062144 0 0.0006213600000000001 0 0.00062146 3.3 0.00062138 3.3 0.00062148 0 0.0006214 0 0.0006215 3.3 0.00062142 3.3 0.00062152 0 0.00062144 0 0.00062154 3.3 0.00062146 3.3 0.00062156 0 0.00062148 0 0.0006215799999999999 3.3 0.0006215000000000001 3.3 0.0006216 0 0.0006215200000000001 0 0.00062162 3.3 0.0006215400000000001 3.3 0.00062164 0 0.0006215600000000001 0 0.00062166 3.3 0.00062158 3.3 0.00062168 0 0.0006216 0 0.0006217 3.3 0.00062162 3.3 0.00062172 0 0.00062164 0 0.00062174 3.3 0.00062166 3.3 0.00062176 0 0.00062168 0 0.0006217799999999999 3.3 0.0006217 3.3 0.0006217999999999999 0 0.0006217200000000001 0 0.00062182 3.3 0.0006217400000000001 3.3 0.00062184 0 0.0006217600000000001 0 0.00062186 3.3 0.00062178 3.3 0.00062188 0 0.0006218 0 0.0006219 3.3 0.00062182 3.3 0.00062192 0 0.00062184 0 0.00062194 3.3 0.00062186 3.3 0.00062196 0 0.00062188 0 0.00062198 3.3 0.0006219 3.3 0.0006219999999999999 0 0.0006219200000000001 0 0.00062202 3.3 0.0006219400000000001 3.3 0.00062204 0 0.0006219600000000001 0 0.00062206 3.3 0.0006219800000000001 3.3 0.00062208 0 0.000622 0 0.0006221 3.3 0.00062202 3.3 0.00062212 0 0.00062204 0 0.00062214 3.3 0.00062206 3.3 0.00062216 0 0.00062208 0 0.00062218 3.3 0.0006221 3.3 0.0006221999999999999 0 0.00062212 0 0.0006222199999999999 3.3 0.0006221400000000001 3.3 0.00062224 0 0.0006221600000000001 0 0.00062226 3.3 0.0006221800000000001 3.3 0.00062228 0 0.0006222 0 0.0006223 3.3 0.00062222 3.3 0.00062232 0 0.00062224 0 0.00062234 3.3 0.00062226 3.3 0.00062236 0 0.00062228 0 0.00062238 3.3 0.0006223 3.3 0.0006224 0 0.00062232 0 0.0006224199999999999 3.3 0.0006223400000000001 3.3 0.00062244 0 0.0006223600000000001 0 0.00062246 3.3 0.0006223800000000001 3.3 0.00062248 0 0.0006224000000000001 0 0.0006225 3.3 0.00062242 3.3 0.00062252 0 0.00062244 0 0.00062254 3.3 0.00062246 3.3 0.00062256 0 0.00062248 0 0.00062258 3.3 0.0006225 3.3 0.0006226 0 0.00062252 0 0.0006226199999999999 3.3 0.00062254 3.3 0.0006226399999999999 0 0.0006225600000000001 0 0.00062266 3.3 0.0006225800000000001 3.3 0.00062268 0 0.0006226000000000001 0 0.0006227 3.3 0.00062262 3.3 0.00062272 0 0.00062264 0 0.00062274 3.3 0.00062266 3.3 0.00062276 0 0.00062268 0 0.00062278 3.3 0.0006227 3.3 0.0006228 0 0.00062272 0 0.00062282 3.3 0.00062274 3.3 0.0006228399999999999 0 0.0006227600000000001 0 0.00062286 3.3 0.0006227800000000001 3.3 0.00062288 0 0.0006228000000000001 0 0.0006229 3.3 0.0006228200000000001 3.3 0.00062292 0 0.00062284 0 0.00062294 3.3 0.00062286 3.3 0.00062296 0 0.00062288 0 0.00062298 3.3 0.0006229 3.3 0.000623 0 0.00062292 0 0.00062302 3.3 0.00062294 3.3 0.0006230399999999999 0 0.00062296 0 0.0006230599999999999 3.3 0.0006229800000000001 3.3 0.00062308 0 0.0006230000000000001 0 0.0006231 3.3 0.0006230200000000001 3.3 0.00062312 0 0.00062304 0 0.00062314 3.3 0.00062306 3.3 0.00062316 0 0.00062308 0 0.00062318 3.3 0.0006231 3.3 0.0006232 0 0.00062312 0 0.00062322 3.3 0.00062314 3.3 0.00062324 0 0.00062316 0 0.0006232599999999999 3.3 0.0006231800000000001 3.3 0.00062328 0 0.0006232000000000001 0 0.0006233 3.3 0.0006232200000000001 3.3 0.00062332 0 0.0006232400000000001 0 0.00062334 3.3 0.00062326 3.3 0.00062336 0 0.00062328 0 0.00062338 3.3 0.0006233 3.3 0.0006234 0 0.00062332 0 0.00062342 3.3 0.00062334 3.3 0.00062344 0 0.00062336 0 0.0006234599999999999 3.3 0.0006233800000000001 3.3 0.00062348 0 0.0006234000000000001 0 0.0006235 3.3 0.0006234200000000001 3.3 0.00062352 0 0.0006234400000000001 0 0.00062354 3.3 0.00062346 3.3 0.00062356 0 0.00062348 0 0.00062358 3.3 0.0006235 3.3 0.0006236 0 0.00062352 0 0.00062362 3.3 0.00062354 3.3 0.00062364 0 0.00062356 0 0.00062366 3.3 0.00062358 3.3 0.0006236799999999999 0 0.0006236000000000001 0 0.0006237 3.3 0.0006236200000000001 3.3 0.00062372 0 0.0006236400000000001 0 0.00062374 3.3 0.0006236600000000001 3.3 0.00062376 0 0.00062368 0 0.00062378 3.3 0.0006237 3.3 0.0006238 0 0.00062372 0 0.00062382 3.3 0.00062374 3.3 0.00062384 0 0.00062376 0 0.00062386 3.3 0.00062378 3.3 0.0006238799999999999 0 0.0006238000000000001 0 0.0006239 3.3 0.0006238200000000001 3.3 0.00062392 0 0.0006238400000000001 0 0.00062394 3.3 0.0006238600000000001 3.3 0.00062396 0 0.00062388 0 0.00062398 3.3 0.0006239 3.3 0.000624 0 0.00062392 0 0.00062402 3.3 0.00062394 3.3 0.00062404 0 0.00062396 0 0.00062406 3.3 0.00062398 3.3 0.00062408 0 0.000624 0 0.0006240999999999999 3.3 0.0006240200000000001 3.3 0.00062412 0 0.0006240400000000001 0 0.00062414 3.3 0.0006240600000000001 3.3 0.00062416 0 0.0006240800000000001 0 0.00062418 3.3 0.0006241 3.3 0.0006242 0 0.00062412 0 0.00062422 3.3 0.00062414 3.3 0.00062424 0 0.00062416 0 0.00062426 3.3 0.00062418 3.3 0.00062428 0 0.0006242 0 0.0006242999999999999 3.3 0.0006242200000000001 3.3 0.00062432 0 0.0006242400000000001 0 0.00062434 3.3 0.0006242600000000001 3.3 0.00062436 0 0.0006242800000000001 0 0.00062438 3.3 0.0006243 3.3 0.0006244 0 0.00062432 0 0.00062442 3.3 0.00062434 3.3 0.00062444 0 0.00062436 0 0.00062446 3.3 0.00062438 3.3 0.00062448 0 0.0006244 0 0.0006245 3.3 0.00062442 3.3 0.0006245199999999999 0 0.0006244400000000001 0 0.00062454 3.3 0.0006244600000000001 3.3 0.00062456 0 0.0006244800000000001 0 0.00062458 3.3 0.0006245000000000001 3.3 0.0006246 0 0.00062452 0 0.00062462 3.3 0.00062454 3.3 0.00062464 0 0.00062456 0 0.00062466 3.3 0.00062458 3.3 0.00062468 0 0.0006246 0 0.0006247 3.3 0.00062462 3.3 0.0006247199999999999 0 0.0006246400000000001 0 0.00062474 3.3 0.0006246600000000001 3.3 0.00062476 0 0.0006246800000000001 0 0.00062478 3.3 0.0006247000000000001 3.3 0.0006248 0 0.00062472 0 0.00062482 3.3 0.00062474 3.3 0.00062484 0 0.00062476 0 0.00062486 3.3 0.00062478 3.3 0.00062488 0 0.0006248 0 0.0006249 3.3 0.00062482 3.3 0.00062492 0 0.00062484 0 0.0006249399999999999 3.3 0.0006248600000000001 3.3 0.00062496 0 0.0006248800000000001 0 0.00062498 3.3 0.0006249000000000001 3.3 0.000625 0 0.0006249200000000001 0 0.00062502 3.3 0.00062494 3.3 0.00062504 0 0.00062496 0 0.00062506 3.3 0.00062498 3.3 0.00062508 0 0.000625 0 0.0006251 3.3 0.00062502 3.3 0.00062512 0 0.00062504 0 0.0006251399999999999 3.3 0.0006250600000000001 3.3 0.00062516 0 0.0006250800000000001 0 0.00062518 3.3 0.0006251000000000001 3.3 0.0006252 0 0.0006251200000000001 0 0.00062522 3.3 0.00062514 3.3 0.00062524 0 0.00062516 0 0.00062526 3.3 0.00062518 3.3 0.00062528 0 0.0006252 0 0.0006253 3.3 0.00062522 3.3 0.00062532 0 0.00062524 0 0.0006253399999999999 3.3 0.00062526 3.3 0.0006253599999999999 0 0.0006252800000000001 0 0.00062538 3.3 0.0006253000000000001 3.3 0.0006254 0 0.0006253200000000001 0 0.00062542 3.3 0.00062534 3.3 0.00062544 0 0.00062536 0 0.00062546 3.3 0.00062538 3.3 0.00062548 0 0.0006254 0 0.0006255 3.3 0.00062542 3.3 0.00062552 0 0.00062544 0 0.00062554 3.3 0.00062546 3.3 0.0006255599999999999 0 0.0006254800000000001 0 0.00062558 3.3 0.0006255000000000001 3.3 0.0006256 0 0.0006255200000000001 0 0.00062562 3.3 0.0006255400000000001 3.3 0.00062564 0 0.00062556 0 0.00062566 3.3 0.00062558 3.3 0.00062568 0 0.0006256 0 0.0006257 3.3 0.00062562 3.3 0.00062572 0 0.00062564 0 0.00062574 3.3 0.00062566 3.3 0.0006257599999999999 0 0.00062568 0 0.0006257799999999999 3.3 0.0006257000000000001 3.3 0.0006258 0 0.0006257200000000001 0 0.00062582 3.3 0.0006257400000000001 3.3 0.00062584 0 0.00062576 0 0.00062586 3.3 0.00062578 3.3 0.00062588 0 0.0006258 0 0.0006259 3.3 0.00062582 3.3 0.00062592 0 0.00062584 0 0.00062594 3.3 0.00062586 3.3 0.00062596 0 0.00062588 0 0.0006259799999999999 3.3 0.0006259000000000001 3.3 0.000626 0 0.0006259200000000001 0 0.00062602 3.3 0.0006259400000000001 3.3 0.00062604 0 0.0006259600000000001 0 0.00062606 3.3 0.00062598 3.3 0.00062608 0 0.000626 0 0.0006261 3.3 0.00062602 3.3 0.00062612 0 0.00062604 0 0.00062614 3.3 0.00062606 3.3 0.00062616 0 0.00062608 0 0.0006261799999999999 3.3 0.0006261 3.3 0.0006261999999999999 0 0.0006261200000000001 0 0.00062622 3.3 0.0006261400000000001 3.3 0.00062624 0 0.0006261600000000001 0 0.00062626 3.3 0.00062618 3.3 0.00062628 0 0.0006262 0 0.0006263 3.3 0.00062622 3.3 0.00062632 0 0.00062624 0 0.00062634 3.3 0.00062626 3.3 0.00062636 0 0.00062628 0 0.00062638 3.3 0.0006263 3.3 0.0006263999999999999 0 0.0006263200000000001 0 0.00062642 3.3 0.0006263400000000001 3.3 0.00062644 0 0.0006263600000000001 0 0.00062646 3.3 0.0006263800000000001 3.3 0.00062648 0 0.0006264 0 0.0006265 3.3 0.00062642 3.3 0.00062652 0 0.00062644 0 0.00062654 3.3 0.00062646 3.3 0.00062656 0 0.00062648 0 0.00062658 3.3 0.0006265 3.3 0.0006265999999999999 0 0.0006265200000000001 0 0.00062662 3.3 0.0006265400000000001 3.3 0.00062664 0 0.0006265600000000001 0 0.00062666 3.3 0.0006265800000000001 3.3 0.00062668 0 0.0006266 0 0.0006267 3.3 0.00062662 3.3 0.00062672 0 0.00062664 0 0.00062674 3.3 0.00062666 3.3 0.00062676 0 0.00062668 0 0.00062678 3.3 0.0006267 3.3 0.0006268 0 0.00062672 0 0.0006268199999999999 3.3 0.0006267400000000001 3.3 0.00062684 0 0.0006267600000000001 0 0.00062686 3.3 0.0006267800000000001 3.3 0.00062688 0 0.0006268000000000001 0 0.0006269 3.3 0.00062682 3.3 0.00062692 0 0.00062684 0 0.00062694 3.3 0.00062686 3.3 0.00062696 0 0.00062688 0 0.00062698 3.3 0.0006269 3.3 0.000627 0 0.00062692 0 0.0006270199999999999 3.3 0.0006269400000000001 3.3 0.00062704 0 0.0006269600000000001 0 0.00062706 3.3 0.0006269800000000001 3.3 0.00062708 0 0.0006270000000000001 0 0.0006271 3.3 0.00062702 3.3 0.00062712 0 0.00062704 0 0.00062714 3.3 0.00062706 3.3 0.00062716 0 0.00062708 0 0.00062718 3.3 0.0006271 3.3 0.0006272 0 0.00062712 0 0.00062722 3.3 0.00062714 3.3 0.0006272399999999999 0 0.0006271600000000001 0 0.00062726 3.3 0.0006271800000000001 3.3 0.00062728 0 0.0006272000000000001 0 0.0006273 3.3 0.0006272200000000001 3.3 0.00062732 0 0.00062724 0 0.00062734 3.3 0.00062726 3.3 0.00062736 0 0.00062728 0 0.00062738 3.3 0.0006273 3.3 0.0006274 0 0.00062732 0 0.00062742 3.3 0.00062734 3.3 0.0006274399999999999 0 0.0006273600000000001 0 0.00062746 3.3 0.0006273800000000001 3.3 0.00062748 0 0.0006274000000000001 0 0.0006275 3.3 0.0006274200000000001 3.3 0.00062752 0 0.00062744 0 0.00062754 3.3 0.00062746 3.3 0.00062756 0 0.00062748 0 0.00062758 3.3 0.0006275 3.3 0.0006276 0 0.00062752 0 0.00062762 3.3 0.00062754 3.3 0.00062764 0 0.00062756 0 0.0006276599999999999 3.3 0.0006275800000000001 3.3 0.00062768 0 0.0006276000000000001 0 0.0006277 3.3 0.0006276200000000001 3.3 0.00062772 0 0.0006276400000000001 0 0.00062774 3.3 0.00062766 3.3 0.00062776 0 0.00062768 0 0.00062778 3.3 0.0006277 3.3 0.0006278 0 0.00062772 0 0.00062782 3.3 0.00062774 3.3 0.00062784 0 0.00062776 0 0.0006278599999999999 3.3 0.0006277800000000001 3.3 0.00062788 0 0.0006278000000000001 0 0.0006279 3.3 0.0006278200000000001 3.3 0.00062792 0 0.0006278400000000001 0 0.00062794 3.3 0.00062786 3.3 0.00062796 0 0.00062788 0 0.00062798 3.3 0.0006279 3.3 0.000628 0 0.00062792 0 0.00062802 3.3 0.00062794 3.3 0.00062804 0 0.00062796 0 0.00062806 3.3 0.00062798 3.3 0.0006280799999999999 0 0.0006280000000000001 0 0.0006281 3.3 0.0006280200000000001 3.3 0.00062812 0 0.0006280400000000001 0 0.00062814 3.3 0.0006280600000000001 3.3 0.00062816 0 0.00062808 0 0.00062818 3.3 0.0006281 3.3 0.0006282 0 0.00062812 0 0.00062822 3.3 0.00062814 3.3 0.00062824 0 0.00062816 0 0.00062826 3.3 0.00062818 3.3 0.0006282799999999999 0 0.0006282000000000001 0 0.0006283 3.3 0.0006282200000000001 3.3 0.00062832 0 0.0006282400000000001 0 0.00062834 3.3 0.0006282600000000001 3.3 0.00062836 0 0.00062828 0 0.00062838 3.3 0.0006283 3.3 0.0006284 0 0.00062832 0 0.00062842 3.3 0.00062834 3.3 0.00062844 0 0.00062836 0 0.00062846 3.3 0.00062838 3.3 0.00062848 0 0.0006284 0 0.0006284999999999999 3.3 0.0006284200000000001 3.3 0.00062852 0 0.0006284400000000001 0 0.00062854 3.3 0.0006284600000000001 3.3 0.00062856 0 0.0006284800000000001 0 0.00062858 3.3 0.0006285 3.3 0.0006286 0 0.00062852 0 0.00062862 3.3 0.00062854 3.3 0.00062864 0 0.00062856 0 0.00062866 3.3 0.00062858 3.3 0.00062868 0 0.0006286 0 0.0006286999999999999 3.3 0.0006286200000000001 3.3 0.00062872 0 0.0006286400000000001 0 0.00062874 3.3 0.0006286600000000001 3.3 0.00062876 0 0.0006286800000000001 0 0.00062878 3.3 0.0006287 3.3 0.0006288 0 0.00062872 0 0.00062882 3.3 0.00062874 3.3 0.00062884 0 0.00062876 0 0.00062886 3.3 0.00062878 3.3 0.00062888 0 0.0006288 0 0.0006288999999999999 3.3 0.00062882 3.3 0.0006289199999999999 0 0.0006288400000000001 0 0.00062894 3.3 0.0006288600000000001 3.3 0.00062896 0 0.0006288800000000001 0 0.00062898 3.3 0.0006289 3.3 0.000629 0 0.00062892 0 0.00062902 3.3 0.00062894 3.3 0.00062904 0 0.00062896 0 0.00062906 3.3 0.00062898 3.3 0.00062908 0 0.000629 0 0.0006291 3.3 0.00062902 3.3 0.0006291199999999999 0 0.0006290400000000001 0 0.00062914 3.3 0.0006290600000000001 3.3 0.00062916 0 0.0006290800000000001 0 0.00062918 3.3 0.0006291000000000001 3.3 0.0006292 0 0.00062912 0 0.00062922 3.3 0.00062914 3.3 0.00062924 0 0.00062916 0 0.00062926 3.3 0.00062918 3.3 0.00062928 0 0.0006292 0 0.0006293 3.3 0.00062922 3.3 0.0006293199999999999 0 0.00062924 0 0.0006293399999999999 3.3 0.0006292600000000001 3.3 0.00062936 0 0.0006292800000000001 0 0.00062938 3.3 0.0006293000000000001 3.3 0.0006294 0 0.00062932 0 0.00062942 3.3 0.00062934 3.3 0.00062944 0 0.00062936 0 0.00062946 3.3 0.00062938 3.3 0.00062948 0 0.0006294 0 0.0006295 3.3 0.00062942 3.3 0.00062952 0 0.00062944 0 0.0006295399999999999 3.3 0.0006294600000000001 3.3 0.00062956 0 0.0006294800000000001 0 0.00062958 3.3 0.0006295000000000001 3.3 0.0006296 0 0.0006295200000000001 0 0.00062962 3.3 0.00062954 3.3 0.00062964 0 0.00062956 0 0.00062966 3.3 0.00062958 3.3 0.00062968 0 0.0006296 0 0.0006297 3.3 0.00062962 3.3 0.00062972 0 0.00062964 0 0.0006297399999999999 3.3 0.00062966 3.3 0.0006297599999999999 0 0.0006296800000000001 0 0.00062978 3.3 0.0006297000000000001 3.3 0.0006298 0 0.0006297200000000001 0 0.00062982 3.3 0.00062974 3.3 0.00062984 0 0.00062976 0 0.00062986 3.3 0.00062978 3.3 0.00062988 0 0.0006298 0 0.0006299 3.3 0.00062982 3.3 0.00062992 0 0.00062984 0 0.00062994 3.3 0.00062986 3.3 0.0006299599999999999 0 0.0006298800000000001 0 0.00062998 3.3 0.0006299000000000001 3.3 0.00063 0 0.0006299200000000001 0 0.00063002 3.3 0.0006299400000000001 3.3 0.00063004 0 0.00062996 0 0.00063006 3.3 0.00062998 3.3 0.00063008 0 0.00063 0 0.0006301 3.3 0.00063002 3.3 0.00063012 0 0.00063004 0 0.00063014 3.3 0.00063006 3.3 0.0006301599999999999 0 0.0006300800000000001 0 0.00063018 3.3 0.0006301000000000001 3.3 0.0006302 0 0.0006301200000000001 0 0.00063022 3.3 0.0006301400000000001 3.3 0.00063024 0 0.00063016 0 0.00063026 3.3 0.00063018 3.3 0.00063028 0 0.0006302 0 0.0006303 3.3 0.00063022 3.3 0.00063032 0 0.00063024 0 0.00063034 3.3 0.00063026 3.3 0.00063036 0 0.00063028 0 0.0006303799999999999 3.3 0.0006303000000000001 3.3 0.0006304 0 0.0006303200000000001 0 0.00063042 3.3 0.0006303400000000001 3.3 0.00063044 0 0.0006303600000000001 0 0.00063046 3.3 0.00063038 3.3 0.00063048 0 0.0006304 0 0.0006305 3.3 0.00063042 3.3 0.00063052 0 0.00063044 0 0.00063054 3.3 0.00063046 3.3 0.00063056 0 0.00063048 0 0.0006305799999999999 3.3 0.0006305000000000001 3.3 0.0006306 0 0.0006305200000000001 0 0.00063062 3.3 0.0006305400000000001 3.3 0.00063064 0 0.0006305600000000001 0 0.00063066 3.3 0.00063058 3.3 0.00063068 0 0.0006306 0 0.0006307 3.3 0.00063062 3.3 0.00063072 0 0.00063064 0 0.00063074 3.3 0.00063066 3.3 0.00063076 0 0.00063068 0 0.00063078 3.3 0.0006307 3.3 0.0006307999999999999 0 0.0006307200000000001 0 0.00063082 3.3 0.0006307400000000001 3.3 0.00063084 0 0.0006307600000000001 0 0.00063086 3.3 0.0006307800000000001 3.3 0.00063088 0 0.0006308 0 0.0006309 3.3 0.00063082 3.3 0.00063092 0 0.00063084 0 0.00063094 3.3 0.00063086 3.3 0.00063096 0 0.00063088 0 0.00063098 3.3 0.0006309 3.3 0.0006309999999999999 0 0.0006309200000000001 0 0.00063102 3.3 0.0006309400000000001 3.3 0.00063104 0 0.0006309600000000001 0 0.00063106 3.3 0.0006309800000000001 3.3 0.00063108 0 0.000631 0 0.0006311 3.3 0.00063102 3.3 0.00063112 0 0.00063104 0 0.00063114 3.3 0.00063106 3.3 0.00063116 0 0.00063108 0 0.00063118 3.3 0.0006311 3.3 0.0006312 0 0.00063112 0 0.0006312199999999999 3.3 0.0006311400000000001 3.3 0.00063124 0 0.0006311600000000001 0 0.00063126 3.3 0.0006311800000000001 3.3 0.00063128 0 0.0006312000000000001 0 0.0006313 3.3 0.00063122 3.3 0.00063132 0 0.00063124 0 0.00063134 3.3 0.00063126 3.3 0.00063136 0 0.00063128 0 0.00063138 3.3 0.0006313 3.3 0.0006314 0 0.00063132 0 0.0006314199999999999 3.3 0.0006313400000000001 3.3 0.00063144 0 0.0006313600000000001 0 0.00063146 3.3 0.0006313800000000001 3.3 0.00063148 0 0.0006314000000000001 0 0.0006315 3.3 0.00063142 3.3 0.00063152 0 0.00063144 0 0.00063154 3.3 0.00063146 3.3 0.00063156 0 0.00063148 0 0.00063158 3.3 0.0006315 3.3 0.0006316 0 0.00063152 0 0.00063162 3.3 0.00063154 3.3 0.0006316399999999999 0 0.0006315600000000001 0 0.00063166 3.3 0.0006315800000000001 3.3 0.00063168 0 0.0006316000000000001 0 0.0006317 3.3 0.0006316200000000001 3.3 0.00063172 0 0.00063164 0 0.00063174 3.3 0.00063166 3.3 0.00063176 0 0.00063168 0 0.00063178 3.3 0.0006317 3.3 0.0006318 0 0.00063172 0 0.00063182 3.3 0.00063174 3.3 0.0006318399999999999 0 0.0006317600000000001 0 0.00063186 3.3 0.0006317800000000001 3.3 0.00063188 0 0.0006318000000000001 0 0.0006319 3.3 0.0006318200000000001 3.3 0.00063192 0 0.00063184 0 0.00063194 3.3 0.00063186 3.3 0.00063196 0 0.00063188 0 0.00063198 3.3 0.0006319 3.3 0.000632 0 0.00063192 0 0.00063202 3.3 0.00063194 3.3 0.0006320399999999999 0 0.00063196 0 0.0006320599999999999 3.3 0.0006319800000000001 3.3 0.00063208 0 0.0006320000000000001 0 0.0006321 3.3 0.0006320200000000001 3.3 0.00063212 0 0.00063204 0 0.00063214 3.3 0.00063206 3.3 0.00063216 0 0.00063208 0 0.00063218 3.3 0.0006321 3.3 0.0006322 0 0.00063212 0 0.00063222 3.3 0.00063214 3.3 0.00063224 0 0.00063216 0 0.0006322599999999999 3.3 0.0006321800000000001 3.3 0.00063228 0 0.0006322000000000001 0 0.0006323 3.3 0.0006322200000000001 3.3 0.00063232 0 0.0006322400000000001 0 0.00063234 3.3 0.00063226 3.3 0.00063236 0 0.00063228 0 0.00063238 3.3 0.0006323 3.3 0.0006324 0 0.00063232 0 0.00063242 3.3 0.00063234 3.3 0.00063244 0 0.00063236 0 0.0006324599999999999 3.3 0.00063238 3.3 0.0006324799999999999 0 0.0006324000000000001 0 0.0006325 3.3 0.0006324200000000001 3.3 0.00063252 0 0.0006324400000000001 0 0.00063254 3.3 0.00063246 3.3 0.00063256 0 0.00063248 0 0.00063258 3.3 0.0006325 3.3 0.0006326 0 0.00063252 0 0.00063262 3.3 0.00063254 3.3 0.00063264 0 0.00063256 0 0.00063266 3.3 0.00063258 3.3 0.0006326799999999999 0 0.0006326000000000001 0 0.0006327 3.3 0.0006326200000000001 3.3 0.00063272 0 0.0006326400000000001 0 0.00063274 3.3 0.0006326600000000001 3.3 0.00063276 0 0.00063268 0 0.00063278 3.3 0.0006327 3.3 0.0006328 0 0.00063272 0 0.00063282 3.3 0.00063274 3.3 0.00063284 0 0.00063276 0 0.00063286 3.3 0.00063278 3.3 0.0006328799999999999 0 0.0006328 0 0.0006328999999999999 3.3 0.0006328200000000001 3.3 0.00063292 0 0.0006328400000000001 0 0.00063294 3.3 0.0006328600000000001 3.3 0.00063296 0 0.00063288 0 0.00063298 3.3 0.0006329 3.3 0.000633 0 0.00063292 0 0.00063302 3.3 0.00063294 3.3 0.00063304 0 0.00063296 0 0.00063306 3.3 0.00063298 3.3 0.00063308 0 0.000633 0 0.0006330999999999999 3.3 0.0006330200000000001 3.3 0.00063312 0 0.0006330400000000001 0 0.00063314 3.3 0.0006330600000000001 3.3 0.00063316 0 0.0006330800000000001 0 0.00063318 3.3 0.0006331 3.3 0.0006332 0 0.00063312 0 0.00063322 3.3 0.00063314 3.3 0.00063324 0 0.00063316 0 0.00063326 3.3 0.00063318 3.3 0.00063328 0 0.0006332 0 0.0006332999999999999 3.3 0.00063322 3.3 0.0006333199999999999 0 0.0006332400000000001 0 0.00063334 3.3 0.0006332600000000001 3.3 0.00063336 0 0.0006332800000000001 0 0.00063338 3.3 0.0006333 3.3 0.0006334 0 0.00063332 0 0.00063342 3.3 0.00063334 3.3 0.00063344 0 0.00063336 0 0.00063346 3.3 0.00063338 3.3 0.00063348 0 0.0006334 0 0.0006335 3.3 0.00063342 3.3 0.0006335199999999999 0 0.0006334400000000001 0 0.00063354 3.3 0.0006334600000000001 3.3 0.00063356 0 0.0006334800000000001 0 0.00063358 3.3 0.0006335000000000001 3.3 0.0006336 0 0.00063352 0 0.00063362 3.3 0.00063354 3.3 0.00063364 0 0.00063356 0 0.00063366 3.3 0.00063358 3.3 0.00063368 0 0.0006336 0 0.0006337 3.3 0.00063362 3.3 0.0006337199999999999 0 0.0006336400000000001 0 0.00063374 3.3 0.0006336600000000001 3.3 0.00063376 0 0.0006336800000000001 0 0.00063378 3.3 0.0006337000000000001 3.3 0.0006338 0 0.00063372 0 0.00063382 3.3 0.00063374 3.3 0.00063384 0 0.00063376 0 0.00063386 3.3 0.00063378 3.3 0.00063388 0 0.0006338 0 0.0006339 3.3 0.00063382 3.3 0.00063392 0 0.00063384 0 0.0006339399999999999 3.3 0.0006338600000000001 3.3 0.00063396 0 0.0006338800000000001 0 0.00063398 3.3 0.0006339000000000001 3.3 0.000634 0 0.0006339200000000001 0 0.00063402 3.3 0.00063394 3.3 0.00063404 0 0.00063396 0 0.00063406 3.3 0.00063398 3.3 0.00063408 0 0.000634 0 0.0006341 3.3 0.00063402 3.3 0.00063412 0 0.00063404 0 0.0006341399999999999 3.3 0.0006340600000000001 3.3 0.00063416 0 0.0006340800000000001 0 0.00063418 3.3 0.0006341000000000001 3.3 0.0006342 0 0.0006341200000000001 0 0.00063422 3.3 0.00063414 3.3 0.00063424 0 0.00063416 0 0.00063426 3.3 0.00063418 3.3 0.00063428 0 0.0006342 0 0.0006343 3.3 0.00063422 3.3 0.00063432 0 0.00063424 0 0.00063434 3.3 0.00063426 3.3 0.0006343599999999999 0 0.0006342800000000001 0 0.00063438 3.3 0.0006343000000000001 3.3 0.0006344 0 0.0006343200000000001 0 0.00063442 3.3 0.0006343400000000001 3.3 0.00063444 0 0.00063436 0 0.00063446 3.3 0.00063438 3.3 0.00063448 0 0.0006344 0 0.0006345 3.3 0.00063442 3.3 0.00063452 0 0.00063444 0 0.00063454 3.3 0.00063446 3.3 0.0006345599999999999 0 0.0006344800000000001 0 0.00063458 3.3 0.0006345000000000001 3.3 0.0006346 0 0.0006345200000000001 0 0.00063462 3.3 0.0006345400000000001 3.3 0.00063464 0 0.00063456 0 0.00063466 3.3 0.00063458 3.3 0.00063468 0 0.0006346 0 0.0006347 3.3 0.00063462 3.3 0.00063472 0 0.00063464 0 0.00063474 3.3 0.00063466 3.3 0.00063476 0 0.00063468 0 0.0006347799999999999 3.3 0.0006347000000000001 3.3 0.0006348 0 0.0006347200000000001 0 0.00063482 3.3 0.0006347400000000001 3.3 0.00063484 0 0.0006347600000000001 0 0.00063486 3.3 0.00063478 3.3 0.00063488 0 0.0006348 0 0.0006349 3.3 0.00063482 3.3 0.00063492 0 0.00063484 0 0.00063494 3.3 0.00063486 3.3 0.00063496 0 0.00063488 0 0.0006349799999999999 3.3 0.0006349000000000001 3.3 0.000635 0 0.0006349200000000001 0 0.00063502 3.3 0.0006349400000000001 3.3 0.00063504 0 0.0006349600000000001 0 0.00063506 3.3 0.00063498 3.3 0.00063508 0 0.000635 0 0.0006351 3.3 0.00063502 3.3 0.00063512 0 0.00063504 0 0.00063514 3.3 0.00063506 3.3 0.00063516 0 0.00063508 0 0.00063518 3.3 0.0006351 3.3 0.0006351999999999999 0 0.0006351200000000001 0 0.00063522 3.3 0.0006351400000000001 3.3 0.00063524 0 0.0006351600000000001 0 0.00063526 3.3 0.0006351800000000001 3.3 0.00063528 0 0.0006352 0 0.0006353 3.3 0.00063522 3.3 0.00063532 0 0.00063524 0 0.00063534 3.3 0.00063526 3.3 0.00063536 0 0.00063528 0 0.00063538 3.3 0.0006353 3.3 0.0006353999999999999 0 0.0006353200000000001 0 0.00063542 3.3 0.0006353400000000001 3.3 0.00063544 0 0.0006353600000000001 0 0.00063546 3.3 0.0006353800000000001 3.3 0.00063548 0 0.0006354 0 0.0006355 3.3 0.00063542 3.3 0.00063552 0 0.00063544 0 0.00063554 3.3 0.00063546 3.3 0.00063556 0 0.00063548 0 0.00063558 3.3 0.0006355 3.3 0.0006355999999999999 0 0.00063552 0 0.0006356199999999999 3.3 0.0006355400000000001 3.3 0.00063564 0 0.0006355600000000001 0 0.00063566 3.3 0.0006355800000000001 3.3 0.00063568 0 0.0006356 0 0.0006357 3.3 0.00063562 3.3 0.00063572 0 0.00063564 0 0.00063574 3.3 0.00063566 3.3 0.00063576 0 0.00063568 0 0.00063578 3.3 0.0006357 3.3 0.0006358 0 0.00063572 0 0.0006358199999999999 3.3 0.0006357400000000001 3.3 0.00063584 0 0.0006357600000000001 0 0.00063586 3.3 0.0006357800000000001 3.3 0.00063588 0 0.0006358000000000001 0 0.0006359 3.3 0.00063582 3.3 0.00063592 0 0.00063584 0 0.00063594 3.3 0.00063586 3.3 0.00063596 0 0.00063588 0 0.00063598 3.3 0.0006359 3.3 0.000636 0 0.00063592 0 0.0006360199999999999 3.3 0.00063594 3.3 0.0006360399999999999 0 0.0006359600000000001 0 0.00063606 3.3 0.0006359800000000001 3.3 0.00063608 0 0.0006360000000000001 0 0.0006361 3.3 0.00063602 3.3 0.00063612 0 0.00063604 0 0.00063614 3.3 0.00063606 3.3 0.00063616 0 0.00063608 0 0.00063618 3.3 0.0006361 3.3 0.0006362 0 0.00063612 0 0.00063622 3.3 0.00063614 3.3 0.0006362399999999999 0 0.0006361600000000001 0 0.00063626 3.3 0.0006361800000000001 3.3 0.00063628 0 0.0006362000000000001 0 0.0006363 3.3 0.0006362200000000001 3.3 0.00063632 0 0.00063624 0 0.00063634 3.3 0.00063626 3.3 0.00063636 0 0.00063628 0 0.00063638 3.3 0.0006363 3.3 0.0006364 0 0.00063632 0 0.00063642 3.3 0.00063634 3.3 0.0006364399999999999 0 0.00063636 0 0.0006364599999999999 3.3 0.0006363800000000001 3.3 0.00063648 0 0.0006364000000000001 0 0.0006365 3.3 0.0006364200000000001 3.3 0.00063652 0 0.00063644 0 0.00063654 3.3 0.00063646 3.3 0.00063656 0 0.00063648 0 0.00063658 3.3 0.0006365 3.3 0.0006366 0 0.00063652 0 0.00063662 3.3 0.00063654 3.3 0.00063664 0 0.00063656 0 0.0006366599999999999 3.3 0.0006365800000000001 3.3 0.00063668 0 0.0006366000000000001 0 0.0006367 3.3 0.0006366200000000001 3.3 0.00063672 0 0.0006366400000000001 0 0.00063674 3.3 0.00063666 3.3 0.00063676 0 0.00063668 0 0.00063678 3.3 0.0006367 3.3 0.0006368 0 0.00063672 0 0.00063682 3.3 0.00063674 3.3 0.00063684 0 0.00063676 0 0.0006368599999999999 3.3 0.00063678 3.3 0.0006368799999999999 0 0.0006368000000000001 0 0.0006369 3.3 0.0006368200000000001 3.3 0.00063692 0 0.0006368400000000001 0 0.00063694 3.3 0.00063686 3.3 0.00063696 0 0.00063688 0 0.00063698 3.3 0.0006369 3.3 0.000637 0 0.00063692 0 0.00063702 3.3 0.00063694 3.3 0.00063704 0 0.00063696 0 0.00063706 3.3 0.00063698 3.3 0.0006370799999999999 0 0.0006370000000000001 0 0.0006371 3.3 0.0006370200000000001 3.3 0.00063712 0 0.0006370400000000001 0 0.00063714 3.3 0.0006370600000000001 3.3 0.00063716 0 0.00063708 0 0.00063718 3.3 0.0006371 3.3 0.0006372 0 0.00063712 0 0.00063722 3.3 0.00063714 3.3 0.00063724 0 0.00063716 0 0.00063726 3.3 0.00063718 3.3 0.0006372799999999999 0 0.0006372000000000001 0 0.0006373 3.3 0.0006372200000000001 3.3 0.00063732 0 0.0006372400000000001 0 0.00063734 3.3 0.0006372600000000001 3.3 0.00063736 0 0.00063728 0 0.00063738 3.3 0.0006373 3.3 0.0006374 0 0.00063732 0 0.00063742 3.3 0.00063734 3.3 0.00063744 0 0.00063736 0 0.00063746 3.3 0.00063738 3.3 0.00063748 0 0.0006374 0 0.0006374999999999999 3.3 0.0006374200000000001 3.3 0.00063752 0 0.0006374400000000001 0 0.00063754 3.3 0.0006374600000000001 3.3 0.00063756 0 0.0006374800000000001 0 0.00063758 3.3 0.0006375 3.3 0.0006376 0 0.00063752 0 0.00063762 3.3 0.00063754 3.3 0.00063764 0 0.00063756 0 0.00063766 3.3 0.00063758 3.3 0.00063768 0 0.0006376 0 0.0006376999999999999 3.3 0.0006376200000000001 3.3 0.00063772 0 0.0006376400000000001 0 0.00063774 3.3 0.0006376600000000001 3.3 0.00063776 0 0.0006376800000000001 0 0.00063778 3.3 0.0006377 3.3 0.0006378 0 0.00063772 0 0.00063782 3.3 0.00063774 3.3 0.00063784 0 0.00063776 0 0.00063786 3.3 0.00063778 3.3 0.00063788 0 0.0006378 0 0.0006379 3.3 0.00063782 3.3 0.0006379199999999999 0 0.0006378400000000001 0 0.00063794 3.3 0.0006378600000000001 3.3 0.00063796 0 0.0006378800000000001 0 0.00063798 3.3 0.0006379000000000001 3.3 0.000638 0 0.00063792 0 0.00063802 3.3 0.00063794 3.3 0.00063804 0 0.00063796 0 0.00063806 3.3 0.00063798 3.3 0.00063808 0 0.000638 0 0.0006381 3.3 0.00063802 3.3 0.0006381199999999999 0 0.0006380400000000001 0 0.00063814 3.3 0.0006380600000000001 3.3 0.00063816 0 0.0006380800000000001 0 0.00063818 3.3 0.0006381000000000001 3.3 0.0006382 0 0.00063812 0 0.00063822 3.3 0.00063814 3.3 0.00063824 0 0.00063816 0 0.00063826 3.3 0.00063818 3.3 0.00063828 0 0.0006382 0 0.0006383 3.3 0.00063822 3.3 0.00063832 0 0.00063824 0 0.0006383399999999999 3.3 0.0006382600000000001 3.3 0.00063836 0 0.0006382800000000001 0 0.00063838 3.3 0.0006383000000000001 3.3 0.0006384 0 0.0006383200000000001 0 0.00063842 3.3 0.00063834 3.3 0.00063844 0 0.00063836 0 0.00063846 3.3 0.00063838 3.3 0.00063848 0 0.0006384 0 0.0006385 3.3 0.00063842 3.3 0.00063852 0 0.00063844 0 0.0006385399999999999 3.3 0.0006384600000000001 3.3 0.00063856 0 0.0006384800000000001 0 0.00063858 3.3 0.0006385000000000001 3.3 0.0006386 0 0.0006385200000000001 0 0.00063862 3.3 0.00063854 3.3 0.00063864 0 0.00063856 0 0.00063866 3.3 0.00063858 3.3 0.00063868 0 0.0006386 0 0.0006387 3.3 0.00063862 3.3 0.00063872 0 0.00063864 0 0.00063874 3.3 0.00063866 3.3 0.0006387599999999999 0 0.0006386800000000001 0 0.00063878 3.3 0.0006387000000000001 3.3 0.0006388 0 0.0006387200000000001 0 0.00063882 3.3 0.0006387400000000001 3.3 0.00063884 0 0.00063876 0 0.00063886 3.3 0.00063878 3.3 0.00063888 0 0.0006388 0 0.0006389 3.3 0.00063882 3.3 0.00063892 0 0.00063884 0 0.00063894 3.3 0.00063886 3.3 0.0006389599999999999 0 0.0006388800000000001 0 0.00063898 3.3 0.0006389000000000001 3.3 0.000639 0 0.0006389200000000001 0 0.00063902 3.3 0.0006389400000000001 3.3 0.00063904 0 0.00063896 0 0.00063906 3.3 0.00063898 3.3 0.00063908 0 0.000639 0 0.0006391 3.3 0.00063902 3.3 0.00063912 0 0.00063904 0 0.00063914 3.3 0.00063906 3.3 0.0006391599999999999 0 0.00063908 0 0.0006391799999999999 3.3 0.0006391000000000001 3.3 0.0006392 0 0.0006391200000000001 0 0.00063922 3.3 0.0006391400000000001 3.3 0.00063924 0 0.00063916 0 0.00063926 3.3 0.00063918 3.3 0.00063928 0 0.0006392 0 0.0006393 3.3 0.00063922 3.3 0.00063932 0 0.00063924 0 0.00063934 3.3 0.00063926 3.3 0.00063936 0 0.00063928 0 0.0006393799999999999 3.3 0.0006393000000000001 3.3 0.0006394 0 0.0006393200000000001 0 0.00063942 3.3 0.0006393400000000001 3.3 0.00063944 0 0.0006393600000000001 0 0.00063946 3.3 0.00063938 3.3 0.00063948 0 0.0006394 0 0.0006395 3.3 0.00063942 3.3 0.00063952 0 0.00063944 0 0.00063954 3.3 0.00063946 3.3 0.00063956 0 0.00063948 0 0.0006395799999999999 3.3 0.0006395 3.3 0.0006395999999999999 0 0.0006395200000000001 0 0.00063962 3.3 0.0006395400000000001 3.3 0.00063964 0 0.0006395600000000001 0 0.00063966 3.3 0.00063958 3.3 0.00063968 0 0.0006396 0 0.0006397 3.3 0.00063962 3.3 0.00063972 0 0.00063964 0 0.00063974 3.3 0.00063966 3.3 0.00063976 0 0.00063968 0 0.00063978 3.3 0.0006397 3.3 0.0006397999999999999 0 0.0006397200000000001 0 0.00063982 3.3 0.0006397400000000001 3.3 0.00063984 0 0.0006397600000000001 0 0.00063986 3.3 0.0006397800000000001 3.3 0.00063988 0 0.0006398 0 0.0006399 3.3 0.00063982 3.3 0.00063992 0 0.00063984 0 0.00063994 3.3 0.00063986 3.3 0.00063996 0 0.00063988 0 0.00063998 3.3 0.0006399 3.3 0.0006399999999999999 0 0.00063992 0 0.0006400199999999999 3.3 0.0006399400000000001 3.3 0.00064004 0 0.0006399600000000001 0 0.00064006 3.3 0.0006399800000000001 3.3 0.00064008 0 0.00064 0 0.0006401 3.3 0.00064002 3.3 0.00064012 0 0.00064004 0 0.00064014 3.3 0.00064006 3.3 0.00064016 0 0.00064008 0 0.00064018 3.3 0.0006401 3.3 0.0006402 0 0.00064012 0 0.0006402199999999999 3.3 0.0006401400000000001 3.3 0.00064024 0 0.0006401600000000001 0 0.00064026 3.3 0.0006401800000000001 3.3 0.00064028 0 0.0006402000000000001 0 0.0006403 3.3 0.00064022 3.3 0.00064032 0 0.00064024 0 0.00064034 3.3 0.00064026 3.3 0.00064036 0 0.00064028 0 0.00064038 3.3 0.0006403 3.3 0.0006404 0 0.00064032 0 0.0006404199999999999 3.3 0.00064034 3.3 0.0006404399999999999 0 0.0006403600000000001 0 0.00064046 3.3 0.0006403800000000001 3.3 0.00064048 0 0.0006404000000000001 0 0.0006405 3.3 0.00064042 3.3 0.00064052 0 0.00064044 0 0.00064054 3.3 0.00064046 3.3 0.00064056 0 0.00064048 0 0.00064058 3.3 0.0006405 3.3 0.0006406 0 0.00064052 0 0.00064062 3.3 0.00064054 3.3 0.0006406399999999999 0 0.0006405600000000001 0 0.00064066 3.3 0.0006405800000000001 3.3 0.00064068 0 0.0006406000000000001 0 0.0006407 3.3 0.0006406200000000001 3.3 0.00064072 0 0.00064064 0 0.00064074 3.3 0.00064066 3.3 0.00064076 0 0.00064068 0 0.00064078 3.3 0.0006407 3.3 0.0006408 0 0.00064072 0 0.00064082 3.3 0.00064074 3.3 0.0006408399999999999 0 0.0006407600000000001 0 0.00064086 3.3 0.0006407800000000001 3.3 0.00064088 0 0.0006408000000000001 0 0.0006409 3.3 0.0006408200000000001 3.3 0.00064092 0 0.00064084 0 0.00064094 3.3 0.00064086 3.3 0.00064096 0 0.00064088 0 0.00064098 3.3 0.0006409 3.3 0.000641 0 0.00064092 0 0.00064102 3.3 0.00064094 3.3 0.00064104 0 0.00064096 0 0.0006410599999999999 3.3 0.0006409800000000001 3.3 0.00064108 0 0.0006410000000000001 0 0.0006411 3.3 0.0006410200000000001 3.3 0.00064112 0 0.0006410400000000001 0 0.00064114 3.3 0.00064106 3.3 0.00064116 0 0.00064108 0 0.00064118 3.3 0.0006411 3.3 0.0006412 0 0.00064112 0 0.00064122 3.3 0.00064114 3.3 0.00064124 0 0.00064116 0 0.0006412599999999999 3.3 0.0006411800000000001 3.3 0.00064128 0 0.0006412000000000001 0 0.0006413 3.3 0.0006412200000000001 3.3 0.00064132 0 0.0006412400000000001 0 0.00064134 3.3 0.00064126 3.3 0.00064136 0 0.00064128 0 0.00064138 3.3 0.0006413 3.3 0.0006414 0 0.00064132 0 0.00064142 3.3 0.00064134 3.3 0.00064144 0 0.00064136 0 0.00064146 3.3 0.00064138 3.3 0.0006414799999999999 0 0.0006414000000000001 0 0.0006415 3.3 0.0006414200000000001 3.3 0.00064152 0 0.0006414400000000001 0 0.00064154 3.3 0.0006414600000000001 3.3 0.00064156 0 0.00064148 0 0.00064158 3.3 0.0006415 3.3 0.0006416 0 0.00064152 0 0.00064162 3.3 0.00064154 3.3 0.00064164 0 0.00064156 0 0.00064166 3.3 0.00064158 3.3 0.0006416799999999999 0 0.0006416000000000001 0 0.0006417 3.3 0.0006416200000000001 3.3 0.00064172 0 0.0006416400000000001 0 0.00064174 3.3 0.0006416600000000001 3.3 0.00064176 0 0.00064168 0 0.00064178 3.3 0.0006417 3.3 0.0006418 0 0.00064172 0 0.00064182 3.3 0.00064174 3.3 0.00064184 0 0.00064176 0 0.00064186 3.3 0.00064178 3.3 0.00064188 0 0.0006418 0 0.0006418999999999999 3.3 0.0006418200000000001 3.3 0.00064192 0 0.0006418400000000001 0 0.00064194 3.3 0.0006418600000000001 3.3 0.00064196 0 0.0006418800000000001 0 0.00064198 3.3 0.0006419 3.3 0.000642 0 0.00064192 0 0.00064202 3.3 0.00064194 3.3 0.00064204 0 0.00064196 0 0.00064206 3.3 0.00064198 3.3 0.00064208 0 0.000642 0 0.0006420999999999999 3.3 0.0006420200000000001 3.3 0.00064212 0 0.0006420400000000001 0 0.00064214 3.3 0.0006420600000000001 3.3 0.00064216 0 0.0006420800000000001 0 0.00064218 3.3 0.0006421 3.3 0.0006422 0 0.00064212 0 0.00064222 3.3 0.00064214 3.3 0.00064224 0 0.00064216 0 0.00064226 3.3 0.00064218 3.3 0.00064228 0 0.0006422 0 0.0006422999999999999 3.3 0.00064222 3.3 0.0006423199999999999 0 0.0006422400000000001 0 0.00064234 3.3 0.0006422600000000001 3.3 0.00064236 0 0.0006422800000000001 0 0.00064238 3.3 0.0006423 3.3 0.0006424 0 0.00064232 0 0.00064242 3.3 0.00064234 3.3 0.00064244 0 0.00064236 0 0.00064246 3.3 0.00064238 3.3 0.00064248 0 0.0006424 0 0.0006425 3.3 0.00064242 3.3 0.0006425199999999999 0 0.0006424400000000001 0 0.00064254 3.3 0.0006424600000000001 3.3 0.00064256 0 0.0006424800000000001 0 0.00064258 3.3 0.0006425000000000001 3.3 0.0006426 0 0.00064252 0 0.00064262 3.3 0.00064254 3.3 0.00064264 0 0.00064256 0 0.00064266 3.3 0.00064258 3.3 0.00064268 0 0.0006426 0 0.0006427 3.3 0.00064262 3.3 0.0006427199999999999 0 0.00064264 0 0.0006427399999999999 3.3 0.0006426600000000001 3.3 0.00064276 0 0.0006426800000000001 0 0.00064278 3.3 0.0006427000000000001 3.3 0.0006428 0 0.00064272 0 0.00064282 3.3 0.00064274 3.3 0.00064284 0 0.00064276 0 0.00064286 3.3 0.00064278 3.3 0.00064288 0 0.0006428 0 0.0006429 3.3 0.00064282 3.3 0.00064292 0 0.00064284 0 0.0006429399999999999 3.3 0.0006428600000000001 3.3 0.00064296 0 0.0006428800000000001 0 0.00064298 3.3 0.0006429000000000001 3.3 0.000643 0 0.0006429200000000001 0 0.00064302 3.3 0.00064294 3.3 0.00064304 0 0.00064296 0 0.00064306 3.3 0.00064298 3.3 0.00064308 0 0.000643 0 0.0006431 3.3 0.00064302 3.3 0.00064312 0 0.00064304 0 0.0006431399999999999 3.3 0.00064306 3.3 0.0006431599999999999 0 0.0006430800000000001 0 0.00064318 3.3 0.0006431000000000001 3.3 0.0006432 0 0.0006431200000000001 0 0.00064322 3.3 0.00064314 3.3 0.00064324 0 0.00064316 0 0.00064326 3.3 0.00064318 3.3 0.00064328 0 0.0006432 0 0.0006433 3.3 0.00064322 3.3 0.00064332 0 0.00064324 0 0.00064334 3.3 0.00064326 3.3 0.0006433599999999999 0 0.0006432800000000001 0 0.00064338 3.3 0.0006433000000000001 3.3 0.0006434 0 0.0006433200000000001 0 0.00064342 3.3 0.0006433400000000001 3.3 0.00064344 0 0.00064336 0 0.00064346 3.3 0.00064338 3.3 0.00064348 0 0.0006434 0 0.0006435 3.3 0.00064342 3.3 0.00064352 0 0.00064344 0 0.00064354 3.3 0.00064346 3.3 0.0006435599999999999 0 0.00064348 0 0.0006435799999999999 3.3 0.0006435000000000001 3.3 0.0006436 0 0.0006435200000000001 0 0.00064362 3.3 0.0006435400000000001 3.3 0.00064364 0 0.00064356 0 0.00064366 3.3 0.00064358 3.3 0.00064368 0 0.0006436 0 0.0006437 3.3 0.00064362 3.3 0.00064372 0 0.00064364 0 0.00064374 3.3 0.00064366 3.3 0.00064376 0 0.00064368 0 0.0006437799999999999 3.3 0.0006437000000000001 3.3 0.0006438 0 0.0006437200000000001 0 0.00064382 3.3 0.0006437400000000001 3.3 0.00064384 0 0.0006437600000000001 0 0.00064386 3.3 0.00064378 3.3 0.00064388 0 0.0006438 0 0.0006439 3.3 0.00064382 3.3 0.00064392 0 0.00064384 0 0.00064394 3.3 0.00064386 3.3 0.00064396 0 0.00064388 0 0.0006439799999999999 3.3 0.0006439000000000001 3.3 0.000644 0 0.0006439200000000001 0 0.00064402 3.3 0.0006439400000000001 3.3 0.00064404 0 0.0006439600000000001 0 0.00064406 3.3 0.00064398 3.3 0.00064408 0 0.000644 0 0.0006441 3.3 0.00064402 3.3 0.00064412 0 0.00064404 0 0.00064414 3.3 0.00064406 3.3 0.00064416 0 0.00064408 0 0.00064418 3.3 0.0006441 3.3 0.0006441999999999999 0 0.0006441200000000001 0 0.00064422 3.3 0.0006441400000000001 3.3 0.00064424 0 0.0006441600000000001 0 0.00064426 3.3 0.0006441800000000001 3.3 0.00064428 0 0.0006442 0 0.0006443 3.3 0.00064422 3.3 0.00064432 0 0.00064424 0 0.00064434 3.3 0.00064426 3.3 0.00064436 0 0.00064428 0 0.00064438 3.3 0.0006443 3.3 0.0006443999999999999 0 0.0006443200000000001 0 0.00064442 3.3 0.0006443400000000001 3.3 0.00064444 0 0.0006443600000000001 0 0.00064446 3.3 0.0006443800000000001 3.3 0.00064448 0 0.0006444 0 0.0006445 3.3 0.00064442 3.3 0.00064452 0 0.00064444 0 0.00064454 3.3 0.00064446 3.3 0.00064456 0 0.00064448 0 0.00064458 3.3 0.0006445 3.3 0.0006446 0 0.00064452 0 0.0006446199999999999 3.3 0.0006445400000000001 3.3 0.00064464 0 0.0006445600000000001 0 0.00064466 3.3 0.0006445800000000001 3.3 0.00064468 0 0.0006446000000000001 0 0.0006447 3.3 0.00064462 3.3 0.00064472 0 0.00064464 0 0.00064474 3.3 0.00064466 3.3 0.00064476 0 0.00064468 0 0.00064478 3.3 0.0006447 3.3 0.0006448 0 0.00064472 0 0.0006448199999999999 3.3 0.0006447400000000001 3.3 0.00064484 0 0.0006447600000000001 0 0.00064486 3.3 0.0006447800000000001 3.3 0.00064488 0 0.0006448000000000001 0 0.0006449 3.3 0.00064482 3.3 0.00064492 0 0.00064484 0 0.00064494 3.3 0.00064486 3.3 0.00064496 0 0.00064488 0 0.00064498 3.3 0.0006449 3.3 0.000645 0 0.00064492 0 0.00064502 3.3 0.00064494 3.3 0.0006450399999999999 0 0.0006449600000000001 0 0.00064506 3.3 0.0006449800000000001 3.3 0.00064508 0 0.0006450000000000001 0 0.0006451 3.3 0.0006450200000000001 3.3 0.00064512 0 0.00064504 0 0.00064514 3.3 0.00064506 3.3 0.00064516 0 0.00064508 0 0.00064518 3.3 0.0006451 3.3 0.0006452 0 0.00064512 0 0.00064522 3.3 0.00064514 3.3 0.0006452399999999999 0 0.0006451600000000001 0 0.00064526 3.3 0.0006451800000000001 3.3 0.00064528 0 0.0006452000000000001 0 0.0006453 3.3 0.0006452200000000001 3.3 0.00064532 0 0.00064524 0 0.00064534 3.3 0.00064526 3.3 0.00064536 0 0.00064528 0 0.00064538 3.3 0.0006453 3.3 0.0006454 0 0.00064532 0 0.00064542 3.3 0.00064534 3.3 0.00064544 0 0.00064536 0 0.0006454599999999999 3.3 0.0006453800000000001 3.3 0.00064548 0 0.0006454000000000001 0 0.0006455 3.3 0.0006454200000000001 3.3 0.00064552 0 0.0006454400000000001 0 0.00064554 3.3 0.00064546 3.3 0.00064556 0 0.00064548 0 0.00064558 3.3 0.0006455 3.3 0.0006456 0 0.00064552 0 0.00064562 3.3 0.00064554 3.3 0.00064564 0 0.00064556 0 0.0006456599999999999 3.3 0.0006455800000000001 3.3 0.00064568 0 0.0006456000000000001 0 0.0006457 3.3 0.0006456200000000001 3.3 0.00064572 0 0.0006456400000000001 0 0.00064574 3.3 0.00064566 3.3 0.00064576 0 0.00064568 0 0.00064578 3.3 0.0006457 3.3 0.0006458 0 0.00064572 0 0.00064582 3.3 0.00064574 3.3 0.00064584 0 0.00064576 0 0.0006458599999999999 3.3 0.00064578 3.3 0.0006458799999999999 0 0.0006458000000000001 0 0.0006459 3.3 0.0006458200000000001 3.3 0.00064592 0 0.0006458400000000001 0 0.00064594 3.3 0.00064586 3.3 0.00064596 0 0.00064588 0 0.00064598 3.3 0.0006459 3.3 0.000646 0 0.00064592 0 0.00064602 3.3 0.00064594 3.3 0.00064604 0 0.00064596 0 0.00064606 3.3 0.00064598 3.3 0.0006460799999999999 0 0.0006460000000000001 0 0.0006461 3.3 0.0006460200000000001 3.3 0.00064612 0 0.0006460400000000001 0 0.00064614 3.3 0.0006460600000000001 3.3 0.00064616 0 0.00064608 0 0.00064618 3.3 0.0006461 3.3 0.0006462 0 0.00064612 0 0.00064622 3.3 0.00064614 3.3 0.00064624 0 0.00064616 0 0.00064626 3.3 0.00064618 3.3 0.0006462799999999999 0 0.0006462 0 0.0006462999999999999 3.3 0.0006462200000000001 3.3 0.00064632 0 0.0006462400000000001 0 0.00064634 3.3 0.0006462600000000001 3.3 0.00064636 0 0.00064628 0 0.00064638 3.3 0.0006463 3.3 0.0006464 0 0.00064632 0 0.00064642 3.3 0.00064634 3.3 0.00064644 0 0.00064636 0 0.00064646 3.3 0.00064638 3.3 0.00064648 0 0.0006464 0 0.0006464999999999999 3.3 0.0006464200000000001 3.3 0.00064652 0 0.0006464400000000001 0 0.00064654 3.3 0.0006464600000000001 3.3 0.00064656 0 0.0006464800000000001 0 0.00064658 3.3 0.0006465 3.3 0.0006466 0 0.00064652 0 0.00064662 3.3 0.00064654 3.3 0.00064664 0 0.00064656 0 0.00064666 3.3 0.00064658 3.3 0.00064668 0 0.0006466 0 0.0006466999999999999 3.3 0.00064662 3.3 0.0006467199999999999 0 0.0006466400000000001 0 0.00064674 3.3 0.0006466600000000001 3.3 0.00064676 0 0.0006466800000000001 0 0.00064678 3.3 0.0006467 3.3 0.0006468 0 0.00064672 0 0.00064682 3.3 0.00064674 3.3 0.00064684 0 0.00064676 0 0.00064686 3.3 0.00064678 3.3 0.00064688 0 0.0006468 0 0.0006469 3.3 0.00064682 3.3 0.0006469199999999999 0 0.0006468400000000001 0 0.00064694 3.3 0.0006468600000000001 3.3 0.00064696 0 0.0006468800000000001 0 0.00064698 3.3 0.0006469000000000001 3.3 0.000647 0 0.00064692 0 0.00064702 3.3 0.00064694 3.3 0.00064704 0 0.00064696 0 0.00064706 3.3 0.00064698 3.3 0.00064708 0 0.000647 0 0.0006471 3.3 0.00064702 3.3 0.0006471199999999999 0 0.00064704 0 0.0006471399999999999 3.3 0.0006470600000000001 3.3 0.00064716 0 0.0006470800000000001 0 0.00064718 3.3 0.0006471000000000001 3.3 0.0006472 0 0.00064712 0 0.00064722 3.3 0.00064714 3.3 0.00064724 0 0.00064716 0 0.00064726 3.3 0.00064718 3.3 0.00064728 0 0.0006472 0 0.0006473 3.3 0.00064722 3.3 0.00064732 0 0.00064724 0 0.0006473399999999999 3.3 0.0006472600000000001 3.3 0.00064736 0 0.0006472800000000001 0 0.00064738 3.3 0.0006473000000000001 3.3 0.0006474 0 0.0006473200000000001 0 0.00064742 3.3 0.00064734 3.3 0.00064744 0 0.00064736 0 0.00064746 3.3 0.00064738 3.3 0.00064748 0 0.0006474 0 0.0006475 3.3 0.00064742 3.3 0.00064752 0 0.00064744 0 0.0006475399999999999 3.3 0.0006474600000000001 3.3 0.00064756 0 0.0006474800000000001 0 0.00064758 3.3 0.0006475000000000001 3.3 0.0006476 0 0.0006475200000000001 0 0.00064762 3.3 0.00064754 3.3 0.00064764 0 0.00064756 0 0.00064766 3.3 0.00064758 3.3 0.00064768 0 0.0006476 0 0.0006477 3.3 0.00064762 3.3 0.00064772 0 0.00064764 0 0.00064774 3.3 0.00064766 3.3 0.0006477599999999999 0 0.0006476800000000001 0 0.00064778 3.3 0.0006477000000000001 3.3 0.0006478 0 0.0006477200000000001 0 0.00064782 3.3 0.0006477400000000001 3.3 0.00064784 0 0.00064776 0 0.00064786 3.3 0.00064778 3.3 0.00064788 0 0.0006478 0 0.0006479 3.3 0.00064782 3.3 0.00064792 0 0.00064784 0 0.00064794 3.3 0.00064786 3.3 0.0006479599999999999 0 0.0006478800000000001 0 0.00064798 3.3 0.0006479000000000001 3.3 0.000648 0 0.0006479200000000001 0 0.00064802 3.3 0.0006479400000000001 3.3 0.00064804 0 0.00064796 0 0.00064806 3.3 0.00064798 3.3 0.00064808 0 0.000648 0 0.0006481 3.3 0.00064802 3.3 0.00064812 0 0.00064804 0 0.00064814 3.3 0.00064806 3.3 0.00064816 0 0.00064808 0 0.0006481799999999999 3.3 0.0006481000000000001 3.3 0.0006482 0 0.0006481200000000001 0 0.00064822 3.3 0.0006481400000000001 3.3 0.00064824 0 0.0006481600000000001 0 0.00064826 3.3 0.00064818 3.3 0.00064828 0 0.0006482 0 0.0006483 3.3 0.00064822 3.3 0.00064832 0 0.00064824 0 0.00064834 3.3 0.00064826 3.3 0.00064836 0 0.00064828 0 0.0006483799999999999 3.3 0.0006483000000000001 3.3 0.0006484 0 0.0006483200000000001 0 0.00064842 3.3 0.0006483400000000001 3.3 0.00064844 0 0.0006483600000000001 0 0.00064846 3.3 0.00064838 3.3 0.00064848 0 0.0006484 0 0.0006485 3.3 0.00064842 3.3 0.00064852 0 0.00064844 0 0.00064854 3.3 0.00064846 3.3 0.00064856 0 0.00064848 0 0.00064858 3.3 0.0006485 3.3 0.0006485999999999999 0 0.0006485200000000001 0 0.00064862 3.3 0.0006485400000000001 3.3 0.00064864 0 0.0006485600000000001 0 0.00064866 3.3 0.0006485800000000001 3.3 0.00064868 0 0.0006486 0 0.0006487 3.3 0.00064862 3.3 0.00064872 0 0.00064864 0 0.00064874 3.3 0.00064866 3.3 0.00064876 0 0.00064868 0 0.00064878 3.3 0.0006487 3.3 0.0006487999999999999 0 0.0006487200000000001 0 0.00064882 3.3 0.0006487400000000001 3.3 0.00064884 0 0.0006487600000000001 0 0.00064886 3.3 0.0006487800000000001 3.3 0.00064888 0 0.0006488 0 0.0006489 3.3 0.00064882 3.3 0.00064892 0 0.00064884 0 0.00064894 3.3 0.00064886 3.3 0.00064896 0 0.00064888 0 0.00064898 3.3 0.0006489 3.3 0.000649 0 0.00064892 0 0.0006490199999999999 3.3 0.0006489400000000001 3.3 0.00064904 0 0.0006489600000000001 0 0.00064906 3.3 0.0006489800000000001 3.3 0.00064908 0 0.0006490000000000001 0 0.0006491 3.3 0.00064902 3.3 0.00064912 0 0.00064904 0 0.00064914 3.3 0.00064906 3.3 0.00064916 0 0.00064908 0 0.00064918 3.3 0.0006491 3.3 0.0006492 0 0.00064912 0 0.0006492199999999999 3.3 0.0006491400000000001 3.3 0.00064924 0 0.0006491600000000001 0 0.00064926 3.3 0.0006491800000000001 3.3 0.00064928 0 0.0006492000000000001 0 0.0006493 3.3 0.00064922 3.3 0.00064932 0 0.00064924 0 0.00064934 3.3 0.00064926 3.3 0.00064936 0 0.00064928 0 0.00064938 3.3 0.0006493 3.3 0.0006494 0 0.00064932 0 0.0006494199999999999 3.3 0.00064934 3.3 0.0006494399999999999 0 0.0006493600000000001 0 0.00064946 3.3 0.0006493800000000001 3.3 0.00064948 0 0.0006494000000000001 0 0.0006495 3.3 0.00064942 3.3 0.00064952 0 0.00064944 0 0.00064954 3.3 0.00064946 3.3 0.00064956 0 0.00064948 0 0.00064958 3.3 0.0006495 3.3 0.0006496 0 0.00064952 0 0.00064962 3.3 0.00064954 3.3 0.0006496399999999999 0 0.0006495600000000001 0 0.00064966 3.3 0.0006495800000000001 3.3 0.00064968 0 0.0006496000000000001 0 0.0006497 3.3 0.0006496200000000001 3.3 0.00064972 0 0.00064964 0 0.00064974 3.3 0.00064966 3.3 0.00064976 0 0.00064968 0 0.00064978 3.3 0.0006497 3.3 0.0006498 0 0.00064972 0 0.00064982 3.3 0.00064974 3.3 0.0006498399999999999 0 0.00064976 0 0.0006498599999999999 3.3 0.0006497800000000001 3.3 0.00064988 0 0.0006498000000000001 0 0.0006499 3.3 0.0006498200000000001 3.3 0.00064992 0 0.00064984 0 0.00064994 3.3 0.00064986 3.3 0.00064996 0 0.00064988 0 0.00064998 3.3 0.0006499 3.3 0.00065 0 0.00064992 0 0.00065002 3.3 0.00064994 3.3 0.00065004 0 0.00064996 0 0.0006500599999999999 3.3 0.0006499800000000001 3.3 0.00065008 0 0.0006500000000000001 0 0.0006501 3.3 0.0006500200000000001 3.3 0.00065012 0 0.0006500400000000001 0 0.00065014 3.3 0.00065006 3.3 0.00065016 0 0.00065008 0 0.00065018 3.3 0.0006501 3.3 0.0006502 0 0.00065012 0 0.00065022 3.3 0.00065014 3.3 0.00065024 0 0.00065016 0 0.0006502599999999999 3.3 0.00065018 3.3 0.0006502799999999999 0 0.0006502000000000001 0 0.0006503 3.3 0.0006502200000000001 3.3 0.00065032 0 0.0006502400000000001 0 0.00065034 3.3 0.00065026 3.3 0.00065036 0 0.00065028 0 0.00065038 3.3 0.0006503 3.3 0.0006504 0 0.00065032 0 0.00065042 3.3 0.00065034 3.3 0.00065044 0 0.00065036 0 0.00065046 3.3 0.00065038 3.3 0.0006504799999999999 0 0.0006504000000000001 0 0.0006505 3.3 0.0006504200000000001 3.3 0.00065052 0 0.0006504400000000001 0 0.00065054 3.3 0.0006504600000000001 3.3 0.00065056 0 0.00065048 0 0.00065058 3.3 0.0006505 3.3 0.0006506 0 0.00065052 0 0.00065062 3.3 0.00065054 3.3 0.00065064 0 0.00065056 0 0.00065066 3.3 0.00065058 3.3 0.0006506799999999999 0 0.0006506 0 0.0006506999999999999 3.3 0.0006506200000000001 3.3 0.00065072 0 0.0006506400000000001 0 0.00065074 3.3 0.0006506600000000001 3.3 0.00065076 0 0.00065068 0 0.00065078 3.3 0.0006507 3.3 0.0006508 0 0.00065072 0 0.00065082 3.3 0.00065074 3.3 0.00065084 0 0.00065076 0 0.00065086 3.3 0.00065078 3.3 0.00065088 0 0.0006508 0 0.0006508999999999999 3.3 0.0006508200000000001 3.3 0.00065092 0 0.0006508400000000001 0 0.00065094 3.3 0.0006508600000000001 3.3 0.00065096 0 0.0006508800000000001 0 0.00065098 3.3 0.0006509 3.3 0.000651 0 0.00065092 0 0.00065102 3.3 0.00065094 3.3 0.00065104 0 0.00065096 0 0.00065106 3.3 0.00065098 3.3 0.00065108 0 0.000651 0 0.0006510999999999999 3.3 0.0006510200000000001 3.3 0.00065112 0 0.0006510400000000001 0 0.00065114 3.3 0.0006510600000000001 3.3 0.00065116 0 0.0006510800000000001 0 0.00065118 3.3 0.0006511 3.3 0.0006512 0 0.00065112 0 0.00065122 3.3 0.00065114 3.3 0.00065124 0 0.00065116 0 0.00065126 3.3 0.00065118 3.3 0.00065128 0 0.0006512 0 0.0006513 3.3 0.00065122 3.3 0.0006513199999999999 0 0.0006512400000000001 0 0.00065134 3.3 0.0006512600000000001 3.3 0.00065136 0 0.0006512800000000001 0 0.00065138 3.3 0.0006513000000000001 3.3 0.0006514 0 0.00065132 0 0.00065142 3.3 0.00065134 3.3 0.00065144 0 0.00065136 0 0.00065146 3.3 0.00065138 3.3 0.00065148 0 0.0006514 0 0.0006515 3.3 0.00065142 3.3 0.0006515199999999999 0 0.0006514400000000001 0 0.00065154 3.3 0.0006514600000000001 3.3 0.00065156 0 0.0006514800000000001 0 0.00065158 3.3 0.0006515000000000001 3.3 0.0006516 0 0.00065152 0 0.00065162 3.3 0.00065154 3.3 0.00065164 0 0.00065156 0 0.00065166 3.3 0.00065158 3.3 0.00065168 0 0.0006516 0 0.0006517 3.3 0.00065162 3.3 0.00065172 0 0.00065164 0 0.0006517399999999999 3.3 0.0006516600000000001 3.3 0.00065176 0 0.0006516800000000001 0 0.00065178 3.3 0.0006517000000000001 3.3 0.0006518 0 0.0006517200000000001 0 0.00065182 3.3 0.00065174 3.3 0.00065184 0 0.00065176 0 0.00065186 3.3 0.00065178 3.3 0.00065188 0 0.0006518 0 0.0006519 3.3 0.00065182 3.3 0.00065192 0 0.00065184 0 0.0006519399999999999 3.3 0.0006518600000000001 3.3 0.00065196 0 0.0006518800000000001 0 0.00065198 3.3 0.0006519000000000001 3.3 0.000652 0 0.0006519200000000001 0 0.00065202 3.3 0.00065194 3.3 0.00065204 0 0.00065196 0 0.00065206 3.3 0.00065198 3.3 0.00065208 0 0.000652 0 0.0006521 3.3 0.00065202 3.3 0.00065212 0 0.00065204 0 0.00065214 3.3 0.00065206 3.3 0.0006521599999999999 0 0.0006520800000000001 0 0.00065218 3.3 0.0006521000000000001 3.3 0.0006522 0 0.0006521200000000001 0 0.00065222 3.3 0.0006521400000000001 3.3 0.00065224 0 0.00065216 0 0.00065226 3.3 0.00065218 3.3 0.00065228 0 0.0006522 0 0.0006523 3.3 0.00065222 3.3 0.00065232 0 0.00065224 0 0.00065234 3.3 0.00065226 3.3 0.0006523599999999999 0 0.0006522800000000001 0 0.00065238 3.3 0.0006523000000000001 3.3 0.0006524 0 0.0006523200000000001 0 0.00065242 3.3 0.0006523400000000001 3.3 0.00065244 0 0.00065236 0 0.00065246 3.3 0.00065238 3.3 0.00065248 0 0.0006524 0 0.0006525 3.3 0.00065242 3.3 0.00065252 0 0.00065244 0 0.00065254 3.3 0.00065246 3.3 0.0006525599999999999 0 0.00065248 0 0.0006525799999999999 3.3 0.0006525000000000001 3.3 0.0006526 0 0.0006525200000000001 0 0.00065262 3.3 0.0006525400000000001 3.3 0.00065264 0 0.00065256 0 0.00065266 3.3 0.00065258 3.3 0.00065268 0 0.0006526 0 0.0006527 3.3 0.00065262 3.3 0.00065272 0 0.00065264 0 0.00065274 3.3 0.00065266 3.3 0.00065276 0 0.00065268 0 0.0006527799999999999 3.3 0.0006527000000000001 3.3 0.0006528 0 0.0006527200000000001 0 0.00065282 3.3 0.0006527400000000001 3.3 0.00065284 0 0.0006527600000000001 0 0.00065286 3.3 0.00065278 3.3 0.00065288 0 0.0006528 0 0.0006529 3.3 0.00065282 3.3 0.00065292 0 0.00065284 0 0.00065294 3.3 0.00065286 3.3 0.00065296 0 0.00065288 0 0.0006529799999999999 3.3 0.0006529 3.3 0.0006529999999999999 0 0.0006529200000000001 0 0.00065302 3.3 0.0006529400000000001 3.3 0.00065304 0 0.0006529600000000001 0 0.00065306 3.3 0.00065298 3.3 0.00065308 0 0.000653 0 0.0006531 3.3 0.00065302 3.3 0.00065312 0 0.00065304 0 0.00065314 3.3 0.00065306 3.3 0.00065316 0 0.00065308 0 0.00065318 3.3 0.0006531 3.3 0.0006531999999999999 0 0.0006531200000000001 0 0.00065322 3.3 0.0006531400000000001 3.3 0.00065324 0 0.0006531600000000001 0 0.00065326 3.3 0.0006531800000000001 3.3 0.00065328 0 0.0006532 0 0.0006533 3.3 0.00065322 3.3 0.00065332 0 0.00065324 0 0.00065334 3.3 0.00065326 3.3 0.00065336 0 0.00065328 0 0.00065338 3.3 0.0006533 3.3 0.0006533999999999999 0 0.00065332 0 0.0006534199999999999 3.3 0.0006533400000000001 3.3 0.00065344 0 0.0006533600000000001 0 0.00065346 3.3 0.0006533800000000001 3.3 0.00065348 0 0.0006534 0 0.0006535 3.3 0.00065342 3.3 0.00065352 0 0.00065344 0 0.00065354 3.3 0.00065346 3.3 0.00065356 0 0.00065348 0 0.00065358 3.3 0.0006535 3.3 0.0006536 0 0.00065352 0 0.0006536199999999999 3.3 0.0006535400000000001 3.3 0.00065364 0 0.0006535600000000001 0 0.00065366 3.3 0.0006535800000000001 3.3 0.00065368 0 0.0006536000000000001 0 0.0006537 3.3 0.00065362 3.3 0.00065372 0 0.00065364 0 0.00065374 3.3 0.00065366 3.3 0.00065376 0 0.00065368 0 0.00065378 3.3 0.0006537 3.3 0.0006538 0 0.00065372 0 0.0006538199999999999 3.3 0.00065374 3.3 0.0006538399999999999 0 0.0006537600000000001 0 0.00065386 3.3 0.0006537800000000001 3.3 0.00065388 0 0.0006538000000000001 0 0.0006539 3.3 0.00065382 3.3 0.00065392 0 0.00065384 0 0.00065394 3.3 0.00065386 3.3 0.00065396 0 0.00065388 0 0.00065398 3.3 0.0006539 3.3 0.000654 0 0.00065392 0 0.00065402 3.3 0.00065394 3.3 0.0006540399999999999 0 0.0006539600000000001 0 0.00065406 3.3 0.0006539800000000001 3.3 0.00065408 0 0.0006540000000000001 0 0.0006541 3.3 0.0006540200000000001 3.3 0.00065412 0 0.00065404 0 0.00065414 3.3 0.00065406 3.3 0.00065416 0 0.00065408 0 0.00065418 3.3 0.0006541 3.3 0.0006542 0 0.00065412 0 0.00065422 3.3 0.00065414 3.3 0.0006542399999999999 0 0.00065416 0 0.0006542599999999999 3.3 0.0006541800000000001 3.3 0.00065428 0 0.0006542000000000001 0 0.0006543 3.3 0.0006542200000000001 3.3 0.00065432 0 0.00065424 0 0.00065434 3.3 0.00065426 3.3 0.00065436 0 0.00065428 0 0.00065438 3.3 0.0006543 3.3 0.0006544 0 0.00065432 0 0.00065442 3.3 0.00065434 3.3 0.00065444 0 0.00065436 0 0.0006544599999999999 3.3 0.0006543800000000001 3.3 0.00065448 0 0.0006544000000000001 0 0.0006545 3.3 0.0006544200000000001 3.3 0.00065452 0 0.0006544400000000001 0 0.00065454 3.3 0.00065446 3.3 0.00065456 0 0.00065448 0 0.00065458 3.3 0.0006545 3.3 0.0006546 0 0.00065452 0 0.00065462 3.3 0.00065454 3.3 0.00065464 0 0.00065456 0 0.0006546599999999999 3.3 0.0006545800000000001 3.3 0.00065468 0 0.0006546000000000001 0 0.0006547 3.3 0.0006546200000000001 3.3 0.00065472 0 0.0006546400000000001 0 0.00065474 3.3 0.00065466 3.3 0.00065476 0 0.00065468 0 0.00065478 3.3 0.0006547 3.3 0.0006548 0 0.00065472 0 0.00065482 3.3 0.00065474 3.3 0.00065484 0 0.00065476 0 0.00065486 3.3 0.00065478 3.3 0.0006548799999999999 0 0.0006548000000000001 0 0.0006549 3.3 0.0006548200000000001 3.3 0.00065492 0 0.0006548400000000001 0 0.00065494 3.3 0.0006548600000000001 3.3 0.00065496 0 0.00065488 0 0.00065498 3.3 0.0006549 3.3 0.000655 0 0.00065492 0 0.00065502 3.3 0.00065494 3.3 0.00065504 0 0.00065496 0 0.00065506 3.3 0.00065498 3.3 0.0006550799999999999 0 0.0006550000000000001 0 0.0006551 3.3 0.0006550200000000001 3.3 0.00065512 0 0.0006550400000000001 0 0.00065514 3.3 0.0006550600000000001 3.3 0.00065516 0 0.00065508 0 0.00065518 3.3 0.0006551 3.3 0.0006552 0 0.00065512 0 0.00065522 3.3 0.00065514 3.3 0.00065524 0 0.00065516 0 0.00065526 3.3 0.00065518 3.3 0.00065528 0 0.0006552 0 0.0006552999999999999 3.3 0.0006552200000000001 3.3 0.00065532 0 0.0006552400000000001 0 0.00065534 3.3 0.0006552600000000001 3.3 0.00065536 0 0.0006552800000000001 0 0.00065538 3.3 0.0006553 3.3 0.0006554 0 0.00065532 0 0.00065542 3.3 0.00065534 3.3 0.00065544 0 0.00065536 0 0.00065546 3.3 0.00065538 3.3 0.00065548 0 0.0006554 0 0.0006554999999999999 3.3 0.0006554200000000001 3.3 0.00065552 0 0.0006554400000000001 0 0.00065554 3.3 0.0006554600000000001 3.3 0.00065556 0 0.0006554800000000001 0 0.00065558 3.3 0.0006555 3.3 0.0006556 0 0.00065552 0 0.00065562 3.3 0.00065554 3.3 0.00065564 0 0.00065556 0 0.00065566 3.3 0.00065558 3.3 0.00065568 0 0.0006556 0 0.0006557 3.3 0.00065562 3.3 0.0006557199999999999 0 0.0006556400000000001 0 0.00065574 3.3 0.0006556600000000001 3.3 0.00065576 0 0.0006556800000000001 0 0.00065578 3.3 0.0006557000000000001 3.3 0.0006558 0 0.00065572 0 0.00065582 3.3 0.00065574 3.3 0.00065584 0 0.00065576 0 0.00065586 3.3 0.00065578 3.3 0.00065588 0 0.0006558 0 0.0006559 3.3 0.00065582 3.3 0.0006559199999999999 0 0.0006558400000000001 0 0.00065594 3.3 0.0006558600000000001 3.3 0.00065596 0 0.0006558800000000001 0 0.00065598 3.3 0.0006559000000000001 3.3 0.000656 0 0.00065592 0 0.00065602 3.3 0.00065594 3.3 0.00065604 0 0.00065596 0 0.00065606 3.3 0.00065598 3.3 0.00065608 0 0.000656 0 0.0006561 3.3 0.00065602 3.3 0.0006561199999999999 0 0.00065604 0 0.0006561399999999999 3.3 0.0006560600000000001 3.3 0.00065616 0 0.0006560800000000001 0 0.00065618 3.3 0.0006561000000000001 3.3 0.0006562 0 0.00065612 0 0.00065622 3.3 0.00065614 3.3 0.00065624 0 0.00065616 0 0.00065626 3.3 0.00065618 3.3 0.00065628 0 0.0006562 0 0.0006563 3.3 0.00065622 3.3 0.00065632 0 0.00065624 0 0.0006563399999999999 3.3 0.0006562600000000001 3.3 0.00065636 0 0.0006562800000000001 0 0.00065638 3.3 0.0006563000000000001 3.3 0.0006564 0 0.0006563200000000001 0 0.00065642 3.3 0.00065634 3.3 0.00065644 0 0.00065636 0 0.00065646 3.3 0.00065638 3.3 0.00065648 0 0.0006564 0 0.0006565 3.3 0.00065642 3.3 0.00065652 0 0.00065644 0 0.0006565399999999999 3.3 0.00065646 3.3 0.0006565599999999999 0 0.0006564800000000001 0 0.00065658 3.3 0.0006565000000000001 3.3 0.0006566 0 0.0006565200000000001 0 0.00065662 3.3 0.00065654 3.3 0.00065664 0 0.00065656 0 0.00065666 3.3 0.00065658 3.3 0.00065668 0 0.0006566 0 0.0006567 3.3 0.00065662 3.3 0.00065672 0 0.00065664 0 0.00065674 3.3 0.00065666 3.3 0.0006567599999999999 0 0.0006566800000000001 0 0.00065678 3.3 0.0006567000000000001 3.3 0.0006568 0 0.0006567200000000001 0 0.00065682 3.3 0.0006567400000000001 3.3 0.00065684 0 0.00065676 0 0.00065686 3.3 0.00065678 3.3 0.00065688 0 0.0006568 0 0.0006569 3.3 0.00065682 3.3 0.00065692 0 0.00065684 0 0.00065694 3.3 0.00065686 3.3 0.0006569599999999999 0 0.00065688 0 0.0006569799999999999 3.3 0.0006569000000000001 3.3 0.000657 0 0.0006569200000000001 0 0.00065702 3.3 0.0006569400000000001 3.3 0.00065704 0 0.00065696 0 0.00065706 3.3 0.00065698 3.3 0.00065708 0 0.000657 0 0.0006571 3.3 0.00065702 3.3 0.00065712 0 0.00065704 0 0.00065714 3.3 0.00065706 3.3 0.00065716 0 0.00065708 0 0.0006571799999999999 3.3 0.0006571000000000001 3.3 0.0006572 0 0.0006571200000000001 0 0.00065722 3.3 0.0006571400000000001 3.3 0.00065724 0 0.0006571600000000001 0 0.00065726 3.3 0.00065718 3.3 0.00065728 0 0.0006572 0 0.0006573 3.3 0.00065722 3.3 0.00065732 0 0.00065724 0 0.00065734 3.3 0.00065726 3.3 0.00065736 0 0.00065728 0 0.0006573799999999999 3.3 0.0006573 3.3 0.0006573999999999999 0 0.0006573200000000001 0 0.00065742 3.3 0.0006573400000000001 3.3 0.00065744 0 0.0006573600000000001 0 0.00065746 3.3 0.00065738 3.3 0.00065748 0 0.0006574 0 0.0006575 3.3 0.00065742 3.3 0.00065752 0 0.00065744 0 0.00065754 3.3 0.00065746 3.3 0.00065756 0 0.00065748 0 0.00065758 3.3 0.0006575 3.3 0.0006575999999999999 0 0.0006575200000000001 0 0.00065762 3.3 0.0006575400000000001 3.3 0.00065764 0 0.0006575600000000001 0 0.00065766 3.3 0.0006575800000000001 3.3 0.00065768 0 0.0006576 0 0.0006577 3.3 0.00065762 3.3 0.00065772 0 0.00065764 0 0.00065774 3.3 0.00065766 3.3 0.00065776 0 0.00065768 0 0.00065778 3.3 0.0006577 3.3 0.0006577999999999999 0 0.00065772 0 0.0006578199999999999 3.3 0.0006577400000000001 3.3 0.00065784 0 0.0006577600000000001 0 0.00065786 3.3 0.0006577800000000001 3.3 0.00065788 0 0.0006578 0 0.0006579 3.3 0.00065782 3.3 0.00065792 0 0.00065784 0 0.00065794 3.3 0.00065786 3.3 0.00065796 0 0.00065788 0 0.00065798 3.3 0.0006579 3.3 0.000658 0 0.00065792 0 0.0006580199999999999 3.3 0.0006579400000000001 3.3 0.00065804 0 0.0006579600000000001 0 0.00065806 3.3 0.0006579800000000001 3.3 0.00065808 0 0.0006580000000000001 0 0.0006581 3.3 0.00065802 3.3 0.00065812 0 0.00065804 0 0.00065814 3.3 0.00065806 3.3 0.00065816 0 0.00065808 0 0.00065818 3.3 0.0006581 3.3 0.0006582 0 0.00065812 0 0.0006582199999999999 3.3 0.0006581400000000001 3.3 0.00065824 0 0.0006581600000000001 0 0.00065826 3.3 0.0006581800000000001 3.3 0.00065828 0 0.0006582000000000001 0 0.0006583 3.3 0.00065822 3.3 0.00065832 0 0.00065824 0 0.00065834 3.3 0.00065826 3.3 0.00065836 0 0.00065828 0 0.00065838 3.3 0.0006583 3.3 0.0006584 0 0.00065832 0 0.00065842 3.3 0.00065834 3.3 0.0006584399999999999 0 0.0006583600000000001 0 0.00065846 3.3 0.0006583800000000001 3.3 0.00065848 0 0.0006584000000000001 0 0.0006585 3.3 0.0006584200000000001 3.3 0.00065852 0 0.00065844 0 0.00065854 3.3 0.00065846 3.3 0.00065856 0 0.00065848 0 0.00065858 3.3 0.0006585 3.3 0.0006586 0 0.00065852 0 0.00065862 3.3 0.00065854 3.3 0.0006586399999999999 0 0.0006585600000000001 0 0.00065866 3.3 0.0006585800000000001 3.3 0.00065868 0 0.0006586000000000001 0 0.0006587 3.3 0.0006586200000000001 3.3 0.00065872 0 0.00065864 0 0.00065874 3.3 0.00065866 3.3 0.00065876 0 0.00065868 0 0.00065878 3.3 0.0006587 3.3 0.0006588 0 0.00065872 0 0.00065882 3.3 0.00065874 3.3 0.00065884 0 0.00065876 0 0.0006588599999999999 3.3 0.0006587800000000001 3.3 0.00065888 0 0.0006588000000000001 0 0.0006589 3.3 0.0006588200000000001 3.3 0.00065892 0 0.0006588400000000001 0 0.00065894 3.3 0.00065886 3.3 0.00065896 0 0.00065888 0 0.00065898 3.3 0.0006589 3.3 0.000659 0 0.00065892 0 0.00065902 3.3 0.00065894 3.3 0.00065904 0 0.00065896 0 0.0006590599999999999 3.3 0.0006589800000000001 3.3 0.00065908 0 0.0006590000000000001 0 0.0006591 3.3 0.0006590200000000001 3.3 0.00065912 0 0.0006590400000000001 0 0.00065914 3.3 0.00065906 3.3 0.00065916 0 0.00065908 0 0.00065918 3.3 0.0006591 3.3 0.0006592 0 0.00065912 0 0.00065922 3.3 0.00065914 3.3 0.00065924 0 0.00065916 0 0.00065926 3.3 0.00065918 3.3 0.0006592799999999999 0 0.0006592000000000001 0 0.0006593 3.3 0.0006592200000000001 3.3 0.00065932 0 0.0006592400000000001 0 0.00065934 3.3 0.0006592600000000001 3.3 0.00065936 0 0.00065928 0 0.00065938 3.3 0.0006593 3.3 0.0006594 0 0.00065932 0 0.00065942 3.3 0.00065934 3.3 0.00065944 0 0.00065936 0 0.00065946 3.3 0.00065938 3.3 0.0006594799999999999 0 0.0006594000000000001 0 0.0006595 3.3 0.0006594200000000001 3.3 0.00065952 0 0.0006594400000000001 0 0.00065954 3.3 0.0006594600000000001 3.3 0.00065956 0 0.00065948 0 0.00065958 3.3 0.0006595 3.3 0.0006596 0 0.00065952 0 0.00065962 3.3 0.00065954 3.3 0.00065964 0 0.00065956 0 0.00065966 3.3 0.00065958 3.3 0.0006596799999999999 0 0.0006596 0 0.0006596999999999999 3.3 0.0006596200000000001 3.3 0.00065972 0 0.0006596400000000001 0 0.00065974 3.3 0.0006596600000000001 3.3 0.00065976 0 0.00065968 0 0.00065978 3.3 0.0006597 3.3 0.0006598 0 0.00065972 0 0.00065982 3.3 0.00065974 3.3 0.00065984 0 0.00065976 0 0.00065986 3.3 0.00065978 3.3 0.00065988 0 0.0006598 0 0.0006598999999999999 3.3 0.0006598200000000001 3.3 0.00065992 0 0.0006598400000000001 0 0.00065994 3.3 0.0006598600000000001 3.3 0.00065996 0 0.0006598800000000001 0 0.00065998 3.3 0.0006599 3.3 0.00066 0 0.00065992 0 0.00066002 3.3 0.00065994 3.3 0.00066004 0 0.00065996 0 0.00066006 3.3 0.00065998 3.3 0.00066008 0 0.00066 0 0.0006600999999999999 3.3 0.00066002 3.3 0.0006601199999999999 0 0.0006600400000000001 0 0.00066014 3.3 0.0006600600000000001 3.3 0.00066016 0 0.0006600800000000001 0 0.00066018 3.3 0.0006601 3.3 0.0006602 0 0.00066012 0 0.00066022 3.3 0.00066014 3.3 0.00066024 0 0.00066016 0 0.00066026 3.3 0.00066018 3.3 0.00066028 0 0.0006602 0 0.0006603 3.3 0.00066022 3.3 0.0006603199999999999 0 0.0006602400000000001 0 0.00066034 3.3 0.0006602600000000001 3.3 0.00066036 0 0.0006602800000000001 0 0.00066038 3.3 0.0006603000000000001 3.3 0.0006604 0 0.00066032 0 0.00066042 3.3 0.00066034 3.3 0.00066044 0 0.00066036 0 0.00066046 3.3 0.00066038 3.3 0.00066048 0 0.0006604 0 0.0006605 3.3 0.00066042 3.3 0.0006605199999999999 0 0.00066044 0 0.0006605399999999999 3.3 0.0006604600000000001 3.3 0.00066056 0 0.0006604800000000001 0 0.00066058 3.3 0.0006605000000000001 3.3 0.0006606 0 0.00066052 0 0.00066062 3.3 0.00066054 3.3 0.00066064 0 0.00066056 0 0.00066066 3.3 0.00066058 3.3 0.00066068 0 0.0006606 0 0.0006607 3.3 0.00066062 3.3 0.00066072 0 0.00066064 0 0.0006607399999999999 3.3 0.0006606600000000001 3.3 0.00066076 0 0.0006606800000000001 0 0.00066078 3.3 0.0006607000000000001 3.3 0.0006608 0 0.0006607200000000001 0 0.00066082 3.3 0.00066074 3.3 0.00066084 0 0.00066076 0 0.00066086 3.3 0.00066078 3.3 0.00066088 0 0.0006608 0 0.0006609 3.3 0.00066082 3.3 0.00066092 0 0.00066084 0 0.0006609399999999999 3.3 0.00066086 3.3 0.0006609599999999999 0 0.0006608800000000001 0 0.00066098 3.3 0.0006609000000000001 3.3 0.000661 0 0.0006609200000000001 0 0.00066102 3.3 0.00066094 3.3 0.00066104 0 0.00066096 0 0.00066106 3.3 0.00066098 3.3 0.00066108 0 0.000661 0 0.0006611 3.3 0.00066102 3.3 0.00066112 0 0.00066104 0 0.00066114 3.3 0.00066106 3.3 0.0006611599999999999 0 0.0006610800000000001 0 0.00066118 3.3 0.0006611000000000001 3.3 0.0006612 0 0.0006611200000000001 0 0.00066122 3.3 0.0006611400000000001 3.3 0.00066124 0 0.00066116 0 0.00066126 3.3 0.00066118 3.3 0.00066128 0 0.0006612 0 0.0006613 3.3 0.00066122 3.3 0.00066132 0 0.00066124 0 0.00066134 3.3 0.00066126 3.3 0.0006613599999999999 0 0.0006612800000000001 0 0.00066138 3.3 0.0006613000000000001 3.3 0.0006614 0 0.0006613200000000001 0 0.00066142 3.3 0.0006613400000000001 3.3 0.00066144 0 0.00066136 0 0.00066146 3.3 0.00066138 3.3 0.00066148 0 0.0006614 0 0.0006615 3.3 0.00066142 3.3 0.00066152 0 0.00066144 0 0.00066154 3.3 0.00066146 3.3 0.00066156 0 0.00066148 0 0.0006615799999999999 3.3 0.0006615000000000001 3.3 0.0006616 0 0.0006615200000000001 0 0.00066162 3.3 0.0006615400000000001 3.3 0.00066164 0 0.0006615600000000001 0 0.00066166 3.3 0.00066158 3.3 0.00066168 0 0.0006616 0 0.0006617 3.3 0.00066162 3.3 0.00066172 0 0.00066164 0 0.00066174 3.3 0.00066166 3.3 0.00066176 0 0.00066168 0 0.0006617799999999999 3.3 0.0006617000000000001 3.3 0.0006618 0 0.0006617200000000001 0 0.00066182 3.3 0.0006617400000000001 3.3 0.00066184 0 0.0006617600000000001 0 0.00066186 3.3 0.00066178 3.3 0.00066188 0 0.0006618 0 0.0006619 3.3 0.00066182 3.3 0.00066192 0 0.00066184 0 0.00066194 3.3 0.00066186 3.3 0.00066196 0 0.00066188 0 0.00066198 3.3 0.0006619 3.3 0.0006619999999999999 0 0.0006619200000000001 0 0.00066202 3.3 0.0006619400000000001 3.3 0.00066204 0 0.0006619600000000001 0 0.00066206 3.3 0.0006619800000000001 3.3 0.00066208 0 0.000662 0 0.0006621 3.3 0.00066202 3.3 0.00066212 0 0.00066204 0 0.00066214 3.3 0.00066206 3.3 0.00066216 0 0.00066208 0 0.00066218 3.3 0.0006621 3.3 0.0006621999999999999 0 0.0006621200000000001 0 0.00066222 3.3 0.0006621400000000001 3.3 0.00066224 0 0.0006621600000000001 0 0.00066226 3.3 0.0006621800000000001 3.3 0.00066228 0 0.0006622 0 0.0006623 3.3 0.00066222 3.3 0.00066232 0 0.00066224 0 0.00066234 3.3 0.00066226 3.3 0.00066236 0 0.00066228 0 0.00066238 3.3 0.0006623 3.3 0.0006624 0 0.00066232 0 0.0006624199999999999 3.3 0.0006623400000000001 3.3 0.00066244 0 0.0006623600000000001 0 0.00066246 3.3 0.0006623800000000001 3.3 0.00066248 0 0.0006624000000000001 0 0.0006625 3.3 0.00066242 3.3 0.00066252 0 0.00066244 0 0.00066254 3.3 0.00066246 3.3 0.00066256 0 0.00066248 0 0.00066258 3.3 0.0006625 3.3 0.0006626 0 0.00066252 0 0.0006626199999999999 3.3 0.0006625400000000001 3.3 0.00066264 0 0.0006625600000000001 0 0.00066266 3.3 0.0006625800000000001 3.3 0.00066268 0 0.0006626000000000001 0 0.0006627 3.3 0.00066262 3.3 0.00066272 0 0.00066264 0 0.00066274 3.3 0.00066266 3.3 0.00066276 0 0.00066268 0 0.00066278 3.3 0.0006627 3.3 0.0006628 0 0.00066272 0 0.0006628199999999999 3.3 0.00066274 3.3 0.0006628399999999999 0 0.0006627600000000001 0 0.00066286 3.3 0.0006627800000000001 3.3 0.00066288 0 0.0006628000000000001 0 0.0006629 3.3 0.00066282 3.3 0.00066292 0 0.00066284 0 0.00066294 3.3 0.00066286 3.3 0.00066296 0 0.00066288 0 0.00066298 3.3 0.0006629 3.3 0.000663 0 0.00066292 0 0.00066302 3.3 0.00066294 3.3 0.0006630399999999999 0 0.0006629600000000001 0 0.00066306 3.3 0.0006629800000000001 3.3 0.00066308 0 0.0006630000000000001 0 0.0006631 3.3 0.0006630200000000001 3.3 0.00066312 0 0.00066304 0 0.00066314 3.3 0.00066306 3.3 0.00066316 0 0.00066308 0 0.00066318 3.3 0.0006631 3.3 0.0006632 0 0.00066312 0 0.00066322 3.3 0.00066314 3.3 0.0006632399999999999 0 0.00066316 0 0.0006632599999999999 3.3 0.0006631800000000001 3.3 0.00066328 0 0.0006632000000000001 0 0.0006633 3.3 0.0006632200000000001 3.3 0.00066332 0 0.00066324 0 0.00066334 3.3 0.00066326 3.3 0.00066336 0 0.00066328 0 0.00066338 3.3 0.0006633 3.3 0.0006634 0 0.00066332 0 0.00066342 3.3 0.00066334 3.3 0.00066344 0 0.00066336 0 0.0006634599999999999 3.3 0.0006633800000000001 3.3 0.00066348 0 0.0006634000000000001 0 0.0006635 3.3 0.0006634200000000001 3.3 0.00066352 0 0.0006634400000000001 0 0.00066354 3.3 0.00066346 3.3 0.00066356 0 0.00066348 0 0.00066358 3.3 0.0006635 3.3 0.0006636 0 0.00066352 0 0.00066362 3.3 0.00066354 3.3 0.00066364 0 0.00066356 0 0.0006636599999999999 3.3 0.00066358 3.3 0.0006636799999999999 0 0.0006636000000000001 0 0.0006637 3.3 0.0006636200000000001 3.3 0.00066372 0 0.0006636400000000001 0 0.00066374 3.3 0.00066366 3.3 0.00066376 0 0.00066368 0 0.00066378 3.3 0.0006637 3.3 0.0006638 0 0.00066372 0 0.00066382 3.3 0.00066374 3.3 0.00066384 0 0.00066376 0 0.00066386 3.3 0.00066378 3.3 0.0006638799999999999 0 0.0006638000000000001 0 0.0006639 3.3 0.0006638200000000001 3.3 0.00066392 0 0.0006638400000000001 0 0.00066394 3.3 0.0006638600000000001 3.3 0.00066396 0 0.00066388 0 0.00066398 3.3 0.0006639 3.3 0.000664 0 0.00066392 0 0.00066402 3.3 0.00066394 3.3 0.00066404 0 0.00066396 0 0.00066406 3.3 0.00066398 3.3 0.0006640799999999999 0 0.000664 0 0.0006640999999999999 3.3 0.0006640200000000001 3.3 0.00066412 0 0.0006640400000000001 0 0.00066414 3.3 0.0006640600000000001 3.3 0.00066416 0 0.00066408 0 0.00066418 3.3 0.0006641 3.3 0.0006642 0 0.00066412 0 0.00066422 3.3 0.00066414 3.3 0.00066424 0 0.00066416 0 0.00066426 3.3 0.00066418 3.3 0.00066428 0 0.0006642 0 0.0006642999999999999 3.3 0.0006642200000000001 3.3 0.00066432 0 0.0006642400000000001 0 0.00066434 3.3 0.0006642600000000001 3.3 0.00066436 0 0.0006642800000000001 0 0.00066438 3.3 0.0006643 3.3 0.0006644 0 0.00066432 0 0.00066442 3.3 0.00066434 3.3 0.00066444 0 0.00066436 0 0.00066446 3.3 0.00066438 3.3 0.00066448 0 0.0006644 0 0.0006644999999999999 3.3 0.00066442 3.3 0.0006645199999999999 0 0.0006644400000000001 0 0.00066454 3.3 0.0006644600000000001 3.3 0.00066456 0 0.0006644800000000001 0 0.00066458 3.3 0.0006645 3.3 0.0006646 0 0.00066452 0 0.00066462 3.3 0.00066454 3.3 0.00066464 0 0.00066456 0 0.00066466 3.3 0.00066458 3.3 0.00066468 0 0.0006646 0 0.0006647 3.3 0.00066462 3.3 0.0006647199999999999 0 0.0006646400000000001 0 0.00066474 3.3 0.0006646600000000001 3.3 0.00066476 0 0.0006646800000000001 0 0.00066478 3.3 0.0006647000000000001 3.3 0.0006648 0 0.00066472 0 0.00066482 3.3 0.00066474 3.3 0.00066484 0 0.00066476 0 0.00066486 3.3 0.00066478 3.3 0.00066488 0 0.0006648 0 0.0006649 3.3 0.00066482 3.3 0.0006649199999999999 0 0.0006648400000000001 0 0.00066494 3.3 0.0006648600000000001 3.3 0.00066496 0 0.0006648800000000001 0 0.00066498 3.3 0.0006649000000000001 3.3 0.000665 0 0.00066492 0 0.00066502 3.3 0.00066494 3.3 0.00066504 0 0.00066496 0 0.00066506 3.3 0.00066498 3.3 0.00066508 0 0.000665 0 0.0006651 3.3 0.00066502 3.3 0.00066512 0 0.00066504 0 0.0006651399999999999 3.3 0.0006650600000000001 3.3 0.00066516 0 0.0006650800000000001 0 0.00066518 3.3 0.0006651000000000001 3.3 0.0006652 0 0.0006651200000000001 0 0.00066522 3.3 0.00066514 3.3 0.00066524 0 0.00066516 0 0.00066526 3.3 0.00066518 3.3 0.00066528 0 0.0006652 0 0.0006653 3.3 0.00066522 3.3 0.00066532 0 0.00066524 0 0.0006653399999999999 3.3 0.0006652600000000001 3.3 0.00066536 0 0.0006652800000000001 0 0.00066538 3.3 0.0006653000000000001 3.3 0.0006654 0 0.0006653200000000001 0 0.00066542 3.3 0.00066534 3.3 0.00066544 0 0.00066536 0 0.00066546 3.3 0.00066538 3.3 0.00066548 0 0.0006654 0 0.0006655 3.3 0.00066542 3.3 0.00066552 0 0.00066544 0 0.00066554 3.3 0.00066546 3.3 0.0006655599999999999 0 0.0006654800000000001 0 0.00066558 3.3 0.0006655000000000001 3.3 0.0006656 0 0.0006655200000000001 0 0.00066562 3.3 0.0006655400000000001 3.3 0.00066564 0 0.00066556 0 0.00066566 3.3 0.00066558 3.3 0.00066568 0 0.0006656 0 0.0006657 3.3 0.00066562 3.3 0.00066572 0 0.00066564 0 0.00066574 3.3 0.00066566 3.3 0.0006657599999999999 0 0.0006656800000000001 0 0.00066578 3.3 0.0006657000000000001 3.3 0.0006658 0 0.0006657200000000001 0 0.00066582 3.3 0.0006657400000000001 3.3 0.00066584 0 0.00066576 0 0.00066586 3.3 0.00066578 3.3 0.00066588 0 0.0006658 0 0.0006659 3.3 0.00066582 3.3 0.00066592 0 0.00066584 0 0.00066594 3.3 0.00066586 3.3 0.00066596 0 0.00066588 0 0.0006659799999999999 3.3 0.0006659000000000001 3.3 0.000666 0 0.0006659200000000001 0 0.00066602 3.3 0.0006659400000000001 3.3 0.00066604 0 0.0006659600000000001 0 0.00066606 3.3 0.00066598 3.3 0.00066608 0 0.000666 0 0.0006661 3.3 0.00066602 3.3 0.00066612 0 0.00066604 0 0.00066614 3.3 0.00066606 3.3 0.00066616 0 0.00066608 0 0.0006661799999999999 3.3 0.0006661000000000001 3.3 0.0006662 0 0.0006661200000000001 0 0.00066622 3.3 0.0006661400000000001 3.3 0.00066624 0 0.0006661600000000001 0 0.00066626 3.3 0.00066618 3.3 0.00066628 0 0.0006662 0 0.0006663 3.3 0.00066622 3.3 0.00066632 0 0.00066624 0 0.00066634 3.3 0.00066626 3.3 0.00066636 0 0.00066628 0 0.0006663799999999999 3.3 0.0006663 3.3 0.0006663999999999999 0 0.0006663200000000001 0 0.00066642 3.3 0.0006663400000000001 3.3 0.00066644 0 0.0006663600000000001 0 0.00066646 3.3 0.00066638 3.3 0.00066648 0 0.0006664 0 0.0006665 3.3 0.00066642 3.3 0.00066652 0 0.00066644 0 0.00066654 3.3 0.00066646 3.3 0.00066656 0 0.00066648 0 0.00066658 3.3 0.0006665 3.3 0.0006665999999999999 0 0.0006665200000000001 0 0.00066662 3.3 0.0006665400000000001 3.3 0.00066664 0 0.0006665600000000001 0 0.00066666 3.3 0.0006665800000000001 3.3 0.00066668 0 0.0006666 0 0.0006667 3.3 0.00066662 3.3 0.00066672 0 0.00066664 0 0.00066674 3.3 0.00066666 3.3 0.00066676 0 0.00066668 0 0.00066678 3.3 0.0006667 3.3 0.0006667999999999999 0 0.00066672 0 0.0006668199999999999 3.3 0.0006667400000000001 3.3 0.00066684 0 0.0006667600000000001 0 0.00066686 3.3 0.0006667800000000001 3.3 0.00066688 0 0.0006668 0 0.0006669 3.3 0.00066682 3.3 0.00066692 0 0.00066684 0 0.00066694 3.3 0.00066686 3.3 0.00066696 0 0.00066688 0 0.00066698 3.3 0.0006669 3.3 0.000667 0 0.00066692 0 0.0006670199999999999 3.3 0.0006669400000000001 3.3 0.00066704 0 0.0006669600000000001 0 0.00066706 3.3 0.0006669800000000001 3.3 0.00066708 0 0.0006670000000000001 0 0.0006671 3.3 0.00066702 3.3 0.00066712 0 0.00066704 0 0.00066714 3.3 0.00066706 3.3 0.00066716 0 0.00066708 0 0.00066718 3.3 0.0006671 3.3 0.0006672 0 0.00066712 0 0.0006672199999999999 3.3 0.00066714 3.3 0.0006672399999999999 0 0.0006671600000000001 0 0.00066726 3.3 0.0006671800000000001 3.3 0.00066728 0 0.0006672000000000001 0 0.0006673 3.3 0.00066722 3.3 0.00066732 0 0.00066724 0 0.00066734 3.3 0.00066726 3.3 0.00066736 0 0.00066728 0 0.00066738 3.3 0.0006673 3.3 0.0006674 0 0.00066732 0 0.00066742 3.3 0.00066734 3.3 0.0006674399999999999 0 0.0006673600000000001 0 0.00066746 3.3 0.0006673800000000001 3.3 0.00066748 0 0.0006674000000000001 0 0.0006675 3.3 0.0006674200000000001 3.3 0.00066752 0 0.00066744 0 0.00066754 3.3 0.00066746 3.3 0.00066756 0 0.00066748 0 0.00066758 3.3 0.0006675 3.3 0.0006676 0 0.00066752 0 0.00066762 3.3 0.00066754 3.3 0.0006676399999999999 0 0.00066756 0 0.0006676599999999999 3.3 0.0006675800000000001 3.3 0.00066768 0 0.0006676000000000001 0 0.0006677 3.3 0.0006676200000000001 3.3 0.00066772 0 0.00066764 0 0.00066774 3.3 0.00066766 3.3 0.00066776 0 0.00066768 0 0.00066778 3.3 0.0006677 3.3 0.0006678 0 0.00066772 0 0.00066782 3.3 0.00066774 3.3 0.00066784 0 0.00066776 0 0.0006678599999999999 3.3 0.0006677800000000001 3.3 0.00066788 0 0.0006678000000000001 0 0.0006679 3.3 0.0006678200000000001 3.3 0.00066792 0 0.0006678400000000001 0 0.00066794 3.3 0.00066786 3.3 0.00066796 0 0.00066788 0 0.00066798 3.3 0.0006679 3.3 0.000668 0 0.00066792 0 0.00066802 3.3 0.00066794 3.3 0.00066804 0 0.00066796 0 0.0006680599999999999 3.3 0.00066798 3.3 0.0006680799999999999 0 0.0006680000000000001 0 0.0006681 3.3 0.0006680200000000001 3.3 0.00066812 0 0.0006680400000000001 0 0.00066814 3.3 0.00066806 3.3 0.00066816 0 0.00066808 0 0.00066818 3.3 0.0006681 3.3 0.0006682 0 0.00066812 0 0.00066822 3.3 0.00066814 3.3 0.00066824 0 0.00066816 0 0.00066826 3.3 0.00066818 3.3 0.0006682799999999999 0 0.0006682000000000001 0 0.0006683 3.3 0.0006682200000000001 3.3 0.00066832 0 0.0006682400000000001 0 0.00066834 3.3 0.0006682600000000001 3.3 0.00066836 0 0.00066828 0 0.00066838 3.3 0.0006683 3.3 0.0006684 0 0.00066832 0 0.00066842 3.3 0.00066834 3.3 0.00066844 0 0.00066836 0 0.00066846 3.3 0.00066838 3.3 0.0006684799999999999 0 0.0006684000000000001 0 0.0006685 3.3 0.0006684200000000001 3.3 0.00066852 0 0.0006684400000000001 0 0.00066854 3.3 0.0006684600000000001 3.3 0.00066856 0 0.00066848 0 0.00066858 3.3 0.0006685 3.3 0.0006686 0 0.00066852 0 0.00066862 3.3 0.00066854 3.3 0.00066864 0 0.00066856 0 0.00066866 3.3 0.00066858 3.3 0.00066868 0 0.0006686 0 0.0006686999999999999 3.3 0.0006686200000000001 3.3 0.00066872 0 0.0006686400000000001 0 0.00066874 3.3 0.0006686600000000001 3.3 0.00066876 0 0.0006686800000000001 0 0.00066878 3.3 0.0006687 3.3 0.0006688 0 0.00066872 0 0.00066882 3.3 0.00066874 3.3 0.00066884 0 0.00066876 0 0.00066886 3.3 0.00066878 3.3 0.00066888 0 0.0006688 0 0.0006688999999999999 3.3 0.0006688200000000001 3.3 0.00066892 0 0.0006688400000000001 0 0.00066894 3.3 0.0006688600000000001 3.3 0.00066896 0 0.0006688800000000001 0 0.00066898 3.3 0.0006689 3.3 0.000669 0 0.00066892 0 0.00066902 3.3 0.00066894 3.3 0.00066904 0 0.00066896 0 0.00066906 3.3 0.00066898 3.3 0.00066908 0 0.000669 0 0.0006691 3.3 0.00066902 3.3 0.0006691199999999999 0 0.0006690400000000001 0 0.00066914 3.3 0.0006690600000000001 3.3 0.00066916 0 0.0006690800000000001 0 0.00066918 3.3 0.0006691000000000001 3.3 0.0006692 0 0.00066912 0 0.00066922 3.3 0.00066914 3.3 0.00066924 0 0.00066916 0 0.00066926 3.3 0.00066918 3.3 0.00066928 0 0.0006692 0 0.0006693 3.3 0.00066922 3.3 0.0006693199999999999 0 0.0006692400000000001 0 0.00066934 3.3 0.0006692600000000001 3.3 0.00066936 0 0.0006692800000000001 0 0.00066938 3.3 0.0006693000000000001 3.3 0.0006694 0 0.00066932 0 0.00066942 3.3 0.00066934 3.3 0.00066944 0 0.00066936 0 0.00066946 3.3 0.00066938 3.3 0.00066948 0 0.0006694 0 0.0006695 3.3 0.00066942 3.3 0.00066952 0 0.00066944 0 0.0006695399999999999 3.3 0.0006694600000000001 3.3 0.00066956 0 0.0006694800000000001 0 0.00066958 3.3 0.0006695000000000001 3.3 0.0006696 0 0.0006695200000000001 0 0.00066962 3.3 0.00066954 3.3 0.00066964 0 0.00066956 0 0.00066966 3.3 0.00066958 3.3 0.00066968 0 0.0006696 0 0.0006697 3.3 0.00066962 3.3 0.00066972 0 0.00066964 0 0.0006697399999999999 3.3 0.0006696600000000001 3.3 0.00066976 0 0.0006696800000000001 0 0.00066978 3.3 0.0006697000000000001 3.3 0.0006698 0 0.0006697200000000001 0 0.00066982 3.3 0.00066974 3.3 0.00066984 0 0.00066976 0 0.00066986 3.3 0.00066978 3.3 0.00066988 0 0.0006698 0 0.0006699 3.3 0.00066982 3.3 0.00066992 0 0.00066984 0 0.0006699399999999999 3.3 0.00066986 3.3 0.0006699599999999999 0 0.0006698800000000001 0 0.00066998 3.3 0.0006699000000000001 3.3 0.00067 0 0.0006699200000000001 0 0.00067002 3.3 0.00066994 3.3 0.00067004 0 0.00066996 0 0.00067006 3.3 0.00066998 3.3 0.00067008 0 0.00067 0 0.0006701 3.3 0.00067002 3.3 0.00067012 0 0.00067004 0 0.00067014 3.3 0.00067006 3.3 0.0006701599999999999 0 0.0006700800000000001 0 0.00067018 3.3 0.0006701000000000001 3.3 0.0006702 0 0.0006701200000000001 0 0.00067022 3.3 0.0006701400000000001 3.3 0.00067024 0 0.00067016 0 0.00067026 3.3 0.00067018 3.3 0.00067028 0 0.0006702 0 0.0006703 3.3 0.00067022 3.3 0.00067032 0 0.00067024 0 0.00067034 3.3 0.00067026 3.3 0.0006703599999999999 0 0.00067028 0 0.0006703799999999999 3.3 0.0006703000000000001 3.3 0.0006704 0 0.0006703200000000001 0 0.00067042 3.3 0.0006703400000000001 3.3 0.00067044 0 0.00067036 0 0.00067046 3.3 0.00067038 3.3 0.00067048 0 0.0006704 0 0.0006705 3.3 0.00067042 3.3 0.00067052 0 0.00067044 0 0.00067054 3.3 0.00067046 3.3 0.00067056 0 0.00067048 0 0.0006705799999999999 3.3 0.0006705000000000001 3.3 0.0006706 0 0.0006705200000000001 0 0.00067062 3.3 0.0006705400000000001 3.3 0.00067064 0 0.0006705600000000001 0 0.00067066 3.3 0.00067058 3.3 0.00067068 0 0.0006706 0 0.0006707 3.3 0.00067062 3.3 0.00067072 0 0.00067064 0 0.00067074 3.3 0.00067066 3.3 0.00067076 0 0.00067068 0 0.0006707799999999999 3.3 0.0006707 3.3 0.0006707999999999999 0 0.0006707200000000001 0 0.00067082 3.3 0.0006707400000000001 3.3 0.00067084 0 0.0006707600000000001 0 0.00067086 3.3 0.00067078 3.3 0.00067088 0 0.0006708 0 0.0006709 3.3 0.00067082 3.3 0.00067092 0 0.00067084 0 0.00067094 3.3 0.00067086 3.3 0.00067096 0 0.00067088 0 0.00067098 3.3 0.0006709 3.3 0.0006709999999999999 0 0.0006709200000000001 0 0.00067102 3.3 0.0006709400000000001 3.3 0.00067104 0 0.0006709600000000001 0 0.00067106 3.3 0.0006709800000000001 3.3 0.00067108 0 0.000671 0 0.0006711 3.3 0.00067102 3.3 0.00067112 0 0.00067104 0 0.00067114 3.3 0.00067106 3.3 0.00067116 0 0.00067108 0 0.00067118 3.3 0.0006711 3.3 0.0006711999999999999 0 0.00067112 0 0.0006712199999999999 3.3 0.0006711400000000001 3.3 0.00067124 0 0.0006711600000000001 0 0.00067126 3.3 0.0006711800000000001 3.3 0.00067128 0 0.0006712 0 0.0006713 3.3 0.00067122 3.3 0.00067132 0 0.00067124 0 0.00067134 3.3 0.00067126 3.3 0.00067136 0 0.00067128 0 0.00067138 3.3 0.0006713 3.3 0.0006714 0 0.00067132 0 0.0006714199999999999 3.3 0.0006713400000000001 3.3 0.00067144 0 0.0006713600000000001 0 0.00067146 3.3 0.0006713800000000001 3.3 0.00067148 0 0.0006714000000000001 0 0.0006715 3.3 0.00067142 3.3 0.00067152 0 0.00067144 0 0.00067154 3.3 0.00067146 3.3 0.00067156 0 0.00067148 0 0.00067158 3.3 0.0006715 3.3 0.0006716 0 0.00067152 0 0.0006716199999999999 3.3 0.00067154 3.3 0.0006716399999999999 0 0.0006715600000000001 0 0.00067166 3.3 0.0006715800000000001 3.3 0.00067168 0 0.0006716000000000001 0 0.0006717 3.3 0.00067162 3.3 0.00067172 0 0.00067164 0 0.00067174 3.3 0.00067166 3.3 0.00067176 0 0.00067168 0 0.00067178 3.3 0.0006717 3.3 0.0006718 0 0.00067172 0 0.00067182 3.3 0.00067174 3.3 0.0006718399999999999 0 0.0006717600000000001 0 0.00067186 3.3 0.0006717800000000001 3.3 0.00067188 0 0.0006718000000000001 0 0.0006719 3.3 0.0006718200000000001 3.3 0.00067192 0 0.00067184 0 0.00067194 3.3 0.00067186 3.3 0.00067196 0 0.00067188 0 0.00067198 3.3 0.0006719 3.3 0.000672 0 0.00067192 0 0.00067202 3.3 0.00067194 3.3 0.0006720399999999999 0 0.0006719600000000001 0 0.00067206 3.3 0.0006719800000000001 3.3 0.00067208 0 0.0006720000000000001 0 0.0006721 3.3 0.0006720200000000001 3.3 0.00067212 0 0.00067204 0 0.00067214 3.3 0.00067206 3.3 0.00067216 0 0.00067208 0 0.00067218 3.3 0.0006721 3.3 0.0006722 0 0.00067212 0 0.00067222 3.3 0.00067214 3.3 0.00067224 0 0.00067216 0 0.0006722599999999999 3.3 0.0006721800000000001 3.3 0.00067228 0 0.0006722000000000001 0 0.0006723 3.3 0.0006722200000000001 3.3 0.00067232 0 0.0006722400000000001 0 0.00067234 3.3 0.00067226 3.3 0.00067236 0 0.00067228 0 0.00067238 3.3 0.0006723 3.3 0.0006724 0 0.00067232 0 0.00067242 3.3 0.00067234 3.3 0.00067244 0 0.00067236 0 0.0006724599999999999 3.3 0.0006723800000000001 3.3 0.00067248 0 0.0006724000000000001 0 0.0006725 3.3 0.0006724200000000001 3.3 0.00067252 0 0.0006724400000000001 0 0.00067254 3.3 0.00067246 3.3 0.00067256 0 0.00067248 0 0.00067258 3.3 0.0006725 3.3 0.0006726 0 0.00067252 0 0.00067262 3.3 0.00067254 3.3 0.00067264 0 0.00067256 0 0.00067266 3.3 0.00067258 3.3 0.0006726799999999999 0 0.0006726000000000001 0 0.0006727 3.3 0.0006726200000000001 3.3 0.00067272 0 0.0006726400000000001 0 0.00067274 3.3 0.0006726600000000001 3.3 0.00067276 0 0.00067268 0 0.00067278 3.3 0.0006727 3.3 0.0006728 0 0.00067272 0 0.00067282 3.3 0.00067274 3.3 0.00067284 0 0.00067276 0 0.00067286 3.3 0.00067278 3.3 0.0006728799999999999 0 0.0006728000000000001 0 0.0006729 3.3 0.0006728200000000001 3.3 0.00067292 0 0.0006728400000000001 0 0.00067294 3.3 0.0006728600000000001 3.3 0.00067296 0 0.00067288 0 0.00067298 3.3 0.0006729 3.3 0.000673 0 0.00067292 0 0.00067302 3.3 0.00067294 3.3 0.00067304 0 0.00067296 0 0.00067306 3.3 0.00067298 3.3 0.0006730799999999999 0 0.000673 0 0.0006730999999999999 3.3 0.0006730200000000001 3.3 0.00067312 0 0.0006730400000000001 0 0.00067314 3.3 0.0006730600000000001 3.3 0.00067316 0 0.00067308 0 0.00067318 3.3 0.0006731 3.3 0.0006732 0 0.00067312 0 0.00067322 3.3 0.00067314 3.3 0.00067324 0 0.00067316 0 0.00067326 3.3 0.00067318 3.3 0.00067328 0 0.0006732 0 0.0006732999999999999 3.3 0.0006732200000000001 3.3 0.00067332 0 0.0006732400000000001 0 0.00067334 3.3 0.0006732600000000001 3.3 0.00067336 0 0.0006732800000000001 0 0.00067338 3.3 0.0006733 3.3 0.0006734 0 0.00067332 0 0.00067342 3.3 0.00067334 3.3 0.00067344 0 0.00067336 0 0.00067346 3.3 0.00067338 3.3 0.00067348 0 0.0006734 0 0.0006734999999999999 3.3 0.00067342 3.3 0.0006735199999999999 0 0.0006734400000000001 0 0.00067354 3.3 0.0006734600000000001 3.3 0.00067356 0 0.0006734800000000001 0 0.00067358 3.3 0.0006735 3.3 0.0006736 0 0.00067352 0 0.00067362 3.3 0.00067354 3.3 0.00067364 0 0.00067356 0 0.00067366 3.3 0.00067358 3.3 0.00067368 0 0.0006736 0 0.0006737 3.3 0.00067362 3.3 0.0006737199999999999 0 0.0006736400000000001 0 0.00067374 3.3 0.0006736600000000001 3.3 0.00067376 0 0.0006736800000000001 0 0.00067378 3.3 0.0006737000000000001 3.3 0.0006738 0 0.00067372 0 0.00067382 3.3 0.00067374 3.3 0.00067384 0 0.00067376 0 0.00067386 3.3 0.00067378 3.3 0.00067388 0 0.0006738 0 0.0006739 3.3 0.00067382 3.3 0.0006739199999999999 0 0.00067384 0 0.0006739399999999999 3.3 0.0006738600000000001 3.3 0.00067396 0 0.0006738800000000001 0 0.00067398 3.3 0.0006739000000000001 3.3 0.000674 0 0.00067392 0 0.00067402 3.3 0.00067394 3.3 0.00067404 0 0.00067396 0 0.00067406 3.3 0.00067398 3.3 0.00067408 0 0.000674 0 0.0006741 3.3 0.00067402 3.3 0.00067412 0 0.00067404 0 0.0006741399999999999 3.3 0.0006740600000000001 3.3 0.00067416 0 0.0006740800000000001 0 0.00067418 3.3 0.0006741000000000001 3.3 0.0006742 0 0.0006741200000000001 0 0.00067422 3.3 0.00067414 3.3 0.00067424 0 0.00067416 0 0.00067426 3.3 0.00067418 3.3 0.00067428 0 0.0006742 0 0.0006743 3.3 0.00067422 3.3 0.00067432 0 0.00067424 0 0.0006743399999999999 3.3 0.00067426 3.3 0.0006743599999999999 0 0.0006742800000000001 0 0.00067438 3.3 0.0006743000000000001 3.3 0.0006744 0 0.0006743200000000001 0 0.00067442 3.3 0.00067434 3.3 0.00067444 0 0.00067436 0 0.00067446 3.3 0.00067438 3.3 0.00067448 0 0.0006744 0 0.0006745 3.3 0.00067442 3.3 0.00067452 0 0.00067444 0 0.00067454 3.3 0.00067446 3.3 0.0006745599999999999 0 0.0006744800000000001 0 0.00067458 3.3 0.0006745000000000001 3.3 0.0006746 0 0.0006745200000000001 0 0.00067462 3.3 0.0006745400000000001 3.3 0.00067464 0 0.00067456 0 0.00067466 3.3 0.00067458 3.3 0.00067468 0 0.0006746 0 0.0006747 3.3 0.00067462 3.3 0.00067472 0 0.00067464 0 0.00067474 3.3 0.00067466 3.3 0.0006747599999999999 0 0.00067468 0 0.0006747799999999999 3.3 0.0006747000000000001 3.3 0.0006748 0 0.0006747200000000001 0 0.00067482 3.3 0.0006747400000000001 3.3 0.00067484 0 0.00067476 0 0.00067486 3.3 0.00067478 3.3 0.00067488 0 0.0006748 0 0.0006749 3.3 0.00067482 3.3 0.00067492 0 0.00067484 0 0.00067494 3.3 0.00067486 3.3 0.00067496 0 0.00067488 0 0.0006749799999999999 3.3 0.0006749000000000001 3.3 0.000675 0 0.0006749200000000001 0 0.00067502 3.3 0.0006749400000000001 3.3 0.00067504 0 0.0006749600000000001 0 0.00067506 3.3 0.00067498 3.3 0.00067508 0 0.000675 0 0.0006751 3.3 0.00067502 3.3 0.00067512 0 0.00067504 0 0.00067514 3.3 0.00067506 3.3 0.00067516 0 0.00067508 0 0.0006751799999999999 3.3 0.0006751000000000001 3.3 0.0006752 0 0.0006751200000000001 0 0.00067522 3.3 0.0006751400000000001 3.3 0.00067524 0 0.0006751600000000001 0 0.00067526 3.3 0.00067518 3.3 0.00067528 0 0.0006752 0 0.0006753 3.3 0.00067522 3.3 0.00067532 0 0.00067524 0 0.00067534 3.3 0.00067526 3.3 0.00067536 0 0.00067528 0 0.00067538 3.3 0.0006753 3.3 0.0006753999999999999 0 0.0006753200000000001 0 0.00067542 3.3 0.0006753400000000001 3.3 0.00067544 0 0.0006753600000000001 0 0.00067546 3.3 0.0006753800000000001 3.3 0.00067548 0 0.0006754 0 0.0006755 3.3 0.00067542 3.3 0.00067552 0 0.00067544 0 0.00067554 3.3 0.00067546 3.3 0.00067556 0 0.00067548 0 0.00067558 3.3 0.0006755 3.3 0.0006755999999999999 0 0.0006755200000000001 0 0.00067562 3.3 0.0006755400000000001 3.3 0.00067564 0 0.0006755600000000001 0 0.00067566 3.3 0.0006755800000000001 3.3 0.00067568 0 0.0006756 0 0.0006757 3.3 0.00067562 3.3 0.00067572 0 0.00067564 0 0.00067574 3.3 0.00067566 3.3 0.00067576 0 0.00067568 0 0.00067578 3.3 0.0006757 3.3 0.0006758 0 0.00067572 0 0.0006758199999999999 3.3 0.0006757400000000001 3.3 0.00067584 0 0.0006757600000000001 0 0.00067586 3.3 0.0006757800000000001 3.3 0.00067588 0 0.0006758000000000001 0 0.0006759 3.3 0.00067582 3.3 0.00067592 0 0.00067584 0 0.00067594 3.3 0.00067586 3.3 0.00067596 0 0.00067588 0 0.00067598 3.3 0.0006759 3.3 0.000676 0 0.00067592 0 0.0006760199999999999 3.3 0.0006759400000000001 3.3 0.00067604 0 0.0006759600000000001 0 0.00067606 3.3 0.0006759800000000001 3.3 0.00067608 0 0.0006760000000000001 0 0.0006761 3.3 0.00067602 3.3 0.00067612 0 0.00067604 0 0.00067614 3.3 0.00067606 3.3 0.00067616 0 0.00067608 0 0.00067618 3.3 0.0006761 3.3 0.0006762 0 0.00067612 0 0.00067622 3.3 0.00067614 3.3 0.0006762399999999999 0 0.0006761600000000001 0 0.00067626 3.3 0.0006761800000000001 3.3 0.00067628 0 0.0006762000000000001 0 0.0006763 3.3 0.0006762200000000001 3.3 0.00067632 0 0.00067624 0 0.00067634 3.3 0.00067626 3.3 0.00067636 0 0.00067628 0 0.00067638 3.3 0.0006763 3.3 0.0006764 0 0.00067632 0 0.00067642 3.3 0.00067634 3.3 0.0006764399999999999 0 0.0006763600000000001 0 0.00067646 3.3 0.0006763800000000001 3.3 0.00067648 0 0.0006764000000000001 0 0.0006765 3.3 0.0006764200000000001 3.3 0.00067652 0 0.00067644 0 0.00067654 3.3 0.00067646 3.3 0.00067656 0 0.00067648 0 0.00067658 3.3 0.0006765 3.3 0.0006766 0 0.00067652 0 0.00067662 3.3 0.00067654 3.3 0.0006766399999999999 0 0.00067656 0 0.0006766599999999999 3.3 0.0006765800000000001 3.3 0.00067668 0 0.0006766000000000001 0 0.0006767 3.3 0.0006766200000000001 3.3 0.00067672 0 0.00067664 0 0.00067674 3.3 0.00067666 3.3 0.00067676 0 0.00067668 0 0.00067678 3.3 0.0006767 3.3 0.0006768 0 0.00067672 0 0.00067682 3.3 0.00067674 3.3 0.00067684 0 0.00067676 0 0.0006768599999999999 3.3 0.0006767800000000001 3.3 0.00067688 0 0.0006768000000000001 0 0.0006769 3.3 0.0006768200000000001 3.3 0.00067692 0 0.0006768400000000001 0 0.00067694 3.3 0.00067686 3.3 0.00067696 0 0.00067688 0 0.00067698 3.3 0.0006769 3.3 0.000677 0 0.00067692 0 0.00067702 3.3 0.00067694 3.3 0.00067704 0 0.00067696 0 0.0006770599999999999 3.3 0.00067698 3.3 0.0006770799999999999 0 0.0006770000000000001 0 0.0006771 3.3 0.0006770200000000001 3.3 0.00067712 0 0.0006770400000000001 0 0.00067714 3.3 0.00067706 3.3 0.00067716 0 0.00067708 0 0.00067718 3.3 0.0006771 3.3 0.0006772 0 0.00067712 0 0.00067722 3.3 0.00067714 3.3 0.00067724 0 0.00067716 0 0.00067726 3.3 0.00067718 3.3 0.0006772799999999999 0 0.0006772000000000001 0 0.0006773 3.3 0.0006772200000000001 3.3 0.00067732 0 0.0006772400000000001 0 0.00067734 3.3 0.0006772600000000001 3.3 0.00067736 0 0.00067728 0 0.00067738 3.3 0.0006773 3.3 0.0006774 0 0.00067732 0 0.00067742 3.3 0.00067734 3.3 0.00067744 0 0.00067736 0 0.00067746 3.3 0.00067738 3.3 0.0006774799999999999 0 0.0006774 0 0.0006774999999999999 3.3 0.0006774200000000001 3.3 0.00067752 0 0.0006774400000000001 0 0.00067754 3.3 0.0006774600000000001 3.3 0.00067756 0 0.00067748 0 0.00067758 3.3 0.0006775 3.3 0.0006776 0 0.00067752 0 0.00067762 3.3 0.00067754 3.3 0.00067764 0 0.00067756 0 0.00067766 3.3 0.00067758 3.3 0.00067768 0 0.0006776 0 0.0006776999999999999 3.3 0.0006776200000000001 3.3 0.00067772 0 0.0006776400000000001 0 0.00067774 3.3 0.0006776600000000001 3.3 0.00067776 0 0.0006776800000000001 0 0.00067778 3.3 0.0006777 3.3 0.0006778 0 0.00067772 0 0.00067782 3.3 0.00067774 3.3 0.00067784 0 0.00067776 0 0.00067786 3.3 0.00067778 3.3 0.00067788 0 0.0006778 0 0.0006778999999999999 3.3 0.00067782 3.3 0.0006779199999999999 0 0.0006778400000000001 0 0.00067794 3.3 0.0006778600000000001 3.3 0.00067796 0 0.0006778800000000001 0 0.00067798 3.3 0.0006779 3.3 0.000678 0 0.00067792 0 0.00067802 3.3 0.00067794 3.3 0.00067804 0 0.00067796 0 0.00067806 3.3 0.00067798 3.3 0.00067808 0 0.000678 0 0.0006781 3.3 0.00067802 3.3 0.0006781199999999999 0 0.0006780400000000001 0 0.00067814 3.3 0.0006780600000000001 3.3 0.00067816 0 0.0006780800000000001 0 0.00067818 3.3 0.0006781000000000001 3.3 0.0006782 0 0.00067812 0 0.00067822 3.3 0.00067814 3.3 0.00067824 0 0.00067816 0 0.00067826 3.3 0.00067818 3.3 0.00067828 0 0.0006782 0 0.0006783 3.3 0.00067822 3.3 0.0006783199999999999 0 0.00067824 0 0.0006783399999999999 3.3 0.0006782600000000001 3.3 0.00067836 0 0.0006782800000000001 0 0.00067838 3.3 0.0006783000000000001 3.3 0.0006784 0 0.00067832 0 0.00067842 3.3 0.00067834 3.3 0.00067844 0 0.00067836 0 0.00067846 3.3 0.00067838 3.3 0.00067848 0 0.0006784 0 0.0006785 3.3 0.00067842 3.3 0.00067852 0 0.00067844 0 0.0006785399999999999 3.3 0.0006784600000000001 3.3 0.00067856 0 0.0006784800000000001 0 0.00067858 3.3 0.0006785000000000001 3.3 0.0006786 0 0.0006785200000000001 0 0.00067862 3.3 0.00067854 3.3 0.00067864 0 0.00067856 0 0.00067866 3.3 0.00067858 3.3 0.00067868 0 0.0006786 0 0.0006787 3.3 0.00067862 3.3 0.00067872 0 0.00067864 0 0.0006787399999999999 3.3 0.0006786600000000001 3.3 0.00067876 0 0.0006786800000000001 0 0.00067878 3.3 0.0006787000000000001 3.3 0.0006788 0 0.0006787200000000001 0 0.00067882 3.3 0.00067874 3.3 0.00067884 0 0.00067876 0 0.00067886 3.3 0.00067878 3.3 0.00067888 0 0.0006788 0 0.0006789 3.3 0.00067882 3.3 0.00067892 0 0.00067884 0 0.00067894 3.3 0.00067886 3.3 0.0006789599999999999 0 0.0006788800000000001 0 0.00067898 3.3 0.0006789000000000001 3.3 0.000679 0 0.0006789200000000001 0 0.00067902 3.3 0.0006789400000000001 3.3 0.00067904 0 0.00067896 0 0.00067906 3.3 0.00067898 3.3 0.00067908 0 0.000679 0 0.0006791 3.3 0.00067902 3.3 0.00067912 0 0.00067904 0 0.00067914 3.3 0.00067906 3.3 0.0006791599999999999 0 0.0006790800000000001 0 0.00067918 3.3 0.0006791000000000001 3.3 0.0006792 0 0.0006791200000000001 0 0.00067922 3.3 0.0006791400000000001 3.3 0.00067924 0 0.00067916 0 0.00067926 3.3 0.00067918 3.3 0.00067928 0 0.0006792 0 0.0006793 3.3 0.00067922 3.3 0.00067932 0 0.00067924 0 0.00067934 3.3 0.00067926 3.3 0.00067936 0 0.00067928 0 0.0006793799999999999 3.3 0.0006793000000000001 3.3 0.0006794 0 0.0006793200000000001 0 0.00067942 3.3 0.0006793400000000001 3.3 0.00067944 0 0.0006793600000000001 0 0.00067946 3.3 0.00067938 3.3 0.00067948 0 0.0006794 0 0.0006795 3.3 0.00067942 3.3 0.00067952 0 0.00067944 0 0.00067954 3.3 0.00067946 3.3 0.00067956 0 0.00067948 0 0.0006795799999999999 3.3 0.0006795000000000001 3.3 0.0006796 0 0.0006795200000000001 0 0.00067962 3.3 0.0006795400000000001 3.3 0.00067964 0 0.0006795600000000001 0 0.00067966 3.3 0.00067958 3.3 0.00067968 0 0.0006796 0 0.0006797 3.3 0.00067962 3.3 0.00067972 0 0.00067964 0 0.00067974 3.3 0.00067966 3.3 0.00067976 0 0.00067968 0 0.00067978 3.3 0.0006797 3.3 0.0006797999999999999 0 0.0006797200000000001 0 0.00067982 3.3 0.0006797400000000001 3.3 0.00067984 0 0.0006797600000000001 0 0.00067986 3.3 0.0006797800000000001 3.3 0.00067988 0 0.0006798 0 0.0006799 3.3 0.00067982 3.3 0.00067992 0 0.00067984 0 0.00067994 3.3 0.00067986 3.3 0.00067996 0 0.00067988 0 0.00067998 3.3 0.0006799 3.3 0.0006799999999999999 0 0.0006799200000000001 0 0.00068002 3.3 0.0006799400000000001 3.3 0.00068004 0 0.0006799600000000001 0 0.00068006 3.3 0.0006799800000000001 3.3 0.00068008 0 0.00068 0 0.0006801 3.3 0.00068002 3.3 0.00068012 0 0.00068004 0 0.00068014 3.3 0.00068006 3.3 0.00068016 0 0.00068008 0 0.00068018 3.3 0.0006801 3.3 0.0006801999999999999 0 0.00068012 0 0.0006802199999999999 3.3 0.0006801400000000001 3.3 0.00068024 0 0.0006801600000000001 0 0.00068026 3.3 0.0006801800000000001 3.3 0.00068028 0 0.0006802 0 0.0006803 3.3 0.00068022 3.3 0.00068032 0 0.00068024 0 0.00068034 3.3 0.00068026 3.3 0.00068036 0 0.00068028 0 0.00068038 3.3 0.0006803 3.3 0.0006804 0 0.00068032 0 0.0006804199999999999 3.3 0.0006803400000000001 3.3 0.00068044 0 0.0006803600000000001 0 0.00068046 3.3 0.0006803800000000001 3.3 0.00068048 0 0.0006804000000000001 0 0.0006805 3.3 0.00068042 3.3 0.00068052 0 0.00068044 0 0.00068054 3.3 0.00068046 3.3 0.00068056 0 0.00068048 0 0.00068058 3.3 0.0006805 3.3 0.0006806 0 0.00068052 0 0.0006806199999999999 3.3 0.00068054 3.3 0.0006806399999999999 0 0.0006805600000000001 0 0.00068066 3.3 0.0006805800000000001 3.3 0.00068068 0 0.0006806000000000001 0 0.0006807 3.3 0.00068062 3.3 0.00068072 0 0.00068064 0 0.00068074 3.3 0.00068066 3.3 0.00068076 0 0.00068068 0 0.00068078 3.3 0.0006807 3.3 0.0006808 0 0.00068072 0 0.00068082 3.3 0.00068074 3.3 0.0006808399999999999 0 0.0006807600000000001 0 0.00068086 3.3 0.0006807800000000001 3.3 0.00068088 0 0.0006808000000000001 0 0.0006809 3.3 0.0006808200000000001 3.3 0.00068092 0 0.00068084 0 0.00068094 3.3 0.00068086 3.3 0.00068096 0 0.00068088 0 0.00068098 3.3 0.0006809 3.3 0.000681 0 0.00068092 0 0.00068102 3.3 0.00068094 3.3 0.0006810399999999999 0 0.00068096 0 0.0006810599999999999 3.3 0.0006809800000000001 3.3 0.00068108 0 0.0006810000000000001 0 0.0006811 3.3 0.0006810200000000001 3.3 0.00068112 0 0.00068104 0 0.00068114 3.3 0.00068106 3.3 0.00068116 0 0.00068108 0 0.00068118 3.3 0.0006811 3.3 0.0006812 0 0.00068112 0 0.00068122 3.3 0.00068114 3.3 0.00068124 0 0.00068116 0 0.0006812599999999999 3.3 0.0006811800000000001 3.3 0.00068128 0 0.0006812000000000001 0 0.0006813 3.3 0.0006812200000000001 3.3 0.00068132 0 0.0006812400000000001 0 0.00068134 3.3 0.00068126 3.3 0.00068136 0 0.00068128 0 0.00068138 3.3 0.0006813 3.3 0.0006814 0 0.00068132 0 0.00068142 3.3 0.00068134 3.3 0.00068144 0 0.00068136 0 0.0006814599999999999 3.3 0.00068138 3.3 0.0006814799999999999 0 0.0006814000000000001 0 0.0006815 3.3 0.0006814200000000001 3.3 0.00068152 0 0.0006814400000000001 0 0.00068154 3.3 0.00068146 3.3 0.00068156 0 0.00068148 0 0.00068158 3.3 0.0006815 3.3 0.0006816 0 0.00068152 0 0.00068162 3.3 0.00068154 3.3 0.00068164 0 0.00068156 0 0.00068166 3.3 0.00068158 3.3 0.0006816799999999999 0 0.0006816000000000001 0 0.0006817 3.3 0.0006816200000000001 3.3 0.00068172 0 0.0006816400000000001 0 0.00068174 3.3 0.0006816600000000001 3.3 0.00068176 0 0.00068168 0 0.00068178 3.3 0.0006817 3.3 0.0006818 0 0.00068172 0 0.00068182 3.3 0.00068174 3.3 0.00068184 0 0.00068176 0 0.00068186 3.3 0.00068178 3.3 0.0006818799999999999 0 0.0006818 0 0.0006818999999999999 3.3 0.0006818200000000001 3.3 0.00068192 0 0.0006818400000000001 0 0.00068194 3.3 0.0006818600000000001 3.3 0.00068196 0 0.00068188 0 0.00068198 3.3 0.0006819 3.3 0.000682 0 0.00068192 0 0.00068202 3.3 0.00068194 3.3 0.00068204 0 0.00068196 0 0.00068206 3.3 0.00068198 3.3 0.00068208 0 0.000682 0 0.0006820999999999999 3.3 0.0006820200000000001 3.3 0.00068212 0 0.0006820400000000001 0 0.00068214 3.3 0.0006820600000000001 3.3 0.00068216 0 0.0006820800000000001 0 0.00068218 3.3 0.0006821 3.3 0.0006822 0 0.00068212 0 0.00068222 3.3 0.00068214 3.3 0.00068224 0 0.00068216 0 0.00068226 3.3 0.00068218 3.3 0.00068228 0 0.0006822 0 0.0006822999999999999 3.3 0.0006822200000000001 3.3 0.00068232 0 0.0006822400000000001 0 0.00068234 3.3 0.0006822600000000001 3.3 0.00068236 0 0.0006822800000000001 0 0.00068238 3.3 0.0006823 3.3 0.0006824 0 0.00068232 0 0.00068242 3.3 0.00068234 3.3 0.00068244 0 0.00068236 0 0.00068246 3.3 0.00068238 3.3 0.00068248 0 0.0006824 0 0.0006825 3.3 0.00068242 3.3 0.0006825199999999999 0 0.0006824400000000001 0 0.00068254 3.3 0.0006824600000000001 3.3 0.00068256 0 0.0006824800000000001 0 0.00068258 3.3 0.0006825000000000001 3.3 0.0006826 0 0.00068252 0 0.00068262 3.3 0.00068254 3.3 0.00068264 0 0.00068256 0 0.00068266 3.3 0.00068258 3.3 0.00068268 0 0.0006826 0 0.0006827 3.3 0.00068262 3.3 0.0006827199999999999 0 0.0006826400000000001 0 0.00068274 3.3 0.0006826600000000001 3.3 0.00068276 0 0.0006826800000000001 0 0.00068278 3.3 0.0006827000000000001 3.3 0.0006828 0 0.00068272 0 0.00068282 3.3 0.00068274 3.3 0.00068284 0 0.00068276 0 0.00068286 3.3 0.00068278 3.3 0.00068288 0 0.0006828 0 0.0006829 3.3 0.00068282 3.3 0.00068292 0 0.00068284 0 0.0006829399999999999 3.3 0.0006828600000000001 3.3 0.00068296 0 0.0006828800000000001 0 0.00068298 3.3 0.0006829000000000001 3.3 0.000683 0 0.0006829200000000001 0 0.00068302 3.3 0.00068294 3.3 0.00068304 0 0.00068296 0 0.00068306 3.3 0.00068298 3.3 0.00068308 0 0.000683 0 0.0006831 3.3 0.00068302 3.3 0.00068312 0 0.00068304 0 0.0006831399999999999 3.3 0.0006830600000000001 3.3 0.00068316 0 0.0006830800000000001 0 0.00068318 3.3 0.0006831000000000001 3.3 0.0006832 0 0.0006831200000000001 0 0.00068322 3.3 0.00068314 3.3 0.00068324 0 0.00068316 0 0.00068326 3.3 0.00068318 3.3 0.00068328 0 0.0006832 0 0.0006833 3.3 0.00068322 3.3 0.00068332 0 0.00068324 0 0.0006833399999999999 3.3 0.00068326 3.3 0.0006833599999999999 0 0.0006832800000000001 0 0.00068338 3.3 0.0006833000000000001 3.3 0.0006834 0 0.0006833200000000001 0 0.00068342 3.3 0.00068334 3.3 0.00068344 0 0.00068336 0 0.00068346 3.3 0.00068338 3.3 0.00068348 0 0.0006834 0 0.0006835 3.3 0.00068342 3.3 0.00068352 0 0.00068344 0 0.00068354 3.3 0.00068346 3.3 0.0006835599999999999 0 0.0006834800000000001 0 0.00068358 3.3 0.0006835000000000001 3.3 0.0006836 0 0.0006835200000000001 0 0.00068362 3.3 0.0006835400000000001 3.3 0.00068364 0 0.00068356 0 0.00068366 3.3 0.00068358 3.3 0.00068368 0 0.0006836 0 0.0006837 3.3 0.00068362 3.3 0.00068372 0 0.00068364 0 0.00068374 3.3 0.00068366 3.3 0.0006837599999999999 0 0.00068368 0 0.0006837799999999999 3.3 0.0006837000000000001 3.3 0.0006838 0 0.0006837200000000001 0 0.00068382 3.3 0.0006837400000000001 3.3 0.00068384 0 0.00068376 0 0.00068386 3.3 0.00068378 3.3 0.00068388 0 0.0006838 0 0.0006839 3.3 0.00068382 3.3 0.00068392 0 0.00068384 0 0.00068394 3.3 0.00068386 3.3 0.00068396 0 0.00068388 0 0.0006839799999999999 3.3 0.0006839000000000001 3.3 0.000684 0 0.0006839200000000001 0 0.00068402 3.3 0.0006839400000000001 3.3 0.00068404 0 0.0006839600000000001 0 0.00068406 3.3 0.00068398 3.3 0.00068408 0 0.000684 0 0.0006841 3.3 0.00068402 3.3 0.00068412 0 0.00068404 0 0.00068414 3.3 0.00068406 3.3 0.00068416 0 0.00068408 0 0.0006841799999999999 3.3 0.0006841 3.3 0.0006841999999999999 0 0.0006841200000000001 0 0.00068422 3.3 0.0006841400000000001 3.3 0.00068424 0 0.0006841600000000001 0 0.00068426 3.3 0.00068418 3.3 0.00068428 0 0.0006842 0 0.0006843 3.3 0.00068422 3.3 0.00068432 0 0.00068424 0 0.00068434 3.3 0.00068426 3.3 0.00068436 0 0.00068428 0 0.00068438 3.3 0.0006843 3.3 0.0006843999999999999 0 0.0006843200000000001 0 0.00068442 3.3 0.0006843400000000001 3.3 0.00068444 0 0.0006843600000000001 0 0.00068446 3.3 0.0006843800000000001 3.3 0.00068448 0 0.0006844 0 0.0006845 3.3 0.00068442 3.3 0.00068452 0 0.00068444 0 0.00068454 3.3 0.00068446 3.3 0.00068456 0 0.00068448 0 0.00068458 3.3 0.0006845 3.3 0.0006845999999999999 0 0.00068452 0 0.0006846199999999999 3.3 0.0006845400000000001 3.3 0.00068464 0 0.0006845600000000001 0 0.00068466 3.3 0.0006845800000000001 3.3 0.00068468 0 0.0006846 0 0.0006847 3.3 0.00068462 3.3 0.00068472 0 0.00068464 0 0.00068474 3.3 0.00068466 3.3 0.00068476 0 0.00068468 0 0.00068478 3.3 0.0006847 3.3 0.0006848 0 0.00068472 0 0.0006848199999999999 3.3 0.0006847400000000001 3.3 0.00068484 0 0.0006847600000000001 0 0.00068486 3.3 0.0006847800000000001 3.3 0.00068488 0 0.0006848000000000001 0 0.0006849 3.3 0.00068482 3.3 0.00068492 0 0.00068484 0 0.00068494 3.3 0.00068486 3.3 0.00068496 0 0.00068488 0 0.00068498 3.3 0.0006849 3.3 0.000685 0 0.00068492 0 0.0006850199999999999 3.3 0.00068494 3.3 0.0006850399999999999 0 0.0006849600000000001 0 0.00068506 3.3 0.0006849800000000001 3.3 0.00068508 0 0.0006850000000000001 0 0.0006851 3.3 0.00068502 3.3 0.00068512 0 0.00068504 0 0.00068514 3.3 0.00068506 3.3 0.00068516 0 0.00068508 0 0.00068518 3.3 0.0006851 3.3 0.0006852 0 0.00068512 0 0.00068522 3.3 0.00068514 3.3 0.0006852399999999999 0 0.0006851600000000001 0 0.00068526 3.3 0.0006851800000000001 3.3 0.00068528 0 0.0006852000000000001 0 0.0006853 3.3 0.0006852200000000001 3.3 0.00068532 0 0.00068524 0 0.00068534 3.3 0.00068526 3.3 0.00068536 0 0.00068528 0 0.00068538 3.3 0.0006853 3.3 0.0006854 0 0.00068532 0 0.00068542 3.3 0.00068534 3.3 0.0006854399999999999 0 0.00068536 0 0.0006854599999999999 3.3 0.0006853800000000001 3.3 0.00068548 0 0.0006854000000000001 0 0.0006855 3.3 0.0006854200000000001 3.3 0.00068552 0 0.00068544 0 0.00068554 3.3 0.00068546 3.3 0.00068556 0 0.00068548 0 0.00068558 3.3 0.0006855 3.3 0.0006856 0 0.00068552 0 0.00068562 3.3 0.00068554 3.3 0.00068564 0 0.00068556 0 0.0006856599999999999 3.3 0.0006855800000000001 3.3 0.00068568 0 0.0006856000000000001 0 0.0006857 3.3 0.0006856200000000001 3.3 0.00068572 0 0.0006856400000000001 0 0.00068574 3.3 0.00068566 3.3 0.00068576 0 0.00068568 0 0.00068578 3.3 0.0006857 3.3 0.0006858 0 0.00068572 0 0.00068582 3.3 0.00068574 3.3 0.00068584 0 0.00068576 0 0.0006858599999999999 3.3 0.0006857800000000001 3.3 0.00068588 0 0.0006858000000000001 0 0.0006859 3.3 0.0006858200000000001 3.3 0.00068592 0 0.0006858400000000001 0 0.00068594 3.3 0.00068586 3.3 0.00068596 0 0.00068588 0 0.00068598 3.3 0.0006859 3.3 0.000686 0 0.00068592 0 0.00068602 3.3 0.00068594 3.3 0.00068604 0 0.00068596 0 0.00068606 3.3 0.00068598 3.3 0.0006860799999999999 0 0.0006860000000000001 0 0.0006861 3.3 0.0006860200000000001 3.3 0.00068612 0 0.0006860400000000001 0 0.00068614 3.3 0.0006860600000000001 3.3 0.00068616 0 0.00068608 0 0.00068618 3.3 0.0006861 3.3 0.0006862 0 0.00068612 0 0.00068622 3.3 0.00068614 3.3 0.00068624 0 0.00068616 0 0.00068626 3.3 0.00068618 3.3 0.0006862799999999999 0 0.0006862000000000001 0 0.0006863 3.3 0.0006862200000000001 3.3 0.00068632 0 0.0006862400000000001 0 0.00068634 3.3 0.0006862600000000001 3.3 0.00068636 0 0.00068628 0 0.00068638 3.3 0.0006863 3.3 0.0006864 0 0.00068632 0 0.00068642 3.3 0.00068634 3.3 0.00068644 0 0.00068636 0 0.00068646 3.3 0.00068638 3.3 0.00068648 0 0.0006864 0 0.0006864999999999999 3.3 0.0006864200000000001 3.3 0.00068652 0 0.0006864400000000001 0 0.00068654 3.3 0.0006864600000000001 3.3 0.00068656 0 0.0006864800000000001 0 0.00068658 3.3 0.0006865 3.3 0.0006866 0 0.00068652 0 0.00068662 3.3 0.00068654 3.3 0.00068664 0 0.00068656 0 0.00068666 3.3 0.00068658 3.3 0.00068668 0 0.0006866 0 0.0006866999999999999 3.3 0.0006866200000000001 3.3 0.00068672 0 0.0006866400000000001 0 0.00068674 3.3 0.0006866600000000001 3.3 0.00068676 0 0.0006866800000000001 0 0.00068678 3.3 0.0006867 3.3 0.0006868 0 0.00068672 0 0.00068682 3.3 0.00068674 3.3 0.00068684 0 0.00068676 0 0.00068686 3.3 0.00068678 3.3 0.00068688 0 0.0006868 0 0.0006868999999999999 3.3 0.00068682 3.3 0.0006869199999999999 0 0.0006868400000000001 0 0.00068694 3.3 0.0006868600000000001 3.3 0.00068696 0 0.0006868800000000001 0 0.00068698 3.3 0.0006869 3.3 0.000687 0 0.00068692 0 0.00068702 3.3 0.00068694 3.3 0.00068704 0 0.00068696 0 0.00068706 3.3 0.00068698 3.3 0.00068708 0 0.000687 0 0.0006871 3.3 0.00068702 3.3 0.0006871199999999999 0 0.0006870400000000001 0 0.00068714 3.3 0.0006870600000000001 3.3 0.00068716 0 0.0006870800000000001 0 0.00068718 3.3 0.0006871000000000001 3.3 0.0006872 0 0.00068712 0 0.00068722 3.3 0.00068714 3.3 0.00068724 0 0.00068716 0 0.00068726 3.3 0.00068718 3.3 0.00068728 0 0.0006872 0 0.0006873 3.3 0.00068722 3.3 0.0006873199999999999 0 0.00068724 0 0.0006873399999999999 3.3 0.0006872600000000001 3.3 0.00068736 0 0.0006872800000000001 0 0.00068738 3.3 0.0006873000000000001 3.3 0.0006874 0 0.00068732 0 0.00068742 3.3 0.00068734 3.3 0.00068744 0 0.00068736 0 0.00068746 3.3 0.00068738 3.3 0.00068748 0 0.0006874 0 0.0006875 3.3 0.00068742 3.3 0.00068752 0 0.00068744 0 0.0006875399999999999 3.3 0.0006874600000000001 3.3 0.00068756 0 0.0006874800000000001 0 0.00068758 3.3 0.0006875000000000001 3.3 0.0006876 0 0.0006875200000000001 0 0.00068762 3.3 0.00068754 3.3 0.00068764 0 0.00068756 0 0.00068766 3.3 0.00068758 3.3 0.00068768 0 0.0006876 0 0.0006877 3.3 0.00068762 3.3 0.00068772 0 0.00068764 0 0.0006877399999999999 3.3 0.00068766 3.3 0.0006877599999999999 0 0.0006876800000000001 0 0.00068778 3.3 0.0006877000000000001 3.3 0.0006878 0 0.0006877200000000001 0 0.00068782 3.3 0.00068774 3.3 0.00068784 0 0.00068776 0 0.00068786 3.3 0.00068778 3.3 0.00068788 0 0.0006878 0 0.0006879 3.3 0.00068782 3.3 0.00068792 0 0.00068784 0 0.00068794 3.3 0.00068786 3.3 0.0006879599999999999 0 0.0006878800000000001 0 0.00068798 3.3 0.0006879000000000001 3.3 0.000688 0 0.0006879200000000001 0 0.00068802 3.3 0.0006879400000000001 3.3 0.00068804 0 0.00068796 0 0.00068806 3.3 0.00068798 3.3 0.00068808 0 0.000688 0 0.0006881 3.3 0.00068802 3.3 0.00068812 0 0.00068804 0 0.00068814 3.3 0.00068806 3.3 0.0006881599999999999 0 0.00068808 0 0.0006881799999999999 3.3 0.0006881000000000001 3.3 0.0006882 0 0.0006881200000000001 0 0.00068822 3.3 0.0006881400000000001 3.3 0.00068824 0 0.00068816 0 0.00068826 3.3 0.00068818 3.3 0.00068828 0 0.0006882 0 0.0006883 3.3 0.00068822 3.3 0.00068832 0 0.00068824 0 0.00068834 3.3 0.00068826 3.3 0.00068836 0 0.00068828 0 0.0006883799999999999 3.3 0.0006883000000000001 3.3 0.0006884 0 0.0006883200000000001 0 0.00068842 3.3 0.0006883400000000001 3.3 0.00068844 0 0.0006883600000000001 0 0.00068846 3.3 0.00068838 3.3 0.00068848 0 0.0006884 0 0.0006885 3.3 0.00068842 3.3 0.00068852 0 0.00068844 0 0.00068854 3.3 0.00068846 3.3 0.00068856 0 0.00068848 0 0.0006885799999999999 3.3 0.0006885 3.3 0.0006885999999999999 0 0.0006885200000000001 0 0.00068862 3.3 0.0006885400000000001 3.3 0.00068864 0 0.0006885600000000001 0 0.00068866 3.3 0.00068858 3.3 0.00068868 0 0.0006886 0 0.0006887 3.3 0.00068862 3.3 0.00068872 0 0.00068864 0 0.00068874 3.3 0.00068866 3.3 0.00068876 0 0.00068868 0 0.00068878 3.3 0.0006887 3.3 0.0006887999999999999 0 0.0006887200000000001 0 0.00068882 3.3 0.0006887400000000001 3.3 0.00068884 0 0.0006887600000000001 0 0.00068886 3.3 0.0006887800000000001 3.3 0.00068888 0 0.0006888 0 0.0006889 3.3 0.00068882 3.3 0.00068892 0 0.00068884 0 0.00068894 3.3 0.00068886 3.3 0.00068896 0 0.00068888 0 0.00068898 3.3 0.0006889 3.3 0.0006889999999999999 0 0.00068892 0 0.0006890199999999999 3.3 0.0006889400000000001 3.3 0.00068904 0 0.0006889600000000001 0 0.00068906 3.3 0.0006889800000000001 3.3 0.00068908 0 0.000689 0 0.0006891 3.3 0.00068902 3.3 0.00068912 0 0.00068904 0 0.00068914 3.3 0.00068906 3.3 0.00068916 0 0.00068908 0 0.00068918 3.3 0.0006891 3.3 0.0006892 0 0.00068912 0 0.0006892199999999999 3.3 0.0006891400000000001 3.3 0.00068924 0 0.0006891600000000001 0 0.00068926 3.3 0.0006891800000000001 3.3 0.00068928 0 0.0006892000000000001 0 0.0006893 3.3 0.00068922 3.3 0.00068932 0 0.00068924 0 0.00068934 3.3 0.00068926 3.3 0.00068936 0 0.00068928 0 0.00068938 3.3 0.0006893 3.3 0.0006894 0 0.00068932 0 0.0006894199999999999 3.3 0.0006893400000000001 3.3 0.00068944 0 0.0006893600000000001 0 0.00068946 3.3 0.0006893800000000001 3.3 0.00068948 0 0.0006894000000000001 0 0.0006895 3.3 0.00068942 3.3 0.00068952 0 0.00068944 0 0.00068954 3.3 0.00068946 3.3 0.00068956 0 0.00068948 0 0.00068958 3.3 0.0006895 3.3 0.0006896 0 0.00068952 0 0.00068962 3.3 0.00068954 3.3 0.0006896399999999999 0 0.0006895600000000001 0 0.00068966 3.3 0.0006895800000000001 3.3 0.00068968 0 0.0006896000000000001 0 0.0006897 3.3 0.0006896200000000001 3.3 0.00068972 0 0.00068964 0 0.00068974 3.3 0.00068966 3.3 0.00068976 0 0.00068968 0 0.00068978 3.3 0.0006897 3.3 0.0006898 0 0.00068972 0 0.00068982 3.3 0.00068974 3.3 0.0006898399999999999 0 0.0006897600000000001 0 0.00068986 3.3 0.0006897800000000001 3.3 0.00068988 0 0.0006898000000000001 0 0.0006899 3.3 0.0006898200000000001 3.3 0.00068992 0 0.00068984 0 0.00068994 3.3 0.00068986 3.3 0.00068996 0 0.00068988 0 0.00068998 3.3 0.0006899 3.3 0.00069 0 0.00068992 0 0.00069002 3.3 0.00068994 3.3 0.00069004 0 0.00068996 0 0.0006900599999999999 3.3 0.0006899800000000001 3.3 0.00069008 0 0.0006900000000000001 0 0.0006901 3.3 0.0006900200000000001 3.3 0.00069012 0 0.0006900400000000001 0 0.00069014 3.3 0.00069006 3.3 0.00069016 0 0.00069008 0 0.00069018 3.3 0.0006901 3.3 0.0006902 0 0.00069012 0 0.00069022 3.3 0.00069014 3.3 0.00069024 0 0.00069016 0 0.0006902599999999999 3.3 0.0006901800000000001 3.3 0.00069028 0 0.0006902000000000001 0 0.0006903 3.3 0.0006902200000000001 3.3 0.00069032 0 0.0006902400000000001 0 0.00069034 3.3 0.00069026 3.3 0.00069036 0 0.00069028 0 0.00069038 3.3 0.0006903 3.3 0.0006904 0 0.00069032 0 0.00069042 3.3 0.00069034 3.3 0.00069044 0 0.00069036 0 0.0006904599999999999 3.3 0.00069038 3.3 0.0006904799999999999 0 0.0006904000000000001 0 0.0006905 3.3 0.0006904200000000001 3.3 0.00069052 0 0.0006904400000000001 0 0.00069054 3.3 0.00069046 3.3 0.00069056 0 0.00069048 0 0.00069058 3.3 0.0006905 3.3 0.0006906 0 0.00069052 0 0.00069062 3.3 0.00069054 3.3 0.00069064 0 0.00069056 0 0.00069066 3.3 0.00069058 3.3 0.0006906799999999999 0 0.0006906000000000001 0 0.0006907 3.3 0.0006906200000000001 3.3 0.00069072 0 0.0006906400000000001 0 0.00069074 3.3 0.0006906600000000001 3.3 0.00069076 0 0.00069068 0 0.00069078 3.3 0.0006907 3.3 0.0006908 0 0.00069072 0 0.00069082 3.3 0.00069074 3.3 0.00069084 0 0.00069076 0 0.00069086 3.3 0.00069078 3.3 0.0006908799999999999 0 0.0006908 0 0.0006908999999999999 3.3 0.0006908200000000001 3.3 0.00069092 0 0.0006908400000000001 0 0.00069094 3.3 0.0006908600000000001 3.3 0.00069096 0 0.00069088 0 0.00069098 3.3 0.0006909 3.3 0.000691 0 0.00069092 0 0.00069102 3.3 0.00069094 3.3 0.00069104 0 0.00069096 0 0.00069106 3.3 0.00069098 3.3 0.00069108 0 0.000691 0 0.0006910999999999999 3.3 0.0006910200000000001 3.3 0.00069112 0 0.0006910400000000001 0 0.00069114 3.3 0.0006910600000000001 3.3 0.00069116 0 0.0006910800000000001 0 0.00069118 3.3 0.0006911 3.3 0.0006912 0 0.00069112 0 0.00069122 3.3 0.00069114 3.3 0.00069124 0 0.00069116 0 0.00069126 3.3 0.00069118 3.3 0.00069128 0 0.0006912 0 0.0006912999999999999 3.3 0.00069122 3.3 0.0006913199999999999 0 0.0006912400000000001 0 0.00069134 3.3 0.0006912600000000001 3.3 0.00069136 0 0.0006912800000000001 0 0.00069138 3.3 0.0006913 3.3 0.0006914 0 0.00069132 0 0.00069142 3.3 0.00069134 3.3 0.00069144 0 0.00069136 0 0.00069146 3.3 0.00069138 3.3 0.00069148 0 0.0006914 0 0.0006915 3.3 0.00069142 3.3 0.0006915199999999999 0 0.0006914400000000001 0 0.00069154 3.3 0.0006914600000000001 3.3 0.00069156 0 0.0006914800000000001 0 0.00069158 3.3 0.0006915000000000001 3.3 0.0006916 0 0.00069152 0 0.00069162 3.3 0.00069154 3.3 0.00069164 0 0.00069156 0 0.00069166 3.3 0.00069158 3.3 0.00069168 0 0.0006916 0 0.0006917 3.3 0.00069162 3.3 0.0006917199999999999 0 0.00069164 0 0.0006917399999999999 3.3 0.0006916600000000001 3.3 0.00069176 0 0.0006916800000000001 0 0.00069178 3.3 0.0006917000000000001 3.3 0.0006918 0 0.00069172 0 0.00069182 3.3 0.00069174 3.3 0.00069184 0 0.00069176 0 0.00069186 3.3 0.00069178 3.3 0.00069188 0 0.0006918 0 0.0006919 3.3 0.00069182 3.3 0.00069192 0 0.00069184 0 0.0006919399999999999 3.3 0.0006918600000000001 3.3 0.00069196 0 0.0006918800000000001 0 0.00069198 3.3 0.0006919000000000001 3.3 0.000692 0 0.0006919200000000001 0 0.00069202 3.3 0.00069194 3.3 0.00069204 0 0.00069196 0 0.00069206 3.3 0.00069198 3.3 0.00069208 0 0.000692 0 0.0006921 3.3 0.00069202 3.3 0.00069212 0 0.00069204 0 0.0006921399999999999 3.3 0.00069206 3.3 0.0006921599999999999 0 0.0006920800000000001 0 0.00069218 3.3 0.0006921000000000001 3.3 0.0006922 0 0.0006921200000000001 0 0.00069222 3.3 0.00069214 3.3 0.00069224 0 0.00069216 0 0.00069226 3.3 0.00069218 3.3 0.00069228 0 0.0006922 0 0.0006923 3.3 0.00069222 3.3 0.00069232 0 0.00069224 0 0.00069234 3.3 0.00069226 3.3 0.0006923599999999999 0 0.0006922800000000001 0 0.00069238 3.3 0.0006923000000000001 3.3 0.0006924 0 0.0006923200000000001 0 0.00069242 3.3 0.0006923400000000001 3.3 0.00069244 0 0.00069236 0 0.00069246 3.3 0.00069238 3.3 0.00069248 0 0.0006924 0 0.0006925 3.3 0.00069242 3.3 0.00069252 0 0.00069244 0 0.00069254 3.3 0.00069246 3.3 0.0006925599999999999 0 0.0006924800000000001 0 0.00069258 3.3 0.0006925000000000001 3.3 0.0006926 0 0.0006925200000000001 0 0.00069262 3.3 0.0006925400000000001 3.3 0.00069264 0 0.00069256 0 0.00069266 3.3 0.00069258 3.3 0.00069268 0 0.0006926 0 0.0006927 3.3 0.00069262 3.3 0.00069272 0 0.00069264 0 0.00069274 3.3 0.00069266 3.3 0.00069276 0 0.00069268 0 0.0006927799999999999 3.3 0.0006927000000000001 3.3 0.0006928 0 0.0006927200000000001 0 0.00069282 3.3 0.0006927400000000001 3.3 0.00069284 0 0.0006927600000000001 0 0.00069286 3.3 0.00069278 3.3 0.00069288 0 0.0006928 0 0.0006929 3.3 0.00069282 3.3 0.00069292 0 0.00069284 0 0.00069294 3.3 0.00069286 3.3 0.00069296 0 0.00069288 0 0.0006929799999999999 3.3 0.0006929000000000001 3.3 0.000693 0 0.0006929200000000001 0 0.00069302 3.3 0.0006929400000000001 3.3 0.00069304 0 0.0006929600000000001 0 0.00069306 3.3 0.00069298 3.3 0.00069308 0 0.000693 0 0.0006931 3.3 0.00069302 3.3 0.00069312 0 0.00069304 0 0.00069314 3.3 0.00069306 3.3 0.00069316 0 0.00069308 0 0.00069318 3.3 0.0006931 3.3 0.0006931999999999999 0 0.0006931200000000001 0 0.00069322 3.3 0.0006931400000000001 3.3 0.00069324 0 0.0006931600000000001 0 0.00069326 3.3 0.0006931800000000001 3.3 0.00069328 0 0.0006932 0 0.0006933 3.3 0.00069322 3.3 0.00069332 0 0.00069324 0 0.00069334 3.3 0.00069326 3.3 0.00069336 0 0.00069328 0 0.00069338 3.3 0.0006933 3.3 0.0006933999999999999 0 0.0006933200000000001 0 0.00069342 3.3 0.0006933400000000001 3.3 0.00069344 0 0.0006933600000000001 0 0.00069346 3.3 0.0006933800000000001 3.3 0.00069348 0 0.0006934 0 0.0006935 3.3 0.00069342 3.3 0.00069352 0 0.00069344 0 0.00069354 3.3 0.00069346 3.3 0.00069356 0 0.00069348 0 0.00069358 3.3 0.0006935 3.3 0.0006935999999999999 0 0.00069352 0 0.0006936199999999999 3.3 0.0006935400000000001 3.3 0.00069364 0 0.0006935600000000001 0 0.00069366 3.3 0.0006935800000000001 3.3 0.00069368 0 0.0006936 0 0.0006937 3.3 0.00069362 3.3 0.00069372 0 0.00069364 0 0.00069374 3.3 0.00069366 3.3 0.00069376 0 0.00069368 0 0.00069378 3.3 0.0006937 3.3 0.0006938 0 0.00069372 0 0.0006938199999999999 3.3 0.0006937400000000001 3.3 0.00069384 0 0.0006937600000000001 0 0.00069386 3.3 0.0006937800000000001 3.3 0.00069388 0 0.0006938000000000001 0 0.0006939 3.3 0.00069382 3.3 0.00069392 0 0.00069384 0 0.00069394 3.3 0.00069386 3.3 0.00069396 0 0.00069388 0 0.00069398 3.3 0.0006939 3.3 0.000694 0 0.00069392 0 0.0006940199999999999 3.3 0.00069394 3.3 0.0006940399999999999 0 0.0006939600000000001 0 0.00069406 3.3 0.0006939800000000001 3.3 0.00069408 0 0.0006940000000000001 0 0.0006941 3.3 0.00069402 3.3 0.00069412 0 0.00069404 0 0.00069414 3.3 0.00069406 3.3 0.00069416 0 0.00069408 0 0.00069418 3.3 0.0006941 3.3 0.0006942 0 0.00069412 0 0.00069422 3.3 0.00069414 3.3 0.0006942399999999999 0 0.0006941600000000001 0 0.00069426 3.3 0.0006941800000000001 3.3 0.00069428 0 0.0006942000000000001 0 0.0006943 3.3 0.0006942200000000001 3.3 0.00069432 0 0.00069424 0 0.00069434 3.3 0.00069426 3.3 0.00069436 0 0.00069428 0 0.00069438 3.3 0.0006943 3.3 0.0006944 0 0.00069432 0 0.00069442 3.3 0.00069434 3.3 0.0006944399999999999 0 0.00069436 0 0.0006944599999999999 3.3 0.0006943800000000001 3.3 0.00069448 0 0.0006944000000000001 0 0.0006945 3.3 0.0006944200000000001 3.3 0.00069452 0 0.00069444 0 0.00069454 3.3 0.00069446 3.3 0.00069456 0 0.00069448 0 0.00069458 3.3 0.0006945 3.3 0.0006946 0 0.00069452 0 0.00069462 3.3 0.00069454 3.3 0.00069464 0 0.00069456 0 0.0006946599999999999 3.3 0.0006945800000000001 3.3 0.00069468 0 0.0006946000000000001 0 0.0006947 3.3 0.0006946200000000001 3.3 0.00069472 0 0.0006946400000000001 0 0.00069474 3.3 0.00069466 3.3 0.00069476 0 0.00069468 0 0.00069478 3.3 0.0006947 3.3 0.0006948 0 0.00069472 0 0.00069482 3.3 0.00069474 3.3 0.00069484 0 0.00069476 0 0.0006948599999999999 3.3 0.00069478 3.3 0.0006948799999999999 0 0.0006948000000000001 0 0.0006949 3.3 0.0006948200000000001 3.3 0.00069492 0 0.0006948400000000001 0 0.00069494 3.3 0.00069486 3.3 0.00069496 0 0.00069488 0 0.00069498 3.3 0.0006949 3.3 0.000695 0 0.00069492 0 0.00069502 3.3 0.00069494 3.3 0.00069504 0 0.00069496 0 0.00069506 3.3 0.00069498 3.3 0.0006950799999999999 0 0.0006950000000000001 0 0.0006951 3.3 0.0006950200000000001 3.3 0.00069512 0 0.0006950400000000001 0 0.00069514 3.3 0.0006950600000000001 3.3 0.00069516 0 0.00069508 0 0.00069518 3.3 0.0006951 3.3 0.0006952 0 0.00069512 0 0.00069522 3.3 0.00069514 3.3 0.00069524 0 0.00069516 0 0.00069526 3.3 0.00069518 3.3 0.0006952799999999999 0 0.0006952 0 0.0006952999999999999 3.3 0.0006952200000000001 3.3 0.00069532 0 0.0006952400000000001 0 0.00069534 3.3 0.0006952600000000001 3.3 0.00069536 0 0.00069528 0 0.00069538 3.3 0.0006953 3.3 0.0006954 0 0.00069532 0 0.00069542 3.3 0.00069534 3.3 0.00069544 0 0.00069536 0 0.00069546 3.3 0.00069538 3.3 0.00069548 0 0.0006954 0 0.0006954999999999999 3.3 0.0006954200000000001 3.3 0.00069552 0 0.0006954400000000001 0 0.00069554 3.3 0.0006954600000000001 3.3 0.00069556 0 0.0006954800000000001 0 0.00069558 3.3 0.0006955 3.3 0.0006956 0 0.00069552 0 0.00069562 3.3 0.00069554 3.3 0.00069564 0 0.00069556 0 0.00069566 3.3 0.00069558 3.3 0.00069568 0 0.0006956 0 0.0006956999999999999 3.3 0.00069562 3.3 0.0006957199999999999 0 0.0006956400000000001 0 0.00069574 3.3 0.0006956600000000001 3.3 0.00069576 0 0.0006956800000000001 0 0.00069578 3.3 0.0006957 3.3 0.0006958 0 0.00069572 0 0.00069582 3.3 0.00069574 3.3 0.00069584 0 0.00069576 0 0.00069586 3.3 0.00069578 3.3 0.00069588 0 0.0006958 0 0.0006959 3.3 0.00069582 3.3 0.0006959199999999999 0 0.0006958400000000001 0 0.00069594 3.3 0.0006958600000000001 3.3 0.00069596 0 0.0006958800000000001 0 0.00069598 3.3 0.0006959000000000001 3.3 0.000696 0 0.00069592 0 0.00069602 3.3 0.00069594 3.3 0.00069604 0 0.00069596 0 0.00069606 3.3 0.00069598 3.3 0.00069608 0 0.000696 0 0.0006961 3.3 0.00069602 3.3 0.0006961199999999999 0 0.0006960400000000001 0 0.00069614 3.3 0.0006960600000000001 3.3 0.00069616 0 0.0006960800000000001 0 0.00069618 3.3 0.0006961000000000001 3.3 0.0006962 0 0.00069612 0 0.00069622 3.3 0.00069614 3.3 0.00069624 0 0.00069616 0 0.00069626 3.3 0.00069618 3.3 0.00069628 0 0.0006962 0 0.0006963 3.3 0.00069622 3.3 0.00069632 0 0.00069624 0 0.0006963399999999999 3.3 0.0006962600000000001 3.3 0.00069636 0 0.0006962800000000001 0 0.00069638 3.3 0.0006963000000000001 3.3 0.0006964 0 0.0006963200000000001 0 0.00069642 3.3 0.00069634 3.3 0.00069644 0 0.00069636 0 0.00069646 3.3 0.00069638 3.3 0.00069648 0 0.0006964 0 0.0006965 3.3 0.00069642 3.3 0.00069652 0 0.00069644 0 0.0006965399999999999 3.3 0.0006964600000000001 3.3 0.00069656 0 0.0006964800000000001 0 0.00069658 3.3 0.0006965000000000001 3.3 0.0006966 0 0.0006965200000000001 0 0.00069662 3.3 0.00069654 3.3 0.00069664 0 0.00069656 0 0.00069666 3.3 0.00069658 3.3 0.00069668 0 0.0006966 0 0.0006967 3.3 0.00069662 3.3 0.00069672 0 0.00069664 0 0.00069674 3.3 0.00069666 3.3 0.0006967599999999999 0 0.0006966800000000001 0 0.00069678 3.3 0.0006967000000000001 3.3 0.0006968 0 0.0006967200000000001 0 0.00069682 3.3 0.0006967400000000001 3.3 0.00069684 0 0.00069676 0 0.00069686 3.3 0.00069678 3.3 0.00069688 0 0.0006968 0 0.0006969 3.3 0.00069682 3.3 0.00069692 0 0.00069684 0 0.00069694 3.3 0.00069686 3.3 0.0006969599999999999 0 0.0006968800000000001 0 0.00069698 3.3 0.0006969000000000001 3.3 0.000697 0 0.0006969200000000001 0 0.00069702 3.3 0.0006969400000000001 3.3 0.00069704 0 0.00069696 0 0.00069706 3.3 0.00069698 3.3 0.00069708 0 0.000697 0 0.0006971 3.3 0.00069702 3.3 0.00069712 0 0.00069704 0 0.00069714 3.3 0.00069706 3.3 0.0006971599999999999 0 0.00069708 0 0.0006971799999999999 3.3 0.0006971000000000001 3.3 0.0006972 0 0.0006971200000000001 0 0.00069722 3.3 0.0006971400000000001 3.3 0.00069724 0 0.00069716 0 0.00069726 3.3 0.00069718 3.3 0.00069728 0 0.0006972 0 0.0006973 3.3 0.00069722 3.3 0.00069732 0 0.00069724 0 0.00069734 3.3 0.00069726 3.3 0.00069736 0 0.00069728 0 0.0006973799999999999 3.3 0.0006973000000000001 3.3 0.0006974 0 0.0006973200000000001 0 0.00069742 3.3 0.0006973400000000001 3.3 0.00069744 0 0.0006973600000000001 0 0.00069746 3.3 0.00069738 3.3 0.00069748 0 0.0006974 0 0.0006975 3.3 0.00069742 3.3 0.00069752 0 0.00069744 0 0.00069754 3.3 0.00069746 3.3 0.00069756 0 0.00069748 0 0.0006975799999999999 3.3 0.0006975 3.3 0.0006975999999999999 0 0.0006975200000000001 0 0.00069762 3.3 0.0006975400000000001 3.3 0.00069764 0 0.0006975600000000001 0 0.00069766 3.3 0.00069758 3.3 0.00069768 0 0.0006976 0 0.0006977 3.3 0.00069762 3.3 0.00069772 0 0.00069764 0 0.00069774 3.3 0.00069766 3.3 0.00069776 0 0.00069768 0 0.00069778 3.3 0.0006977 3.3 0.0006977999999999999 0 0.0006977200000000001 0 0.00069782 3.3 0.0006977400000000001 3.3 0.00069784 0 0.0006977600000000001 0 0.00069786 3.3 0.0006977800000000001 3.3 0.00069788 0 0.0006978 0 0.0006979 3.3 0.00069782 3.3 0.00069792 0 0.00069784 0 0.00069794 3.3 0.00069786 3.3 0.00069796 0 0.00069788 0 0.00069798 3.3 0.0006979 3.3 0.0006979999999999999 0 0.00069792 0 0.0006980199999999999 3.3 0.0006979400000000001 3.3 0.00069804 0 0.0006979600000000001 0 0.00069806 3.3 0.0006979800000000001 3.3 0.00069808 0 0.000698 0 0.0006981 3.3 0.00069802 3.3 0.00069812 0 0.00069804 0 0.00069814 3.3 0.00069806 3.3 0.00069816 0 0.00069808 0 0.00069818 3.3 0.0006981 3.3 0.0006982 0 0.00069812 0 0.0006982199999999999 3.3 0.0006981400000000001 3.3 0.00069824 0 0.0006981600000000001 0 0.00069826 3.3 0.0006981800000000001 3.3 0.00069828 0 0.0006982000000000001 0 0.0006983 3.3 0.00069822 3.3 0.00069832 0 0.00069824 0 0.00069834 3.3 0.00069826 3.3 0.00069836 0 0.00069828 0 0.00069838 3.3 0.0006983 3.3 0.0006984 0 0.00069832 0 0.0006984199999999999 3.3 0.00069834 3.3 0.0006984399999999999 0 0.0006983600000000001 0 0.00069846 3.3 0.0006983800000000001 3.3 0.00069848 0 0.0006984000000000001 0 0.0006985 3.3 0.00069842 3.3 0.00069852 0 0.00069844 0 0.00069854 3.3 0.00069846 3.3 0.00069856 0 0.00069848 0 0.00069858 3.3 0.0006985 3.3 0.0006986 0 0.00069852 0 0.00069862 3.3 0.00069854 3.3 0.0006986399999999999 0 0.0006985600000000001 0 0.00069866 3.3 0.0006985800000000001 3.3 0.00069868 0 0.0006986000000000001 0 0.0006987 3.3 0.0006986200000000001 3.3 0.00069872 0 0.00069864 0 0.00069874 3.3 0.00069866 3.3 0.00069876 0 0.00069868 0 0.00069878 3.3 0.0006987 3.3 0.0006988 0 0.00069872 0 0.00069882 3.3 0.00069874 3.3 0.0006988399999999999 0 0.00069876 0 0.0006988599999999999 3.3 0.0006987800000000001 3.3 0.00069888 0 0.0006988000000000001 0 0.0006989 3.3 0.0006988200000000001 3.3 0.00069892 0 0.00069884 0 0.00069894 3.3 0.00069886 3.3 0.00069896 0 0.00069888 0 0.00069898 3.3 0.0006989 3.3 0.000699 0 0.00069892 0 0.00069902 3.3 0.00069894 3.3 0.00069904 0 0.00069896 0 0.0006990599999999999 3.3 0.0006989800000000001 3.3 0.00069908 0 0.0006990000000000001 0 0.0006991 3.3 0.0006990200000000001 3.3 0.00069912 0 0.0006990400000000001 0 0.00069914 3.3 0.00069906 3.3 0.00069916 0 0.00069908 0 0.00069918 3.3 0.0006991 3.3 0.0006992 0 0.00069912 0 0.00069922 3.3 0.00069914 3.3 0.00069924 0 0.00069916 0 0.0006992599999999999 3.3 0.00069918 3.3 0.0006992799999999999 0 0.0006992000000000001 0 0.0006993 3.3 0.0006992200000000001 3.3 0.00069932 0 0.0006992400000000001 0 0.00069934 3.3 0.00069926 3.3 0.00069936 0 0.00069928 0 0.00069938 3.3 0.0006993 3.3 0.0006994 0 0.00069932 0 0.00069942 3.3 0.00069934 3.3 0.00069944 0 0.00069936 0 0.00069946 3.3 0.00069938 3.3 0.0006994799999999999 0 0.0006994000000000001 0 0.0006995 3.3 0.0006994200000000001 3.3 0.00069952 0 0.0006994400000000001 0 0.00069954 3.3 0.0006994600000000001 3.3 0.00069956 0 0.00069948 0 0.00069958 3.3 0.0006995 3.3 0.0006996 0 0.00069952 0 0.00069962 3.3 0.00069954 3.3 0.00069964 0 0.00069956 0 0.00069966 3.3 0.00069958 3.3 0.0006996799999999999 0 0.0006996000000000001 0 0.0006997 3.3 0.0006996200000000001 3.3 0.00069972 0 0.0006996400000000001 0 0.00069974 3.3 0.0006996600000000001 3.3 0.00069976 0 0.00069968 0 0.00069978 3.3 0.0006997 3.3 0.0006998 0 0.00069972 0 0.00069982 3.3 0.00069974 3.3 0.00069984 0 0.00069976 0 0.00069986 3.3 0.00069978 3.3 0.00069988 0 0.0006998 0 0.0006998999999999999 3.3 0.0006998200000000001 3.3 0.00069992 0 0.0006998400000000001 0 0.00069994 3.3 0.0006998600000000001 3.3 0.00069996 0 0.0006998800000000001 0 0.00069998 3.3 0.0006999 3.3 0.0007 0 0.00069992 0 0.00070002 3.3 0.00069994 3.3 0.00070004 0 0.00069996 0 0.00070006 3.3 0.00069998 3.3 0.00070008 0 0.0007 0 0.0007000999999999999 3.3 0.0007000200000000001 3.3 0.00070012 0 0.0007000400000000001 0 0.00070014 3.3 0.0007000600000000001 3.3 0.00070016 0 0.0007000800000000001 0 0.00070018 3.3 0.0007001 3.3 0.0007002 0 0.00070012 0 0.00070022 3.3 0.00070014 3.3 0.00070024 0 0.00070016 0 0.00070026 3.3 0.00070018 3.3 0.00070028 0 0.0007002 0 0.0007003 3.3 0.00070022 3.3 0.0007003199999999999 0 0.0007002400000000001 0 0.00070034 3.3 0.0007002600000000001 3.3 0.00070036 0 0.0007002800000000001 0 0.00070038 3.3 0.0007003000000000001 3.3 0.0007004 0 0.00070032 0 0.00070042 3.3 0.00070034 3.3 0.00070044 0 0.00070036 0 0.00070046 3.3 0.00070038 3.3 0.00070048 0 0.0007004 0 0.0007005 3.3 0.00070042 3.3 0.0007005199999999999 0 0.0007004400000000001 0 0.00070054 3.3 0.0007004600000000001 3.3 0.00070056 0 0.0007004800000000001 0 0.00070058 3.3 0.0007005000000000001 3.3 0.0007006 0 0.00070052 0 0.00070062 3.3 0.00070054 3.3 0.00070064 0 0.00070056 0 0.00070066 3.3 0.00070058 3.3 0.00070068 0 0.0007006 0 0.0007007 3.3 0.00070062 3.3 0.0007007199999999999 0 0.00070064 0 0.0007007399999999999 3.3 0.0007006600000000001 3.3 0.00070076 0 0.0007006800000000001 0 0.00070078 3.3 0.0007007000000000001 3.3 0.0007008 0 0.00070072 0 0.00070082 3.3 0.00070074 3.3 0.00070084 0 0.00070076 0 0.00070086 3.3 0.00070078 3.3 0.00070088 0 0.0007008 0 0.0007009 3.3 0.00070082 3.3 0.00070092 0 0.00070084 0 0.0007009399999999999 3.3 0.0007008600000000001 3.3 0.00070096 0 0.0007008800000000001 0 0.00070098 3.3 0.0007009000000000001 3.3 0.000701 0 0.0007009200000000001 0 0.00070102 3.3 0.00070094 3.3 0.00070104 0 0.00070096 0 0.00070106 3.3 0.00070098 3.3 0.00070108 0 0.000701 0 0.0007011 3.3 0.00070102 3.3 0.00070112 0 0.00070104 0 0.0007011399999999999 3.3 0.00070106 3.3 0.0007011599999999999 0 0.0007010800000000001 0 0.00070118 3.3 0.0007011000000000001 3.3 0.0007012 0 0.0007011200000000001 0 0.00070122 3.3 0.00070114 3.3 0.00070124 0 0.00070116 0 0.00070126 3.3 0.00070118 3.3 0.00070128 0 0.0007012 0 0.0007013 3.3 0.00070122 3.3 0.00070132 0 0.00070124 0 0.00070134 3.3 0.00070126 3.3 0.0007013599999999999 0 0.0007012800000000001 0 0.00070138 3.3 0.0007013000000000001 3.3 0.0007014 0 0.0007013200000000001 0 0.00070142 3.3 0.0007013400000000001 3.3 0.00070144 0 0.00070136 0 0.00070146 3.3 0.00070138 3.3 0.00070148 0 0.0007014 0 0.0007015 3.3 0.00070142 3.3 0.00070152 0 0.00070144 0 0.00070154 3.3 0.00070146 3.3 0.0007015599999999999 0 0.00070148 0 0.0007015799999999999 3.3 0.0007015000000000001 3.3 0.0007016 0 0.0007015200000000001 0 0.00070162 3.3 0.0007015400000000001 3.3 0.00070164 0 0.00070156 0 0.00070166 3.3 0.00070158 3.3 0.00070168 0 0.0007016 0 0.0007017 3.3 0.00070162 3.3 0.00070172 0 0.00070164 0 0.00070174 3.3 0.00070166 3.3 0.00070176 0 0.00070168 0 0.0007017799999999999 3.3 0.0007017000000000001 3.3 0.0007018 0 0.0007017200000000001 0 0.00070182 3.3 0.0007017400000000001 3.3 0.00070184 0 0.0007017600000000001 0 0.00070186 3.3 0.00070178 3.3 0.00070188 0 0.0007018 0 0.0007019 3.3 0.00070182 3.3 0.00070192 0 0.00070184 0 0.00070194 3.3 0.00070186 3.3 0.00070196 0 0.00070188 0 0.0007019799999999999 3.3 0.0007019 3.3 0.0007019999999999999 0 0.0007019200000000001 0 0.00070202 3.3 0.0007019400000000001 3.3 0.00070204 0 0.0007019600000000001 0 0.00070206 3.3 0.00070198 3.3 0.00070208 0 0.000702 0 0.0007021 3.3 0.00070202 3.3 0.00070212 0 0.00070204 0 0.00070214 3.3 0.00070206 3.3 0.00070216 0 0.00070208 0 0.00070218 3.3 0.0007021 3.3 0.0007021999999999999 0 0.0007021200000000001 0 0.00070222 3.3 0.0007021400000000001 3.3 0.00070224 0 0.0007021600000000001 0 0.00070226 3.3 0.0007021800000000001 3.3 0.00070228 0 0.0007022 0 0.0007023 3.3 0.00070222 3.3 0.00070232 0 0.00070224 0 0.00070234 3.3 0.00070226 3.3 0.00070236 0 0.00070228 0 0.00070238 3.3 0.0007023 3.3 0.0007023999999999999 0 0.00070232 0 0.0007024199999999999 3.3 0.0007023400000000001 3.3 0.00070244 0 0.0007023600000000001 0 0.00070246 3.3 0.0007023800000000001 3.3 0.00070248 0 0.0007024 0 0.0007025 3.3 0.00070242 3.3 0.00070252 0 0.00070244 0 0.00070254 3.3 0.00070246 3.3 0.00070256 0 0.00070248 0 0.00070258 3.3 0.0007025 3.3 0.0007026 0 0.00070252 0 0.0007026199999999999 3.3 0.0007025400000000001 3.3 0.00070264 0 0.0007025600000000001 0 0.00070266 3.3 0.0007025800000000001 3.3 0.00070268 0 0.0007026000000000001 0 0.0007027 3.3 0.00070262 3.3 0.00070272 0 0.00070264 0 0.00070274 3.3 0.00070266 3.3 0.00070276 0 0.00070268 0 0.00070278 3.3 0.0007027 3.3 0.0007028 0 0.00070272 0 0.0007028199999999999 3.3 0.00070274 3.3 0.0007028399999999999 0 0.0007027600000000001 0 0.00070286 3.3 0.0007027800000000001 3.3 0.00070288 0 0.0007028000000000001 0 0.0007029 3.3 0.00070282 3.3 0.00070292 0 0.00070284 0 0.00070294 3.3 0.00070286 3.3 0.00070296 0 0.00070288 0 0.00070298 3.3 0.0007029 3.3 0.000703 0 0.00070292 0 0.00070302 3.3 0.00070294 3.3 0.0007030399999999999 0 0.0007029600000000001 0 0.00070306 3.3 0.0007029800000000001 3.3 0.00070308 0 0.0007030000000000001 0 0.0007031 3.3 0.0007030200000000001 3.3 0.00070312 0 0.00070304 0 0.00070314 3.3 0.00070306 3.3 0.00070316 0 0.00070308 0 0.00070318 3.3 0.0007031 3.3 0.0007032 0 0.00070312 0 0.00070322 3.3 0.00070314 3.3 0.0007032399999999999 0 0.0007031600000000001 0 0.00070326 3.3 0.0007031800000000001 3.3 0.00070328 0 0.0007032000000000001 0 0.0007033 3.3 0.0007032200000000001 3.3 0.00070332 0 0.00070324 0 0.00070334 3.3 0.00070326 3.3 0.00070336 0 0.00070328 0 0.00070338 3.3 0.0007033 3.3 0.0007034 0 0.00070332 0 0.00070342 3.3 0.00070334 3.3 0.00070344 0 0.00070336 0 0.0007034599999999999 3.3 0.0007033800000000001 3.3 0.00070348 0 0.0007034000000000001 0 0.0007035 3.3 0.0007034200000000001 3.3 0.00070352 0 0.0007034400000000001 0 0.00070354 3.3 0.00070346 3.3 0.00070356 0 0.00070348 0 0.00070358 3.3 0.0007035 3.3 0.0007036 0 0.00070352 0 0.00070362 3.3 0.00070354 3.3 0.00070364 0 0.00070356 0 0.0007036599999999999 3.3 0.0007035800000000001 3.3 0.00070368 0 0.0007036000000000001 0 0.0007037 3.3 0.0007036200000000001 3.3 0.00070372 0 0.0007036400000000001 0 0.00070374 3.3 0.00070366 3.3 0.00070376 0 0.00070368 0 0.00070378 3.3 0.0007037 3.3 0.0007038 0 0.00070372 0 0.00070382 3.3 0.00070374 3.3 0.00070384 0 0.00070376 0 0.0007038599999999999 3.3 0.00070378 3.3 0.0007038799999999999 0 0.0007038000000000001 0 0.0007039 3.3 0.0007038200000000001 3.3 0.00070392 0 0.0007038400000000001 0 0.00070394 3.3 0.00070386 3.3 0.00070396 0 0.00070388 0 0.00070398 3.3 0.0007039 3.3 0.000704 0 0.00070392 0 0.00070402 3.3 0.00070394 3.3 0.00070404 0 0.00070396 0 0.00070406 3.3 0.00070398 3.3 0.0007040799999999999 0 0.0007040000000000001 0 0.0007041 3.3 0.0007040200000000001 3.3 0.00070412 0 0.0007040400000000001 0 0.00070414 3.3 0.0007040600000000001 3.3 0.00070416 0 0.00070408 0 0.00070418 3.3 0.0007041 3.3 0.0007042 0 0.00070412 0 0.00070422 3.3 0.00070414 3.3 0.00070424 0 0.00070416 0 0.00070426 3.3 0.00070418 3.3 0.0007042799999999999 0 0.0007042 0 0.0007042999999999999 3.3 0.0007042200000000001 3.3 0.00070432 0 0.0007042400000000001 0 0.00070434 3.3 0.0007042600000000001 3.3 0.00070436 0 0.00070428 0 0.00070438 3.3 0.0007043 3.3 0.0007044 0 0.00070432 0 0.00070442 3.3 0.00070434 3.3 0.00070444 0 0.00070436 0 0.00070446 3.3 0.00070438 3.3 0.00070448 0 0.0007044 0 0.0007044999999999999 3.3 0.0007044200000000001 3.3 0.00070452 0 0.0007044400000000001 0 0.00070454 3.3 0.0007044600000000001 3.3 0.00070456 0 0.0007044800000000001 0 0.00070458 3.3 0.0007045 3.3 0.0007046 0 0.00070452 0 0.00070462 3.3 0.00070454 3.3 0.00070464 0 0.00070456 0 0.00070466 3.3 0.00070458 3.3 0.00070468 0 0.0007046 0 0.0007046999999999999 3.3 0.00070462 3.3 0.0007047199999999999 0 0.0007046400000000001 0 0.00070474 3.3 0.0007046600000000001 3.3 0.00070476 0 0.0007046800000000001 0 0.00070478 3.3 0.0007047 3.3 0.0007048 0 0.00070472 0 0.00070482 3.3 0.00070474 3.3 0.00070484 0 0.00070476 0 0.00070486 3.3 0.00070478 3.3 0.00070488 0 0.0007048 0 0.0007049 3.3 0.00070482 3.3 0.0007049199999999999 0 0.0007048400000000001 0 0.00070494 3.3 0.0007048600000000001 3.3 0.00070496 0 0.0007048800000000001 0 0.00070498 3.3 0.0007049000000000001 3.3 0.000705 0 0.00070492 0 0.00070502 3.3 0.00070494 3.3 0.00070504 0 0.00070496 0 0.00070506 3.3 0.00070498 3.3 0.00070508 0 0.000705 0 0.0007051 3.3 0.00070502 3.3 0.0007051199999999999 0 0.00070504 0 0.0007051399999999999 3.3 0.0007050600000000001 3.3 0.00070516 0 0.0007050800000000001 0 0.00070518 3.3 0.0007051000000000001 3.3 0.0007052 0 0.00070512 0 0.00070522 3.3 0.00070514 3.3 0.00070524 0 0.00070516 0 0.00070526 3.3 0.00070518 3.3 0.00070528 0 0.0007052 0 0.0007053 3.3 0.00070522 3.3 0.00070532 0 0.00070524 0 0.0007053399999999999 3.3 0.0007052600000000001 3.3 0.00070536 0 0.0007052800000000001 0 0.00070538 3.3 0.0007053000000000001 3.3 0.0007054 0 0.0007053200000000001 0 0.00070542 3.3 0.00070534 3.3 0.00070544 0 0.00070536 0 0.00070546 3.3 0.00070538 3.3 0.00070548 0 0.0007054 0 0.0007055 3.3 0.00070542 3.3 0.00070552 0 0.00070544 0 0.0007055399999999999 3.3 0.00070546 3.3 0.0007055599999999999 0 0.0007054800000000001 0 0.00070558 3.3 0.0007055000000000001 3.3 0.0007056 0 0.0007055200000000001 0 0.00070562 3.3 0.00070554 3.3 0.00070564 0 0.00070556 0 0.00070566 3.3 0.00070558 3.3 0.00070568 0 0.0007056 0 0.0007057 3.3 0.00070562 3.3 0.00070572 0 0.00070564 0 0.00070574 3.3 0.00070566 3.3 0.0007057599999999999 0 0.0007056800000000001 0 0.00070578 3.3 0.0007057000000000001 3.3 0.0007058 0 0.0007057200000000001 0 0.00070582 3.3 0.0007057400000000001 3.3 0.00070584 0 0.00070576 0 0.00070586 3.3 0.00070578 3.3 0.00070588 0 0.0007058 0 0.0007059 3.3 0.00070582 3.3 0.00070592 0 0.00070584 0 0.00070594 3.3 0.00070586 3.3 0.0007059599999999999 0 0.00070588 0 0.0007059799999999999 3.3 0.0007059000000000001 3.3 0.000706 0 0.0007059200000000001 0 0.00070602 3.3 0.0007059400000000001 3.3 0.00070604 0 0.00070596 0 0.00070606 3.3 0.00070598 3.3 0.00070608 0 0.000706 0 0.0007061 3.3 0.00070602 3.3 0.00070612 0 0.00070604 0 0.00070614 3.3 0.00070606 3.3 0.00070616 0 0.00070608 0 0.0007061799999999999 3.3 0.0007061000000000001 3.3 0.0007062 0 0.0007061200000000001 0 0.00070622 3.3 0.0007061400000000001 3.3 0.00070624 0 0.0007061600000000001 0 0.00070626 3.3 0.00070618 3.3 0.00070628 0 0.0007062 0 0.0007063 3.3 0.00070622 3.3 0.00070632 0 0.00070624 0 0.00070634 3.3 0.00070626 3.3 0.00070636 0 0.00070628 0 0.0007063799999999999 3.3 0.0007063 3.3 0.0007063999999999999 0 0.0007063200000000001 0 0.00070642 3.3 0.0007063400000000001 3.3 0.00070644 0 0.0007063600000000001 0 0.00070646 3.3 0.00070638 3.3 0.00070648 0 0.0007064 0 0.0007065 3.3 0.00070642 3.3 0.00070652 0 0.00070644 0 0.00070654 3.3 0.00070646 3.3 0.00070656 0 0.00070648 0 0.00070658 3.3 0.0007065 3.3 0.0007065999999999999 0 0.0007065200000000001 0 0.00070662 3.3 0.0007065400000000001 3.3 0.00070664 0 0.0007065600000000001 0 0.00070666 3.3 0.0007065800000000001 3.3 0.00070668 0 0.0007066 0 0.0007067 3.3 0.00070662 3.3 0.00070672 0 0.00070664 0 0.00070674 3.3 0.00070666 3.3 0.00070676 0 0.00070668 0 0.00070678 3.3 0.0007067 3.3 0.0007067999999999999 0 0.0007067200000000001 0 0.00070682 3.3 0.0007067400000000001 3.3 0.00070684 0 0.0007067600000000001 0 0.00070686 3.3 0.0007067800000000001 3.3 0.00070688 0 0.0007068 0 0.0007069 3.3 0.00070682 3.3 0.00070692 0 0.00070684 0 0.00070694 3.3 0.00070686 3.3 0.00070696 0 0.00070688 0 0.00070698 3.3 0.0007069 3.3 0.000707 0 0.00070692 0 0.0007070199999999999 3.3 0.0007069400000000001 3.3 0.00070704 0 0.0007069600000000001 0 0.00070706 3.3 0.0007069800000000001 3.3 0.00070708 0 0.0007070000000000001 0 0.0007071 3.3 0.00070702 3.3 0.00070712 0 0.00070704 0 0.00070714 3.3 0.00070706 3.3 0.00070716 0 0.00070708 0 0.00070718 3.3 0.0007071 3.3 0.0007072 0 0.00070712 0 0.0007072199999999999 3.3 0.0007071400000000001 3.3 0.00070724 0 0.0007071600000000001 0 0.00070726 3.3 0.0007071800000000001 3.3 0.00070728 0 0.0007072000000000001 0 0.0007073 3.3 0.00070722 3.3 0.00070732 0 0.00070724 0 0.00070734 3.3 0.00070726 3.3 0.00070736 0 0.00070728 0 0.00070738 3.3 0.0007073 3.3 0.0007074 0 0.00070732 0 0.0007074199999999999 3.3 0.00070734 3.3 0.0007074399999999999 0 0.0007073600000000001 0 0.00070746 3.3 0.0007073800000000001 3.3 0.00070748 0 0.0007074000000000001 0 0.0007075 3.3 0.00070742 3.3 0.00070752 0 0.00070744 0 0.00070754 3.3 0.00070746 3.3 0.00070756 0 0.00070748 0 0.00070758 3.3 0.0007075 3.3 0.0007076 0 0.00070752 0 0.00070762 3.3 0.00070754 3.3 0.0007076399999999999 0 0.0007075600000000001 0 0.00070766 3.3 0.0007075800000000001 3.3 0.00070768 0 0.0007076000000000001 0 0.0007077 3.3 0.0007076200000000001 3.3 0.00070772 0 0.00070764 0 0.00070774 3.3 0.00070766 3.3 0.00070776 0 0.00070768 0 0.00070778 3.3 0.0007077 3.3 0.0007078 0 0.00070772 0 0.00070782 3.3 0.00070774 3.3 0.0007078399999999999 0 0.00070776 0 0.0007078599999999999 3.3 0.0007077800000000001 3.3 0.00070788 0 0.0007078000000000001 0 0.0007079 3.3 0.0007078200000000001 3.3 0.00070792 0 0.00070784 0 0.00070794 3.3 0.00070786 3.3 0.00070796 0 0.00070788 0 0.00070798 3.3 0.0007079 3.3 0.000708 0 0.00070792 0 0.00070802 3.3 0.00070794 3.3 0.00070804 0 0.00070796 0 0.0007080599999999999 3.3 0.0007079800000000001 3.3 0.00070808 0 0.0007080000000000001 0 0.0007081 3.3 0.0007080200000000001 3.3 0.00070812 0 0.0007080400000000001 0 0.00070814 3.3 0.00070806 3.3 0.00070816 0 0.00070808 0 0.00070818 3.3 0.0007081 3.3 0.0007082 0 0.00070812 0 0.00070822 3.3 0.00070814 3.3 0.00070824 0 0.00070816 0 0.0007082599999999999 3.3 0.00070818 3.3 0.0007082799999999999 0 0.0007082000000000001 0 0.0007083 3.3 0.0007082200000000001 3.3 0.00070832 0 0.0007082400000000001 0 0.00070834 3.3 0.00070826 3.3 0.00070836 0 0.00070828 0 0.00070838 3.3 0.0007083 3.3 0.0007084 0 0.00070832 0 0.00070842 3.3 0.00070834 3.3 0.00070844 0 0.00070836 0 0.00070846 3.3 0.00070838 3.3 0.0007084799999999999 0 0.0007084000000000001 0 0.0007085 3.3 0.0007084200000000001 3.3 0.00070852 0 0.0007084400000000001 0 0.00070854 3.3 0.0007084600000000001 3.3 0.00070856 0 0.00070848 0 0.00070858 3.3 0.0007085 3.3 0.0007086 0 0.00070852 0 0.00070862 3.3 0.00070854 3.3 0.00070864 0 0.00070856 0 0.00070866 3.3 0.00070858 3.3 0.0007086799999999999 0 0.0007086 0 0.0007086999999999999 3.3 0.0007086200000000001 3.3 0.00070872 0 0.0007086400000000001 0 0.00070874 3.3 0.0007086600000000001 3.3 0.00070876 0 0.00070868 0 0.00070878 3.3 0.0007087 3.3 0.0007088 0 0.00070872 0 0.00070882 3.3 0.00070874 3.3 0.00070884 0 0.00070876 0 0.00070886 3.3 0.00070878 3.3 0.00070888 0 0.0007088 0 0.0007088999999999999 3.3 0.0007088200000000001 3.3 0.00070892 0 0.0007088400000000001 0 0.00070894 3.3 0.0007088600000000001 3.3 0.00070896 0 0.0007088800000000001 0 0.00070898 3.3 0.0007089 3.3 0.000709 0 0.00070892 0 0.00070902 3.3 0.00070894 3.3 0.00070904 0 0.00070896 0 0.00070906 3.3 0.00070898 3.3 0.00070908 0 0.000709 0 0.0007090999999999999 3.3 0.00070902 3.3 0.0007091199999999999 0 0.0007090400000000001 0 0.00070914 3.3 0.0007090600000000001 3.3 0.00070916 0 0.0007090800000000001 0 0.00070918 3.3 0.0007091 3.3 0.0007092 0 0.00070912 0 0.00070922 3.3 0.00070914 3.3 0.00070924 0 0.00070916 0 0.00070926 3.3 0.00070918 3.3 0.00070928 0 0.0007092 0 0.0007093 3.3 0.00070922 3.3 0.0007093199999999999 0 0.0007092400000000001 0 0.00070934 3.3 0.0007092600000000001 3.3 0.00070936 0 0.0007092800000000001 0 0.00070938 3.3 0.0007093000000000001 3.3 0.0007094 0 0.00070932 0 0.00070942 3.3 0.00070934 3.3 0.00070944 0 0.00070936 0 0.00070946 3.3 0.00070938 3.3 0.00070948 0 0.0007094 0 0.0007095 3.3 0.00070942 3.3 0.0007095199999999999 0 0.00070944 0 0.0007095399999999999 3.3 0.0007094600000000001 3.3 0.00070956 0 0.0007094800000000001 0 0.00070958 3.3 0.0007095000000000001 3.3 0.0007096 0 0.00070952 0 0.00070962 3.3 0.00070954 3.3 0.00070964 0 0.00070956 0 0.00070966 3.3 0.00070958 3.3 0.00070968 0 0.0007096 0 0.0007097 3.3 0.00070962 3.3 0.00070972 0 0.00070964 0 0.0007097399999999999 3.3 0.0007096600000000001 3.3 0.00070976 0 0.0007096800000000001 0 0.00070978 3.3 0.0007097000000000001 3.3 0.0007098 0 0.0007097200000000001 0 0.00070982 3.3 0.00070974 3.3 0.00070984 0 0.00070976 0 0.00070986 3.3 0.00070978 3.3 0.00070988 0 0.0007098 0 0.0007099 3.3 0.00070982 3.3 0.00070992 0 0.00070984 0 0.0007099399999999999 3.3 0.0007098600000000001 3.3 0.00070996 0 0.0007098800000000001 0 0.00070998 3.3 0.0007099000000000001 3.3 0.00071 0 0.0007099200000000001 0 0.00071002 3.3 0.00070994 3.3 0.00071004 0 0.00070996 0 0.00071006 3.3 0.00070998 3.3 0.00071008 0 0.00071 0 0.0007101 3.3 0.00071002 3.3 0.00071012 0 0.00071004 0 0.00071014 3.3 0.00071006 3.3 0.0007101599999999999 0 0.0007100800000000001 0 0.00071018 3.3 0.0007101000000000001 3.3 0.0007102 0 0.0007101200000000001 0 0.00071022 3.3 0.0007101400000000001 3.3 0.00071024 0 0.00071016 0 0.00071026 3.3 0.00071018 3.3 0.00071028 0 0.0007102 0 0.0007103 3.3 0.00071022 3.3 0.00071032 0 0.00071024 0 0.00071034 3.3 0.00071026 3.3 0.0007103599999999999 0 0.0007102800000000001 0 0.00071038 3.3 0.0007103000000000001 3.3 0.0007104 0 0.0007103200000000001 0 0.00071042 3.3 0.0007103400000000001 3.3 0.00071044 0 0.00071036 0 0.00071046 3.3 0.00071038 3.3 0.00071048 0 0.0007104 0 0.0007105 3.3 0.00071042 3.3 0.00071052 0 0.00071044 0 0.00071054 3.3 0.00071046 3.3 0.00071056 0 0.00071048 0 0.0007105799999999999 3.3 0.0007105000000000001 3.3 0.0007106 0 0.0007105200000000001 0 0.00071062 3.3 0.0007105400000000001 3.3 0.00071064 0 0.0007105600000000001 0 0.00071066 3.3 0.00071058 3.3 0.00071068 0 0.0007106 0 0.0007107 3.3 0.00071062 3.3 0.00071072 0 0.00071064 0 0.00071074 3.3 0.00071066 3.3 0.00071076 0 0.00071068 0 0.0007107799999999999 3.3 0.0007107000000000001 3.3 0.0007108 0 0.0007107200000000001 0 0.00071082 3.3 0.0007107400000000001 3.3 0.00071084 0 0.0007107600000000001 0 0.00071086 3.3 0.00071078 3.3 0.00071088 0 0.0007108 0 0.0007109 3.3 0.00071082 3.3 0.00071092 0 0.00071084 0 0.00071094 3.3 0.00071086 3.3 0.00071096 0 0.00071088 0 0.0007109799999999999 3.3 0.0007109 3.3 0.0007109999999999999 0 0.0007109200000000001 0 0.00071102 3.3 0.0007109400000000001 3.3 0.00071104 0 0.0007109600000000001 0 0.00071106 3.3 0.00071098 3.3 0.00071108 0 0.000711 0 0.0007111 3.3 0.00071102 3.3 0.00071112 0 0.00071104 0 0.00071114 3.3 0.00071106 3.3 0.00071116 0 0.00071108 0 0.00071118 3.3 0.0007111 3.3 0.0007111999999999999 0 0.0007111200000000001 0 0.00071122 3.3 0.0007111400000000001 3.3 0.00071124 0 0.0007111600000000001 0 0.00071126 3.3 0.0007111800000000001 3.3 0.00071128 0 0.0007112 0 0.0007113 3.3 0.00071122 3.3 0.00071132 0 0.00071124 0 0.00071134 3.3 0.00071126 3.3 0.00071136 0 0.00071128 0 0.00071138 3.3 0.0007113 3.3 0.0007113999999999999 0 0.00071132 0 0.0007114199999999999 3.3 0.0007113400000000001 3.3 0.00071144 0 0.0007113600000000001 0 0.00071146 3.3 0.0007113800000000001 3.3 0.00071148 0 0.0007114 0 0.0007115 3.3 0.00071142 3.3 0.00071152 0 0.00071144 0 0.00071154 3.3 0.00071146 3.3 0.00071156 0 0.00071148 0 0.00071158 3.3 0.0007115 3.3 0.0007116 0 0.00071152 0 0.0007116199999999999 3.3 0.0007115400000000001 3.3 0.00071164 0 0.0007115600000000001 0 0.00071166 3.3 0.0007115800000000001 3.3 0.00071168 0 0.0007116000000000001 0 0.0007117 3.3 0.00071162 3.3 0.00071172 0 0.00071164 0 0.00071174 3.3 0.00071166 3.3 0.00071176 0 0.00071168 0 0.00071178 3.3 0.0007117 3.3 0.0007118 0 0.00071172 0 0.0007118199999999999 3.3 0.00071174 3.3 0.0007118399999999999 0 0.0007117600000000001 0 0.00071186 3.3 0.0007117800000000001 3.3 0.00071188 0 0.0007118000000000001 0 0.0007119 3.3 0.00071182 3.3 0.00071192 0 0.00071184 0 0.00071194 3.3 0.00071186 3.3 0.00071196 0 0.00071188 0 0.00071198 3.3 0.0007119 3.3 0.000712 0 0.00071192 0 0.00071202 3.3 0.00071194 3.3 0.0007120399999999999 0 0.0007119600000000001 0 0.00071206 3.3 0.0007119800000000001 3.3 0.00071208 0 0.0007120000000000001 0 0.0007121 3.3 0.0007120200000000001 3.3 0.00071212 0 0.00071204 0 0.00071214 3.3 0.00071206 3.3 0.00071216 0 0.00071208 0 0.00071218 3.3 0.0007121 3.3 0.0007122 0 0.00071212 0 0.00071222 3.3 0.00071214 3.3 0.0007122399999999999 0 0.00071216 0 0.0007122599999999999 3.3 0.0007121800000000001 3.3 0.00071228 0 0.0007122000000000001 0 0.0007123 3.3 0.0007122200000000001 3.3 0.00071232 0 0.00071224 0 0.00071234 3.3 0.00071226 3.3 0.00071236 0 0.00071228 0 0.00071238 3.3 0.0007123 3.3 0.0007124 0 0.00071232 0 0.00071242 3.3 0.00071234 3.3 0.00071244 0 0.00071236 0 0.0007124599999999999 3.3 0.0007123800000000001 3.3 0.00071248 0 0.0007124000000000001 0 0.0007125 3.3 0.0007124200000000001 3.3 0.00071252 0 0.0007124400000000001 0 0.00071254 3.3 0.00071246 3.3 0.00071256 0 0.00071248 0 0.00071258 3.3 0.0007125 3.3 0.0007126 0 0.00071252 0 0.00071262 3.3 0.00071254 3.3 0.00071264 0 0.00071256 0 0.0007126599999999999 3.3 0.00071258 3.3 0.0007126799999999999 0 0.0007126000000000001 0 0.0007127 3.3 0.0007126200000000001 3.3 0.00071272 0 0.0007126400000000001 0 0.00071274 3.3 0.00071266 3.3 0.00071276 0 0.00071268 0 0.00071278 3.3 0.0007127 3.3 0.0007128 0 0.00071272 0 0.00071282 3.3 0.00071274 3.3 0.00071284 0 0.00071276 0 0.00071286 3.3 0.00071278 3.3 0.0007128799999999999 0 0.0007128000000000001 0 0.0007129 3.3 0.0007128200000000001 3.3 0.00071292 0 0.0007128400000000001 0 0.00071294 3.3 0.0007128600000000001 3.3 0.00071296 0 0.00071288 0 0.00071298 3.3 0.0007129 3.3 0.000713 0 0.00071292 0 0.00071302 3.3 0.00071294 3.3 0.00071304 0 0.00071296 0 0.00071306 3.3 0.00071298 3.3 0.0007130799999999999 0 0.000713 0 0.0007130999999999999 3.3 0.0007130200000000001 3.3 0.00071312 0 0.0007130400000000001 0 0.00071314 3.3 0.0007130600000000001 3.3 0.00071316 0 0.00071308 0 0.00071318 3.3 0.0007131 3.3 0.0007132 0 0.00071312 0 0.00071322 3.3 0.00071314 3.3 0.00071324 0 0.00071316 0 0.00071326 3.3 0.00071318 3.3 0.00071328 0 0.0007132 0 0.0007132999999999999 3.3 0.0007132200000000001 3.3 0.00071332 0 0.0007132400000000001 0 0.00071334 3.3 0.0007132600000000001 3.3 0.00071336 0 0.0007132800000000001 0 0.00071338 3.3 0.0007133 3.3 0.0007134 0 0.00071332 0 0.00071342 3.3 0.00071334 3.3 0.00071344 0 0.00071336 0 0.00071346 3.3 0.00071338 3.3 0.00071348 0 0.0007134 0 0.0007134999999999999 3.3 0.0007134200000000001 3.3 0.00071352 0 0.0007134400000000001 0 0.00071354 3.3 0.0007134600000000001 3.3 0.00071356 0 0.0007134800000000001 0 0.00071358 3.3 0.0007135 3.3 0.0007136 0 0.00071352 0 0.00071362 3.3 0.00071354 3.3 0.00071364 0 0.00071356 0 0.00071366 3.3 0.00071358 3.3 0.00071368 0 0.0007136 0 0.0007137 3.3 0.00071362 3.3 0.0007137199999999999 0 0.0007136400000000001 0 0.00071374 3.3 0.0007136600000000001 3.3 0.00071376 0 0.0007136800000000001 0 0.00071378 3.3 0.0007137000000000001 3.3 0.0007138 0 0.00071372 0 0.00071382 3.3 0.00071374 3.3 0.00071384 0 0.00071376 0 0.00071386 3.3 0.00071378 3.3 0.00071388 0 0.0007138 0 0.0007139 3.3 0.00071382 3.3 0.0007139199999999999 0 0.0007138400000000001 0 0.00071394 3.3 0.0007138600000000001 3.3 0.00071396 0 0.0007138800000000001 0 0.00071398 3.3 0.0007139000000000001 3.3 0.000714 0 0.00071392 0 0.00071402 3.3 0.00071394 3.3 0.00071404 0 0.00071396 0 0.00071406 3.3 0.00071398 3.3 0.00071408 0 0.000714 0 0.0007141 3.3 0.00071402 3.3 0.0007141199999999999 0 0.00071404 0 0.0007141399999999999 3.3 0.0007140600000000001 3.3 0.00071416 0 0.0007140800000000001 0 0.00071418 3.3 0.0007141000000000001 3.3 0.0007142 0 0.00071412 0 0.00071422 3.3 0.00071414 3.3 0.00071424 0 0.00071416 0 0.00071426 3.3 0.00071418 3.3 0.00071428 0 0.0007142 0 0.0007143 3.3 0.00071422 3.3 0.00071432 0 0.00071424 0 0.0007143399999999999 3.3 0.0007142600000000001 3.3 0.00071436 0 0.0007142800000000001 0 0.00071438 3.3 0.0007143000000000001 3.3 0.0007144 0 0.0007143200000000001 0 0.00071442 3.3 0.00071434 3.3 0.00071444 0 0.00071436 0 0.00071446 3.3 0.00071438 3.3 0.00071448 0 0.0007144 0 0.0007145 3.3 0.00071442 3.3 0.00071452 0 0.00071444 0 0.0007145399999999999 3.3 0.00071446 3.3 0.0007145599999999999 0 0.0007144800000000001 0 0.00071458 3.3 0.0007145000000000001 3.3 0.0007146 0 0.0007145200000000001 0 0.00071462 3.3 0.00071454 3.3 0.00071464 0 0.00071456 0 0.00071466 3.3 0.00071458 3.3 0.00071468 0 0.0007146 0 0.0007147 3.3 0.00071462 3.3 0.00071472 0 0.00071464 0 0.00071474 3.3 0.00071466 3.3 0.0007147599999999999 0 0.0007146800000000001 0 0.00071478 3.3 0.0007147000000000001 3.3 0.0007148 0 0.0007147200000000001 0 0.00071482 3.3 0.0007147400000000001 3.3 0.00071484 0 0.00071476 0 0.00071486 3.3 0.00071478 3.3 0.00071488 0 0.0007148 0 0.0007149 3.3 0.00071482 3.3 0.00071492 0 0.00071484 0 0.00071494 3.3 0.00071486 3.3 0.0007149599999999999 0 0.00071488 0 0.0007149799999999999 3.3 0.0007149000000000001 3.3 0.000715 0 0.0007149200000000001 0 0.00071502 3.3 0.0007149400000000001 3.3 0.00071504 0 0.00071496 0 0.00071506 3.3 0.00071498 3.3 0.00071508 0 0.000715 0 0.0007151 3.3 0.00071502 3.3 0.00071512 0 0.00071504 0 0.00071514 3.3 0.00071506 3.3 0.00071516 0 0.00071508 0 0.0007151799999999999 3.3 0.0007151000000000001 3.3 0.0007152 0 0.0007151200000000001 0 0.00071522 3.3 0.0007151400000000001 3.3 0.00071524 0 0.0007151600000000001 0 0.00071526 3.3 0.00071518 3.3 0.00071528 0 0.0007152 0 0.0007153 3.3 0.00071522 3.3 0.00071532 0 0.00071524 0 0.00071534 3.3 0.00071526 3.3 0.00071536 0 0.00071528 0 0.0007153799999999999 3.3 0.0007153 3.3 0.0007153999999999999 0 0.0007153200000000001 0 0.00071542 3.3 0.0007153400000000001 3.3 0.00071544 0 0.0007153600000000001 0 0.00071546 3.3 0.00071538 3.3 0.00071548 0 0.0007154 0 0.0007155 3.3 0.00071542 3.3 0.00071552 0 0.00071544 0 0.00071554 3.3 0.00071546 3.3 0.00071556 0 0.00071548 0 0.00071558 3.3 0.0007155 3.3 0.0007155999999999999 0 0.0007155200000000001 0 0.00071562 3.3 0.0007155400000000001 3.3 0.00071564 0 0.0007155600000000001 0 0.00071566 3.3 0.0007155800000000001 3.3 0.00071568 0 0.0007156 0 0.0007157 3.3 0.00071562 3.3 0.00071572 0 0.00071564 0 0.00071574 3.3 0.00071566 3.3 0.00071576 0 0.00071568 0 0.00071578 3.3 0.0007157 3.3 0.0007157999999999999 0 0.00071572 0 0.0007158199999999999 3.3 0.0007157400000000001 3.3 0.00071584 0 0.0007157600000000001 0 0.00071586 3.3 0.0007157800000000001 3.3 0.00071588 0 0.0007158 0 0.0007159 3.3 0.00071582 3.3 0.00071592 0 0.00071584 0 0.00071594 3.3 0.00071586 3.3 0.00071596 0 0.00071588 0 0.00071598 3.3 0.0007159 3.3 0.000716 0 0.00071592 0 0.0007160199999999999 3.3 0.0007159400000000001 3.3 0.00071604 0 0.0007159600000000001 0 0.00071606 3.3 0.0007159800000000001 3.3 0.00071608 0 0.0007160000000000001 0 0.0007161 3.3 0.00071602 3.3 0.00071612 0 0.00071604 0 0.00071614 3.3 0.00071606 3.3 0.00071616 0 0.00071608 0 0.00071618 3.3 0.0007161 3.3 0.0007162 0 0.00071612 0 0.0007162199999999999 3.3 0.00071614 3.3 0.0007162399999999999 0 0.0007161600000000001 0 0.00071626 3.3 0.0007161800000000001 3.3 0.00071628 0 0.0007162000000000001 0 0.0007163 3.3 0.00071622 3.3 0.00071632 0 0.00071624 0 0.00071634 3.3 0.00071626 3.3 0.00071636 0 0.00071628 0 0.00071638 3.3 0.0007163 3.3 0.0007164 0 0.00071632 0 0.00071642 3.3 0.00071634 3.3 0.0007164399999999999 0 0.0007163600000000001 0 0.00071646 3.3 0.0007163800000000001 3.3 0.00071648 0 0.0007164000000000001 0 0.0007165 3.3 0.0007164200000000001 3.3 0.00071652 0 0.00071644 0 0.00071654 3.3 0.00071646 3.3 0.00071656 0 0.00071648 0 0.00071658 3.3 0.0007165 3.3 0.0007166 0 0.00071652 0 0.00071662 3.3 0.00071654 3.3 0.0007166399999999999 0 0.00071656 0 0.0007166599999999999 3.3 0.0007165800000000001 3.3 0.00071668 0 0.0007166000000000001 0 0.0007167 3.3 0.0007166200000000001 3.3 0.00071672 0 0.00071664 0 0.00071674 3.3 0.00071666 3.3 0.00071676 0 0.00071668 0 0.00071678 3.3 0.0007167 3.3 0.0007168 0 0.00071672 0 0.00071682 3.3 0.00071674 3.3 0.00071684 0 0.00071676 0 0.0007168599999999999 3.3 0.0007167800000000001 3.3 0.00071688 0 0.0007168000000000001 0 0.0007169 3.3 0.0007168200000000001 3.3 0.00071692 0 0.0007168400000000001 0 0.00071694 3.3 0.00071686 3.3 0.00071696 0 0.00071688 0 0.00071698 3.3 0.0007169 3.3 0.000717 0 0.00071692 0 0.00071702 3.3 0.00071694 3.3 0.00071704 0 0.00071696 0 0.0007170599999999999 3.3 0.0007169800000000001 3.3 0.00071708 0 0.0007170000000000001 0 0.0007171 3.3 0.0007170200000000001 3.3 0.00071712 0 0.0007170400000000001 0 0.00071714 3.3 0.00071706 3.3 0.00071716 0 0.00071708 0 0.00071718 3.3 0.0007171 3.3 0.0007172 0 0.00071712 0 0.00071722 3.3 0.00071714 3.3 0.00071724 0 0.00071716 0 0.00071726 3.3 0.00071718 3.3 0.0007172799999999999 0 0.0007172000000000001 0 0.0007173 3.3 0.0007172200000000001 3.3 0.00071732 0 0.0007172400000000001 0 0.00071734 3.3 0.0007172600000000001 3.3 0.00071736 0 0.00071728 0 0.00071738 3.3 0.0007173 3.3 0.0007174 0 0.00071732 0 0.00071742 3.3 0.00071734 3.3 0.00071744 0 0.00071736 0 0.00071746 3.3 0.00071738 3.3 0.0007174799999999999 0 0.0007174000000000001 0 0.0007175 3.3 0.0007174200000000001 3.3 0.00071752 0 0.0007174400000000001 0 0.00071754 3.3 0.0007174600000000001 3.3 0.00071756 0 0.00071748 0 0.00071758 3.3 0.0007175 3.3 0.0007176 0 0.00071752 0 0.00071762 3.3 0.00071754 3.3 0.00071764 0 0.00071756 0 0.00071766 3.3 0.00071758 3.3 0.0007176799999999999 0 0.0007176 0 0.0007176999999999999 3.3 0.0007176200000000001 3.3 0.00071772 0 0.0007176400000000001 0 0.00071774 3.3 0.0007176600000000001 3.3 0.00071776 0 0.00071768 0 0.00071778 3.3 0.0007177 3.3 0.0007178 0 0.00071772 0 0.00071782 3.3 0.00071774 3.3 0.00071784 0 0.00071776 0 0.00071786 3.3 0.00071778 3.3 0.00071788 0 0.0007178 0 0.0007178999999999999 3.3 0.0007178200000000001 3.3 0.00071792 0 0.0007178400000000001 0 0.00071794 3.3 0.0007178600000000001 3.3 0.00071796 0 0.0007178800000000001 0 0.00071798 3.3 0.0007179 3.3 0.000718 0 0.00071792 0 0.00071802 3.3 0.00071794 3.3 0.00071804 0 0.00071796 0 0.00071806 3.3 0.00071798 3.3 0.00071808 0 0.000718 0 0.0007180999999999999 3.3 0.00071802 3.3 0.0007181199999999999 0 0.0007180400000000001 0 0.00071814 3.3 0.0007180600000000001 3.3 0.00071816 0 0.0007180800000000001 0 0.00071818 3.3 0.0007181 3.3 0.0007182 0 0.00071812 0 0.00071822 3.3 0.00071814 3.3 0.00071824 0 0.00071816 0 0.00071826 3.3 0.00071818 3.3 0.00071828 0 0.0007182 0 0.0007183 3.3 0.00071822 3.3 0.0007183199999999999 0 0.0007182400000000001 0 0.00071834 3.3 0.0007182600000000001 3.3 0.00071836 0 0.0007182800000000001 0 0.00071838 3.3 0.0007183000000000001 3.3 0.0007184 0 0.00071832 0 0.00071842 3.3 0.00071834 3.3 0.00071844 0 0.00071836 0 0.00071846 3.3 0.00071838 3.3 0.00071848 0 0.0007184 0 0.0007185 3.3 0.00071842 3.3 0.0007185199999999999 0 0.00071844 0 0.0007185399999999999 3.3 0.0007184600000000001 3.3 0.00071856 0 0.0007184800000000001 0 0.00071858 3.3 0.0007185000000000001 3.3 0.0007186 0 0.00071852 0 0.00071862 3.3 0.00071854 3.3 0.00071864 0 0.00071856 0 0.00071866 3.3 0.00071858 3.3 0.00071868 0 0.0007186 0 0.0007187 3.3 0.00071862 3.3 0.00071872 0 0.00071864 0 0.0007187399999999999 3.3 0.0007186600000000001 3.3 0.00071876 0 0.0007186800000000001 0 0.00071878 3.3 0.0007187000000000001 3.3 0.0007188 0 0.0007187200000000001 0 0.00071882 3.3 0.00071874 3.3 0.00071884 0 0.00071876 0 0.00071886 3.3 0.00071878 3.3 0.00071888 0 0.0007188 0 0.0007189 3.3 0.00071882 3.3 0.00071892 0 0.00071884 0 0.0007189399999999999 3.3 0.00071886 3.3 0.0007189599999999999 0 0.0007188800000000001 0 0.00071898 3.3 0.0007189000000000001 3.3 0.000719 0 0.0007189200000000001 0 0.00071902 3.3 0.00071894 3.3 0.00071904 0 0.00071896 0 0.00071906 3.3 0.00071898 3.3 0.00071908 0 0.000719 0 0.0007191 3.3 0.00071902 3.3 0.00071912 0 0.00071904 0 0.00071914 3.3 0.00071906 3.3 0.0007191599999999999 0 0.0007190800000000001 0 0.00071918 3.3 0.0007191000000000001 3.3 0.0007192 0 0.0007191200000000001 0 0.00071922 3.3 0.0007191400000000001 3.3 0.00071924 0 0.00071916 0 0.00071926 3.3 0.00071918 3.3 0.00071928 0 0.0007192 0 0.0007193 3.3 0.00071922 3.3 0.00071932 0 0.00071924 0 0.00071934 3.3 0.00071926 3.3 0.0007193599999999999 0 0.00071928 0 0.0007193799999999999 3.3 0.0007193000000000001 3.3 0.0007194 0 0.0007193200000000001 0 0.00071942 3.3 0.0007193400000000001 3.3 0.00071944 0 0.00071936 0 0.00071946 3.3 0.00071938 3.3 0.00071948 0 0.0007194 0 0.0007195 3.3 0.00071942 3.3 0.00071952 0 0.00071944 0 0.00071954 3.3 0.00071946 3.3 0.00071956 0 0.00071948 0 0.0007195799999999999 3.3 0.0007195000000000001 3.3 0.0007196 0 0.0007195200000000001 0 0.00071962 3.3 0.0007195400000000001 3.3 0.00071964 0 0.0007195600000000001 0 0.00071966 3.3 0.00071958 3.3 0.00071968 0 0.0007196 0 0.0007197 3.3 0.00071962 3.3 0.00071972 0 0.00071964 0 0.00071974 3.3 0.00071966 3.3 0.00071976 0 0.00071968 0 0.0007197799999999999 3.3 0.0007197 3.3 0.0007197999999999999 0 0.0007197200000000001 0 0.00071982 3.3 0.0007197400000000001 3.3 0.00071984 0 0.0007197600000000001 0 0.00071986 3.3 0.00071978 3.3 0.00071988 0 0.0007198 0 0.0007199 3.3 0.00071982 3.3 0.00071992 0 0.00071984 0 0.00071994 3.3 0.00071986 3.3 0.00071996 0 0.00071988 0 0.00071998 3.3 0.0007199 3.3 0.0007199999999999999 0 0.0007199200000000001 0 0.00072002 3.3 0.0007199400000000001 3.3 0.00072004 0 0.0007199600000000001 0 0.00072006 3.3 0.0007199800000000001 3.3 0.00072008 0 0.00072 0 0.0007201 3.3 0.00072002 3.3 0.00072012 0 0.00072004 0 0.00072014 3.3 0.00072006 3.3 0.00072016 0 0.00072008 0 0.00072018 3.3 0.0007201 3.3 0.0007201999999999999 0 0.00072012 0 0.0007202199999999999 3.3 0.0007201400000000001 3.3 0.00072024 0 0.0007201600000000001 0 0.00072026 3.3 0.0007201800000000001 3.3 0.00072028 0 0.0007202 0 0.0007203 3.3 0.00072022 3.3 0.00072032 0 0.00072024 0 0.00072034 3.3 0.00072026 3.3 0.00072036 0 0.00072028 0 0.00072038 3.3 0.0007203 3.3 0.0007204 0 0.00072032 0 0.0007204199999999999 3.3 0.0007203400000000001 3.3 0.00072044 0 0.0007203600000000001 0 0.00072046 3.3 0.0007203800000000001 3.3 0.00072048 0 0.0007204000000000001 0 0.0007205 3.3 0.00072042 3.3 0.00072052 0 0.00072044 0 0.00072054 3.3 0.00072046 3.3 0.00072056 0 0.00072048 0 0.00072058 3.3 0.0007205 3.3 0.0007206 0 0.00072052 0 0.0007206199999999999 3.3 0.0007205400000000001 3.3 0.00072064 0 0.0007205600000000001 0 0.00072066 3.3 0.0007205800000000001 3.3 0.00072068 0 0.0007206000000000001 0 0.0007207 3.3 0.00072062 3.3 0.00072072 0 0.00072064 0 0.00072074 3.3 0.00072066 3.3 0.00072076 0 0.00072068 0 0.00072078 3.3 0.0007207 3.3 0.0007208 0 0.00072072 0 0.00072082 3.3 0.00072074 3.3 0.0007208399999999999 0 0.0007207600000000001 0 0.00072086 3.3 0.0007207800000000001 3.3 0.00072088 0 0.0007208000000000001 0 0.0007209 3.3 0.0007208200000000001 3.3 0.00072092 0 0.00072084 0 0.00072094 3.3 0.00072086 3.3 0.00072096 0 0.00072088 0 0.00072098 3.3 0.0007209 3.3 0.000721 0 0.00072092 0 0.00072102 3.3 0.00072094 3.3 0.0007210399999999999 0 0.0007209600000000001 0 0.00072106 3.3 0.0007209800000000001 3.3 0.00072108 0 0.0007210000000000001 0 0.0007211 3.3 0.0007210200000000001 3.3 0.00072112 0 0.00072104 0 0.00072114 3.3 0.00072106 3.3 0.00072116 0 0.00072108 0 0.00072118 3.3 0.0007211 3.3 0.0007212 0 0.00072112 0 0.00072122 3.3 0.00072114 3.3 0.0007212399999999999 0 0.00072116 0 0.0007212599999999999 3.3 0.0007211800000000001 3.3 0.00072128 0 0.0007212000000000001 0 0.0007213 3.3 0.0007212200000000001 3.3 0.00072132 0 0.00072124 0 0.00072134 3.3 0.00072126 3.3 0.00072136 0 0.00072128 0 0.00072138 3.3 0.0007213 3.3 0.0007214 0 0.00072132 0 0.00072142 3.3 0.00072134 3.3 0.00072144 0 0.00072136 0 0.0007214599999999999 3.3 0.0007213800000000001 3.3 0.00072148 0 0.0007214000000000001 0 0.0007215 3.3 0.0007214200000000001 3.3 0.00072152 0 0.0007214400000000001 0 0.00072154 3.3 0.00072146 3.3 0.00072156 0 0.00072148 0 0.00072158 3.3 0.0007215 3.3 0.0007216 0 0.00072152 0 0.00072162 3.3 0.00072154 3.3 0.00072164 0 0.00072156 0 0.0007216599999999999 3.3 0.00072158 3.3 0.0007216799999999999 0 0.0007216000000000001 0 0.0007217 3.3 0.0007216200000000001 3.3 0.00072172 0 0.0007216400000000001 0 0.00072174 3.3 0.00072166 3.3 0.00072176 0 0.00072168 0 0.00072178 3.3 0.0007217 3.3 0.0007218 0 0.00072172 0 0.00072182 3.3 0.00072174 3.3 0.00072184 0 0.00072176 0 0.00072186 3.3 0.00072178 3.3 0.0007218799999999999 0 0.0007218000000000001 0 0.0007219 3.3 0.0007218200000000001 3.3 0.00072192 0 0.0007218400000000001 0 0.00072194 3.3 0.0007218600000000001 3.3 0.00072196 0 0.00072188 0 0.00072198 3.3 0.0007219 3.3 0.000722 0 0.00072192 0 0.00072202 3.3 0.00072194 3.3 0.00072204 0 0.00072196 0 0.00072206 3.3 0.00072198 3.3 0.0007220799999999999 0 0.000722 0 0.0007220999999999999 3.3 0.0007220200000000001 3.3 0.00072212 0 0.0007220400000000001 0 0.00072214 3.3 0.0007220600000000001 3.3 0.00072216 0 0.00072208 0 0.00072218 3.3 0.0007221 3.3 0.0007222 0 0.00072212 0 0.00072222 3.3 0.00072214 3.3 0.00072224 0 0.00072216 0 0.00072226 3.3 0.00072218 3.3 0.00072228 0 0.0007222 0 0.0007222999999999999 3.3 0.0007222200000000001 3.3 0.00072232 0 0.0007222400000000001 0 0.00072234 3.3 0.0007222600000000001 3.3 0.00072236 0 0.0007222800000000001 0 0.00072238 3.3 0.0007223 3.3 0.0007224 0 0.00072232 0 0.00072242 3.3 0.00072234 3.3 0.00072244 0 0.00072236 0 0.00072246 3.3 0.00072238 3.3 0.00072248 0 0.0007224 0 0.0007224999999999999 3.3 0.00072242 3.3 0.0007225199999999999 0 0.0007224400000000001 0 0.00072254 3.3 0.0007224600000000001 3.3 0.00072256 0 0.0007224800000000001 0 0.00072258 3.3 0.0007225 3.3 0.0007226 0 0.00072252 0 0.00072262 3.3 0.00072254 3.3 0.00072264 0 0.00072256 0 0.00072266 3.3 0.00072258 3.3 0.00072268 0 0.0007226 0 0.0007227 3.3 0.00072262 3.3 0.0007227199999999999 0 0.0007226400000000001 0 0.00072274 3.3 0.0007226600000000001 3.3 0.00072276 0 0.0007226800000000001 0 0.00072278 3.3 0.0007227000000000001 3.3 0.0007228 0 0.00072272 0 0.00072282 3.3 0.00072274 3.3 0.00072284 0 0.00072276 0 0.00072286 3.3 0.00072278 3.3 0.00072288 0 0.0007228 0 0.0007229 3.3 0.00072282 3.3 0.0007229199999999999 0 0.00072284 0 0.0007229399999999999 3.3 0.0007228600000000001 3.3 0.00072296 0 0.0007228800000000001 0 0.00072298 3.3 0.0007229000000000001 3.3 0.000723 0 0.00072292 0 0.00072302 3.3 0.00072294 3.3 0.00072304 0 0.00072296 0 0.00072306 3.3 0.00072298 3.3 0.00072308 0 0.000723 0 0.0007231 3.3 0.00072302 3.3 0.00072312 0 0.00072304 0 0.0007231399999999999 3.3 0.0007230600000000001 3.3 0.00072316 0 0.0007230800000000001 0 0.00072318 3.3 0.0007231000000000001 3.3 0.0007232 0 0.0007231200000000001 0 0.00072322 3.3 0.00072314 3.3 0.00072324 0 0.00072316 0 0.00072326 3.3 0.00072318 3.3 0.00072328 0 0.0007232 0 0.0007233 3.3 0.00072322 3.3 0.00072332 0 0.00072324 0 0.0007233399999999999 3.3 0.00072326 3.3 0.0007233599999999999 0 0.0007232800000000001 0 0.00072338 3.3 0.0007233000000000001 3.3 0.0007234 0 0.0007233200000000001 0 0.00072342 3.3 0.00072334 3.3 0.00072344 0 0.00072336 0 0.00072346 3.3 0.00072338 3.3 0.00072348 0 0.0007234 0 0.0007235 3.3 0.00072342 3.3 0.00072352 0 0.00072344 0 0.00072354 3.3 0.00072346 3.3 0.0007235599999999999 0 0.0007234800000000001 0 0.00072358 3.3 0.0007235000000000001 3.3 0.0007236 0 0.0007235200000000001 0 0.00072362 3.3 0.0007235400000000001 3.3 0.00072364 0 0.00072356 0 0.00072366 3.3 0.00072358 3.3 0.00072368 0 0.0007236 0 0.0007237 3.3 0.00072362 3.3 0.00072372 0 0.00072364 0 0.00072374 3.3 0.00072366 3.3 0.0007237599999999999 0 0.0007236800000000001 0 0.00072378 3.3 0.0007237000000000001 3.3 0.0007238 0 0.0007237200000000001 0 0.00072382 3.3 0.0007237400000000001 3.3 0.00072384 0 0.00072376 0 0.00072386 3.3 0.00072378 3.3 0.00072388 0 0.0007238 0 0.0007239 3.3 0.00072382 3.3 0.00072392 0 0.00072384 0 0.00072394 3.3 0.00072386 3.3 0.00072396 0 0.00072388 0 0.0007239799999999999 3.3 0.0007239000000000001 3.3 0.000724 0 0.0007239200000000001 0 0.00072402 3.3 0.0007239400000000001 3.3 0.00072404 0 0.0007239600000000001 0 0.00072406 3.3 0.00072398 3.3 0.00072408 0 0.000724 0 0.0007241 3.3 0.00072402 3.3 0.00072412 0 0.00072404 0 0.00072414 3.3 0.00072406 3.3 0.00072416 0 0.00072408 0 0.0007241799999999999 3.3 0.0007241000000000001 3.3 0.0007242 0 0.0007241200000000001 0 0.00072422 3.3 0.0007241400000000001 3.3 0.00072424 0 0.0007241600000000001 0 0.00072426 3.3 0.00072418 3.3 0.00072428 0 0.0007242 0 0.0007243 3.3 0.00072422 3.3 0.00072432 0 0.00072424 0 0.00072434 3.3 0.00072426 3.3 0.00072436 0 0.00072428 0 0.00072438 3.3 0.0007243 3.3 0.0007243999999999999 0 0.0007243200000000001 0 0.00072442 3.3 0.0007243400000000001 3.3 0.00072444 0 0.0007243600000000001 0 0.00072446 3.3 0.0007243800000000001 3.3 0.00072448 0 0.0007244 0 0.0007245 3.3 0.00072442 3.3 0.00072452 0 0.00072444 0 0.00072454 3.3 0.00072446 3.3 0.00072456 0 0.00072448 0 0.00072458 3.3 0.0007245 3.3 0.0007245999999999999 0 0.0007245200000000001 0 0.00072462 3.3 0.0007245400000000001 3.3 0.00072464 0 0.0007245600000000001 0 0.00072466 3.3 0.0007245800000000001 3.3 0.00072468 0 0.0007246 0 0.0007247 3.3 0.00072462 3.3 0.00072472 0 0.00072464 0 0.00072474 3.3 0.00072466 3.3 0.00072476 0 0.00072468 0 0.00072478 3.3 0.0007247 3.3 0.0007247999999999999 0 0.00072472 0 0.0007248199999999999 3.3 0.0007247400000000001 3.3 0.00072484 0 0.0007247600000000001 0 0.00072486 3.3 0.0007247800000000001 3.3 0.00072488 0 0.0007248 0 0.0007249 3.3 0.00072482 3.3 0.00072492 0 0.00072484 0 0.00072494 3.3 0.00072486 3.3 0.00072496 0 0.00072488 0 0.00072498 3.3 0.0007249 3.3 0.000725 0 0.00072492 0 0.0007250199999999999 3.3 0.0007249400000000001 3.3 0.00072504 0 0.0007249600000000001 0 0.00072506 3.3 0.0007249800000000001 3.3 0.00072508 0 0.0007250000000000001 0 0.0007251 3.3 0.00072502 3.3 0.00072512 0 0.00072504 0 0.00072514 3.3 0.00072506 3.3 0.00072516 0 0.00072508 0 0.00072518 3.3 0.0007251 3.3 0.0007252 0 0.00072512 0 0.0007252199999999999 3.3 0.00072514 3.3 0.0007252399999999999 0 0.0007251600000000001 0 0.00072526 3.3 0.0007251800000000001 3.3 0.00072528 0 0.0007252000000000001 0 0.0007253 3.3 0.00072522 3.3 0.00072532 0 0.00072524 0 0.00072534 3.3 0.00072526 3.3 0.00072536 0 0.00072528 0 0.00072538 3.3 0.0007253 3.3 0.0007254 0 0.00072532 0 0.00072542 3.3 0.00072534 3.3 0.0007254399999999999 0 0.0007253600000000001 0 0.00072546 3.3 0.0007253800000000001 3.3 0.00072548 0 0.0007254000000000001 0 0.0007255 3.3 0.0007254200000000001 3.3 0.00072552 0 0.00072544 0 0.00072554 3.3 0.00072546 3.3 0.00072556 0 0.00072548 0 0.00072558 3.3 0.0007255 3.3 0.0007256 0 0.00072552 0 0.00072562 3.3 0.00072554 3.3 0.0007256399999999999 0 0.00072556 0 0.0007256599999999999 3.3 0.0007255800000000001 3.3 0.00072568 0 0.0007256000000000001 0 0.0007257 3.3 0.0007256200000000001 3.3 0.00072572 0 0.00072564 0 0.00072574 3.3 0.00072566 3.3 0.00072576 0 0.00072568 0 0.00072578 3.3 0.0007257 3.3 0.0007258 0 0.00072572 0 0.00072582 3.3 0.00072574 3.3 0.00072584 0 0.00072576 0 0.0007258599999999999 3.3 0.0007257800000000001 3.3 0.00072588 0 0.0007258000000000001 0 0.0007259 3.3 0.0007258200000000001 3.3 0.00072592 0 0.0007258400000000001 0 0.00072594 3.3 0.00072586 3.3 0.00072596 0 0.00072588 0 0.00072598 3.3 0.0007259 3.3 0.000726 0 0.00072592 0 0.00072602 3.3 0.00072594 3.3 0.00072604 0 0.00072596 0 0.0007260599999999999 3.3 0.00072598 3.3 0.0007260799999999999 0 0.0007260000000000001 0 0.0007261 3.3 0.0007260200000000001 3.3 0.00072612 0 0.0007260400000000001 0 0.00072614 3.3 0.00072606 3.3 0.00072616 0 0.00072608 0 0.00072618 3.3 0.0007261 3.3 0.0007262 0 0.00072612 0 0.00072622 3.3 0.00072614 3.3 0.00072624 0 0.00072616 0 0.00072626 3.3 0.00072618 3.3 0.0007262799999999999 0 0.0007262000000000001 0 0.0007263 3.3 0.0007262200000000001 3.3 0.00072632 0 0.0007262400000000001 0 0.00072634 3.3 0.0007262600000000001 3.3 0.00072636 0 0.00072628 0 0.00072638 3.3 0.0007263 3.3 0.0007264 0 0.00072632 0 0.00072642 3.3 0.00072634 3.3 0.00072644 0 0.00072636 0 0.00072646 3.3 0.00072638 3.3 0.0007264799999999999 0 0.0007264 0 0.0007264999999999999 3.3 0.0007264200000000001 3.3 0.00072652 0 0.0007264400000000001 0 0.00072654 3.3 0.0007264600000000001 3.3 0.00072656 0 0.00072648 0 0.00072658 3.3 0.0007265 3.3 0.0007266 0 0.00072652 0 0.00072662 3.3 0.00072654 3.3 0.00072664 0 0.00072656 0 0.00072666 3.3 0.00072658 3.3 0.00072668 0 0.0007266 0 0.0007266999999999999 3.3 0.0007266200000000001 3.3 0.00072672 0 0.0007266400000000001 0 0.00072674 3.3 0.0007266600000000001 3.3 0.00072676 0 0.0007266800000000001 0 0.00072678 3.3 0.0007267 3.3 0.0007268 0 0.00072672 0 0.00072682 3.3 0.00072674 3.3 0.00072684 0 0.00072676 0 0.00072686 3.3 0.00072678 3.3 0.00072688 0 0.0007268 0 0.0007268999999999999 3.3 0.00072682 3.3 0.0007269199999999999 0 0.0007268400000000001 0 0.00072694 3.3 0.0007268600000000001 3.3 0.00072696 0 0.0007268800000000001 0 0.00072698 3.3 0.0007269 3.3 0.000727 0 0.00072692 0 0.00072702 3.3 0.00072694 3.3 0.00072704 0 0.00072696 0 0.00072706 3.3 0.00072698 3.3 0.00072708 0 0.000727 0 0.0007271 3.3 0.00072702 3.3 0.0007271199999999999 0 0.0007270400000000001 0 0.00072714 3.3 0.0007270600000000001 3.3 0.00072716 0 0.0007270800000000001 0 0.00072718 3.3 0.0007271000000000001 3.3 0.0007272 0 0.00072712 0 0.00072722 3.3 0.00072714 3.3 0.00072724 0 0.00072716 0 0.00072726 3.3 0.00072718 3.3 0.00072728 0 0.0007272 0 0.0007273 3.3 0.00072722 3.3 0.0007273199999999999 0 0.0007272400000000001 0 0.00072734 3.3 0.0007272600000000001 3.3 0.00072736 0 0.0007272800000000001 0 0.00072738 3.3 0.0007273000000000001 3.3 0.0007274 0 0.00072732 0 0.00072742 3.3 0.00072734 3.3 0.00072744 0 0.00072736 0 0.00072746 3.3 0.00072738 3.3 0.00072748 0 0.0007274 0 0.0007275 3.3 0.00072742 3.3 0.00072752 0 0.00072744 0 0.0007275399999999999 3.3 0.0007274600000000001 3.3 0.00072756 0 0.0007274800000000001 0 0.00072758 3.3 0.0007275000000000001 3.3 0.0007276 0 0.0007275200000000001 0 0.00072762 3.3 0.00072754 3.3 0.00072764 0 0.00072756 0 0.00072766 3.3 0.00072758 3.3 0.00072768 0 0.0007276 0 0.0007277 3.3 0.00072762 3.3 0.00072772 0 0.00072764 0 0.0007277399999999999 3.3 0.0007276600000000001 3.3 0.00072776 0 0.0007276800000000001 0 0.00072778 3.3 0.0007277000000000001 3.3 0.0007278 0 0.0007277200000000001 0 0.00072782 3.3 0.00072774 3.3 0.00072784 0 0.00072776 0 0.00072786 3.3 0.00072778 3.3 0.00072788 0 0.0007278 0 0.0007279 3.3 0.00072782 3.3 0.00072792 0 0.00072784 0 0.0007279399999999999 3.3 0.00072786 3.3 0.0007279599999999999 0 0.0007278800000000001 0 0.00072798 3.3 0.0007279000000000001 3.3 0.000728 0 0.0007279200000000001 0 0.00072802 3.3 0.00072794 3.3 0.00072804 0 0.00072796 0 0.00072806 3.3 0.00072798 3.3 0.00072808 0 0.000728 0 0.0007281 3.3 0.00072802 3.3 0.00072812 0 0.00072804 0 0.00072814 3.3 0.00072806 3.3 0.0007281599999999999 0 0.0007280800000000001 0 0.00072818 3.3 0.0007281000000000001 3.3 0.0007282 0 0.0007281200000000001 0 0.00072822 3.3 0.0007281400000000001 3.3 0.00072824 0 0.00072816 0 0.00072826 3.3 0.00072818 3.3 0.00072828 0 0.0007282 0 0.0007283 3.3 0.00072822 3.3 0.00072832 0 0.00072824 0 0.00072834 3.3 0.00072826 3.3 0.0007283599999999999 0 0.00072828 0 0.0007283799999999999 3.3 0.0007283000000000001 3.3 0.0007284 0 0.0007283200000000001 0 0.00072842 3.3 0.0007283400000000001 3.3 0.00072844 0 0.00072836 0 0.00072846 3.3 0.00072838 3.3 0.00072848 0 0.0007284 0 0.0007285 3.3 0.00072842 3.3 0.00072852 0 0.00072844 0 0.00072854 3.3 0.00072846 3.3 0.00072856 0 0.00072848 0 0.0007285799999999999 3.3 0.0007285000000000001 3.3 0.0007286 0 0.0007285200000000001 0 0.00072862 3.3 0.0007285400000000001 3.3 0.00072864 0 0.0007285600000000001 0 0.00072866 3.3 0.00072858 3.3 0.00072868 0 0.0007286 0 0.0007287 3.3 0.00072862 3.3 0.00072872 0 0.00072864 0 0.00072874 3.3 0.00072866 3.3 0.00072876 0 0.00072868 0 0.0007287799999999999 3.3 0.0007287 3.3 0.0007287999999999999 0 0.0007287200000000001 0 0.00072882 3.3 0.0007287400000000001 3.3 0.00072884 0 0.0007287600000000001 0 0.00072886 3.3 0.00072878 3.3 0.00072888 0 0.0007288 0 0.0007289 3.3 0.00072882 3.3 0.00072892 0 0.00072884 0 0.00072894 3.3 0.00072886 3.3 0.00072896 0 0.00072888 0 0.00072898 3.3 0.0007289 3.3 0.0007289999999999999 0 0.0007289200000000001 0 0.00072902 3.3 0.0007289400000000001 3.3 0.00072904 0 0.0007289600000000001 0 0.00072906 3.3 0.0007289800000000001 3.3 0.00072908 0 0.000729 0 0.0007291 3.3 0.00072902 3.3 0.00072912 0 0.00072904 0 0.00072914 3.3 0.00072906 3.3 0.00072916 0 0.00072908 0 0.00072918 3.3 0.0007291 3.3 0.0007291999999999999 0 0.00072912 0 0.0007292199999999999 3.3 0.0007291400000000001 3.3 0.00072924 0 0.0007291600000000001 0 0.00072926 3.3 0.0007291800000000001 3.3 0.00072928 0 0.0007292 0 0.0007293 3.3 0.00072922 3.3 0.00072932 0 0.00072924 0 0.00072934 3.3 0.00072926 3.3 0.00072936 0 0.00072928 0 0.00072938 3.3 0.0007293 3.3 0.0007294 0 0.00072932 0 0.0007294199999999999 3.3 0.0007293400000000001 3.3 0.00072944 0 0.0007293600000000001 0 0.00072946 3.3 0.0007293800000000001 3.3 0.00072948 0 0.0007294000000000001 0 0.0007295 3.3 0.00072942 3.3 0.00072952 0 0.00072944 0 0.00072954 3.3 0.00072946 3.3 0.00072956 0 0.00072948 0 0.00072958 3.3 0.0007295 3.3 0.0007296 0 0.00072952 0 0.0007296199999999999 3.3 0.00072954 3.3 0.0007296399999999999 0 0.0007295600000000001 0 0.00072966 3.3 0.0007295800000000001 3.3 0.00072968 0 0.0007296000000000001 0 0.0007297 3.3 0.00072962 3.3 0.00072972 0 0.00072964 0 0.00072974 3.3 0.00072966 3.3 0.00072976 0 0.00072968 0 0.00072978 3.3 0.0007297 3.3 0.0007298 0 0.00072972 0 0.00072982 3.3 0.00072974 3.3 0.0007298399999999999 0 0.0007297600000000001 0 0.00072986 3.3 0.0007297800000000001 3.3 0.00072988 0 0.0007298000000000001 0 0.0007299 3.3 0.0007298200000000001 3.3 0.00072992 0 0.00072984 0 0.00072994 3.3 0.00072986 3.3 0.00072996 0 0.00072988 0 0.00072998 3.3 0.0007299 3.3 0.00073 0 0.00072992 0 0.00073002 3.3 0.00072994 3.3 0.0007300399999999999 0 0.00072996 0 0.0007300599999999999 3.3 0.0007299800000000001 3.3 0.00073008 0 0.0007300000000000001 0 0.0007301 3.3 0.0007300200000000001 3.3 0.00073012 0 0.00073004 0 0.00073014 3.3 0.00073006 3.3 0.00073016 0 0.00073008 0 0.00073018 3.3 0.0007301 3.3 0.0007302 0 0.00073012 0 0.00073022 3.3 0.00073014 3.3 0.00073024 0 0.00073016 0 0.0007302599999999999 3.3 0.0007301800000000001 3.3 0.00073028 0 0.0007302000000000001 0 0.0007303 3.3 0.0007302200000000001 3.3 0.00073032 0 0.0007302400000000001 0 0.00073034 3.3 0.00073026 3.3 0.00073036 0 0.00073028 0 0.00073038 3.3 0.0007303 3.3 0.0007304 0 0.00073032 0 0.00073042 3.3 0.00073034 3.3 0.00073044 0 0.00073036 0 0.0007304599999999999 3.3 0.00073038 3.3 0.0007304799999999999 0 0.0007304000000000001 0 0.0007305 3.3 0.0007304200000000001 3.3 0.00073052 0 0.0007304400000000001 0 0.00073054 3.3 0.00073046 3.3 0.00073056 0 0.00073048 0 0.00073058 3.3 0.0007305 3.3 0.0007306 0 0.00073052 0 0.00073062 3.3 0.00073054 3.3 0.00073064 0 0.00073056 0 0.00073066 3.3 0.00073058 3.3 0.0007306799999999999 0 0.0007306000000000001 0 0.0007307 3.3 0.0007306200000000001 3.3 0.00073072 0 0.0007306400000000001 0 0.00073074 3.3 0.0007306600000000001 3.3 0.00073076 0 0.00073068 0 0.00073078 3.3 0.0007307 3.3 0.0007308 0 0.00073072 0 0.00073082 3.3 0.00073074 3.3 0.00073084 0 0.00073076 0 0.00073086 3.3 0.00073078 3.3 0.0007308799999999999 0 0.0007308000000000001 0 0.0007309 3.3 0.0007308200000000001 3.3 0.00073092 0 0.0007308400000000001 0 0.00073094 3.3 0.0007308600000000001 3.3 0.00073096 0 0.00073088 0 0.00073098 3.3 0.0007309 3.3 0.000731 0 0.00073092 0 0.00073102 3.3 0.00073094 3.3 0.00073104 0 0.00073096 0 0.00073106 3.3 0.00073098 3.3 0.00073108 0 0.000731 0 0.0007310999999999999 3.3 0.0007310200000000001 3.3 0.00073112 0 0.0007310400000000001 0 0.00073114 3.3 0.0007310600000000001 3.3 0.00073116 0 0.0007310800000000001 0 0.00073118 3.3 0.0007311 3.3 0.0007312 0 0.00073112 0 0.00073122 3.3 0.00073114 3.3 0.00073124 0 0.00073116 0 0.00073126 3.3 0.00073118 3.3 0.00073128 0 0.0007312 0 0.0007312999999999999 3.3 0.0007312200000000001 3.3 0.00073132 0 0.0007312400000000001 0 0.00073134 3.3 0.0007312600000000001 3.3 0.00073136 0 0.0007312800000000001 0 0.00073138 3.3 0.0007313 3.3 0.0007314 0 0.00073132 0 0.00073142 3.3 0.00073134 3.3 0.00073144 0 0.00073136 0 0.00073146 3.3 0.00073138 3.3 0.00073148 0 0.0007314 0 0.0007314999999999999 3.3 0.00073142 3.3 0.0007315199999999999 0 0.0007314400000000001 0 0.00073154 3.3 0.0007314600000000001 3.3 0.00073156 0 0.0007314800000000001 0 0.00073158 3.3 0.0007315 3.3 0.0007316 0 0.00073152 0 0.00073162 3.3 0.00073154 3.3 0.00073164 0 0.00073156 0 0.00073166 3.3 0.00073158 3.3 0.00073168 0 0.0007316 0 0.0007317 3.3 0.00073162 3.3 0.0007317199999999999 0 0.0007316400000000001 0 0.00073174 3.3 0.0007316600000000001 3.3 0.00073176 0 0.0007316800000000001 0 0.00073178 3.3 0.0007317000000000001 3.3 0.0007318 0 0.00073172 0 0.00073182 3.3 0.00073174 3.3 0.00073184 0 0.00073176 0 0.00073186 3.3 0.00073178 3.3 0.00073188 0 0.0007318 0 0.0007319 3.3 0.00073182 3.3 0.0007319199999999999 0 0.00073184 0 0.0007319399999999999 3.3 0.0007318600000000001 3.3 0.00073196 0 0.0007318800000000001 0 0.00073198 3.3 0.0007319000000000001 3.3 0.000732 0 0.00073192 0 0.00073202 3.3 0.00073194 3.3 0.00073204 0 0.00073196 0 0.00073206 3.3 0.00073198 3.3 0.00073208 0 0.000732 0 0.0007321 3.3 0.00073202 3.3 0.00073212 0 0.00073204 0 0.0007321399999999999 3.3 0.0007320600000000001 3.3 0.00073216 0 0.0007320800000000001 0 0.00073218 3.3 0.0007321000000000001 3.3 0.0007322 0 0.0007321200000000001 0 0.00073222 3.3 0.00073214 3.3 0.00073224 0 0.00073216 0 0.00073226 3.3 0.00073218 3.3 0.00073228 0 0.0007322 0 0.0007323 3.3 0.00073222 3.3 0.00073232 0 0.00073224 0 0.0007323399999999999 3.3 0.00073226 3.3 0.0007323599999999999 0 0.0007322800000000001 0 0.00073238 3.3 0.0007323000000000001 3.3 0.0007324 0 0.0007323200000000001 0 0.00073242 3.3 0.00073234 3.3 0.00073244 0 0.00073236 0 0.00073246 3.3 0.00073238 3.3 0.00073248 0 0.0007324 0 0.0007325 3.3 0.00073242 3.3 0.00073252 0 0.00073244 0 0.00073254 3.3 0.00073246 3.3 0.0007325599999999999 0 0.0007324800000000001 0 0.00073258 3.3 0.0007325000000000001 3.3 0.0007326 0 0.0007325200000000001 0 0.00073262 3.3 0.0007325400000000001 3.3 0.00073264 0 0.00073256 0 0.00073266 3.3 0.00073258 3.3 0.00073268 0 0.0007326 0 0.0007327 3.3 0.00073262 3.3 0.00073272 0 0.00073264 0 0.00073274 3.3 0.00073266 3.3 0.0007327599999999999 0 0.00073268 0 0.0007327799999999999 3.3 0.0007327000000000001 3.3 0.0007328 0 0.0007327200000000001 0 0.00073282 3.3 0.0007327400000000001 3.3 0.00073284 0 0.00073276 0 0.00073286 3.3 0.00073278 3.3 0.00073288 0 0.0007328 0 0.0007329 3.3 0.00073282 3.3 0.00073292 0 0.00073284 0 0.00073294 3.3 0.00073286 3.3 0.00073296 0 0.00073288 0 0.0007329799999999999 3.3 0.0007329000000000001 3.3 0.000733 0 0.0007329200000000001 0 0.00073302 3.3 0.0007329400000000001 3.3 0.00073304 0 0.0007329600000000001 0 0.00073306 3.3 0.00073298 3.3 0.00073308 0 0.000733 0 0.0007331 3.3 0.00073302 3.3 0.00073312 0 0.00073304 0 0.00073314 3.3 0.00073306 3.3 0.00073316 0 0.00073308 0 0.0007331799999999999 3.3 0.0007331 3.3 0.0007331999999999999 0 0.0007331200000000001 0 0.00073322 3.3 0.0007331400000000001 3.3 0.00073324 0 0.0007331600000000001 0 0.00073326 3.3 0.00073318 3.3 0.00073328 0 0.0007332 0 0.0007333 3.3 0.00073322 3.3 0.00073332 0 0.00073324 0 0.00073334 3.3 0.00073326 3.3 0.00073336 0 0.00073328 0 0.00073338 3.3 0.0007333 3.3 0.0007333999999999999 0 0.0007333200000000001 0 0.00073342 3.3 0.0007333400000000001 3.3 0.00073344 0 0.0007333600000000001 0 0.00073346 3.3 0.0007333800000000001 3.3 0.00073348 0 0.0007334 0 0.0007335 3.3 0.00073342 3.3 0.00073352 0 0.00073344 0 0.00073354 3.3 0.00073346 3.3 0.00073356 0 0.00073348 0 0.00073358 3.3 0.0007335 3.3 0.0007335999999999999 0 0.00073352 0 0.0007336199999999999 3.3 0.0007335400000000001 3.3 0.00073364 0 0.0007335600000000001 0 0.00073366 3.3 0.0007335800000000001 3.3 0.00073368 0 0.0007336 0 0.0007337 3.3 0.00073362 3.3 0.00073372 0 0.00073364 0 0.00073374 3.3 0.00073366 3.3 0.00073376 0 0.00073368 0 0.00073378 3.3 0.0007337 3.3 0.0007338 0 0.00073372 0 0.0007338199999999999 3.3 0.0007337400000000001 3.3 0.00073384 0 0.0007337600000000001 0 0.00073386 3.3 0.0007337800000000001 3.3 0.00073388 0 0.0007338000000000001 0 0.0007339 3.3 0.00073382 3.3 0.00073392 0 0.00073384 0 0.00073394 3.3 0.00073386 3.3 0.00073396 0 0.00073388 0 0.00073398 3.3 0.0007339 3.3 0.000734 0 0.00073392 0 0.0007340199999999999 3.3 0.00073394 3.3 0.0007340399999999999 0 0.0007339600000000001 0 0.00073406 3.3 0.0007339800000000001 3.3 0.00073408 0 0.0007340000000000001 0 0.0007341 3.3 0.00073402 3.3 0.00073412 0 0.00073404 0 0.00073414 3.3 0.00073406 3.3 0.00073416 0 0.00073408 0 0.00073418 3.3 0.0007341 3.3 0.0007342 0 0.00073412 0 0.00073422 3.3 0.00073414 3.3 0.0007342399999999999 0 0.0007341600000000001 0 0.00073426 3.3 0.0007341800000000001 3.3 0.00073428 0 0.0007342000000000001 0 0.0007343 3.3 0.0007342200000000001 3.3 0.00073432 0 0.00073424 0 0.00073434 3.3 0.00073426 3.3 0.00073436 0 0.00073428 0 0.00073438 3.3 0.0007343 3.3 0.0007344 0 0.00073432 0 0.00073442 3.3 0.00073434 3.3 0.0007344399999999999 0 0.0007343600000000001 0 0.00073446 3.3 0.0007343800000000001 3.3 0.00073448 0 0.0007344000000000001 0 0.0007345 3.3 0.0007344200000000001 3.3 0.00073452 0 0.00073444 0 0.00073454 3.3 0.00073446 3.3 0.00073456 0 0.00073448 0 0.00073458 3.3 0.0007345 3.3 0.0007346 0 0.00073452 0 0.00073462 3.3 0.00073454 3.3 0.00073464 0 0.00073456 0 0.0007346599999999999 3.3 0.0007345800000000001 3.3 0.00073468 0 0.0007346000000000001 0 0.0007347 3.3 0.0007346200000000001 3.3 0.00073472 0 0.0007346400000000001 0 0.00073474 3.3 0.00073466 3.3 0.00073476 0 0.00073468 0 0.00073478 3.3 0.0007347 3.3 0.0007348 0 0.00073472 0 0.00073482 3.3 0.00073474 3.3 0.00073484 0 0.00073476 0 0.0007348599999999999 3.3 0.0007347800000000001 3.3 0.00073488 0 0.0007348000000000001 0 0.0007349 3.3 0.0007348200000000001 3.3 0.00073492 0 0.0007348400000000001 0 0.00073494 3.3 0.00073486 3.3 0.00073496 0 0.00073488 0 0.00073498 3.3 0.0007349 3.3 0.000735 0 0.00073492 0 0.00073502 3.3 0.00073494 3.3 0.00073504 0 0.00073496 0 0.0007350599999999999 3.3 0.00073498 3.3 0.0007350799999999999 0 0.0007350000000000001 0 0.0007351 3.3 0.0007350200000000001 3.3 0.00073512 0 0.0007350400000000001 0 0.00073514 3.3 0.00073506 3.3 0.00073516 0 0.00073508 0 0.00073518 3.3 0.0007351 3.3 0.0007352 0 0.00073512 0 0.00073522 3.3 0.00073514 3.3 0.00073524 0 0.00073516 0 0.00073526 3.3 0.00073518 3.3 0.0007352799999999999 0 0.0007352000000000001 0 0.0007353 3.3 0.0007352200000000001 3.3 0.00073532 0 0.0007352400000000001 0 0.00073534 3.3 0.0007352600000000001 3.3 0.00073536 0 0.00073528 0 0.00073538 3.3 0.0007353 3.3 0.0007354 0 0.00073532 0 0.00073542 3.3 0.00073534 3.3 0.00073544 0 0.00073536 0 0.00073546 3.3 0.00073538 3.3 0.0007354799999999999 0 0.0007354 0 0.0007354999999999999 3.3 0.0007354200000000001 3.3 0.00073552 0 0.0007354400000000001 0 0.00073554 3.3 0.0007354600000000001 3.3 0.00073556 0 0.00073548 0 0.00073558 3.3 0.0007355 3.3 0.0007356 0 0.00073552 0 0.00073562 3.3 0.00073554 3.3 0.00073564 0 0.00073556 0 0.00073566 3.3 0.00073558 3.3 0.00073568 0 0.0007356 0 0.0007356999999999999 3.3 0.0007356200000000001 3.3 0.00073572 0 0.0007356400000000001 0 0.00073574 3.3 0.0007356600000000001 3.3 0.00073576 0 0.0007356800000000001 0 0.00073578 3.3 0.0007357 3.3 0.0007358 0 0.00073572 0 0.00073582 3.3 0.00073574 3.3 0.00073584 0 0.00073576 0 0.00073586 3.3 0.00073578 3.3 0.00073588 0 0.0007358 0 0.0007358999999999999 3.3 0.00073582 3.3 0.0007359199999999999 0 0.0007358400000000001 0 0.00073594 3.3 0.0007358600000000001 3.3 0.00073596 0 0.0007358800000000001 0 0.00073598 3.3 0.0007359 3.3 0.000736 0 0.00073592 0 0.00073602 3.3 0.00073594 3.3 0.00073604 0 0.00073596 0 0.00073606 3.3 0.00073598 3.3 0.00073608 0 0.000736 0 0.0007361 3.3 0.00073602 3.3 0.0007361199999999999 0 0.0007360400000000001 0 0.00073614 3.3 0.0007360600000000001 3.3 0.00073616 0 0.0007360800000000001 0 0.00073618 3.3 0.0007361000000000001 3.3 0.0007362 0 0.00073612 0 0.00073622 3.3 0.00073614 3.3 0.00073624 0 0.00073616 0 0.00073626 3.3 0.00073618 3.3 0.00073628 0 0.0007362 0 0.0007363 3.3 0.00073622 3.3 0.0007363199999999999 0 0.00073624 0 0.0007363399999999999 3.3 0.0007362600000000001 3.3 0.00073636 0 0.0007362800000000001 0 0.00073638 3.3 0.0007363000000000001 3.3 0.0007364 0 0.00073632 0 0.00073642 3.3 0.00073634 3.3 0.00073644 0 0.00073636 0 0.00073646 3.3 0.00073638 3.3 0.00073648 0 0.0007364 0 0.0007365 3.3 0.00073642 3.3 0.00073652 0 0.00073644 0 0.0007365399999999999 3.3 0.0007364600000000001 3.3 0.00073656 0 0.0007364800000000001 0 0.00073658 3.3 0.0007365000000000001 3.3 0.0007366 0 0.0007365200000000001 0 0.00073662 3.3 0.00073654 3.3 0.00073664 0 0.00073656 0 0.00073666 3.3 0.00073658 3.3 0.00073668 0 0.0007366 0 0.0007367 3.3 0.00073662 3.3 0.00073672 0 0.00073664 0 0.0007367399999999999 3.3 0.00073666 3.3 0.0007367599999999999 0 0.0007366800000000001 0 0.00073678 3.3 0.0007367000000000001 3.3 0.0007368 0 0.0007367200000000001 0 0.00073682 3.3 0.00073674 3.3 0.00073684 0 0.00073676 0 0.00073686 3.3 0.00073678 3.3 0.00073688 0 0.0007368 0 0.0007369 3.3 0.00073682 3.3 0.00073692 0 0.00073684 0 0.00073694 3.3 0.00073686 3.3 0.0007369599999999999 0 0.0007368800000000001 0 0.00073698 3.3 0.0007369000000000001 3.3 0.000737 0 0.0007369200000000001 0 0.00073702 3.3 0.0007369400000000001 3.3 0.00073704 0 0.00073696 0 0.00073706 3.3 0.00073698 3.3 0.00073708 0 0.000737 0 0.0007371 3.3 0.00073702 3.3 0.00073712 0 0.00073704 0 0.00073714 3.3 0.00073706 3.3 0.0007371599999999999 0 0.00073708 0 0.0007371799999999999 3.3 0.0007371000000000001 3.3 0.0007372 0 0.0007371200000000001 0 0.00073722 3.3 0.0007371400000000001 3.3 0.00073724 0 0.00073716 0 0.00073726 3.3 0.00073718 3.3 0.00073728 0 0.0007372 0 0.0007373 3.3 0.00073722 3.3 0.00073732 0 0.00073724 0 0.00073734 3.3 0.00073726 3.3 0.00073736 0 0.00073728 0 0.0007373799999999999 3.3 0.0007373000000000001 3.3 0.0007374 0 0.0007373200000000001 0 0.00073742 3.3 0.0007373400000000001 3.3 0.00073744 0 0.0007373600000000001 0 0.00073746 3.3 0.00073738 3.3 0.00073748 0 0.0007374 0 0.0007375 3.3 0.00073742 3.3 0.00073752 0 0.00073744 0 0.00073754 3.3 0.00073746 3.3 0.00073756 0 0.00073748 0 0.0007375799999999999 3.3 0.0007375 3.3 0.0007375999999999999 0 0.0007375200000000001 0 0.00073762 3.3 0.0007375400000000001 3.3 0.00073764 0 0.0007375600000000001 0 0.00073766 3.3 0.00073758 3.3 0.00073768 0 0.0007376 0 0.0007377 3.3 0.00073762 3.3 0.00073772 0 0.00073764 0 0.00073774 3.3 0.00073766 3.3 0.00073776 0 0.00073768 0 0.00073778 3.3 0.0007377 3.3 0.0007377999999999999 0 0.0007377200000000001 0 0.00073782 3.3 0.0007377400000000001 3.3 0.00073784 0 0.0007377600000000001 0 0.00073786 3.3 0.0007377800000000001 3.3 0.00073788 0 0.0007378 0 0.0007379 3.3 0.00073782 3.3 0.00073792 0 0.00073784 0 0.00073794 3.3 0.00073786 3.3 0.00073796 0 0.00073788 0 0.00073798 3.3 0.0007379 3.3 0.0007379999999999999 0 0.0007379200000000001 0 0.00073802 3.3 0.0007379400000000001 3.3 0.00073804 0 0.0007379600000000001 0 0.00073806 3.3 0.0007379800000000001 3.3 0.00073808 0 0.000738 0 0.0007381 3.3 0.00073802 3.3 0.00073812 0 0.00073804 0 0.00073814 3.3 0.00073806 3.3 0.00073816 0 0.00073808 0 0.00073818 3.3 0.0007381 3.3 0.0007381999999999999 0 0.00073812 0 0.0007382199999999999 3.3 0.0007381400000000001 3.3 0.00073824 0 0.0007381600000000001 0 0.00073826 3.3 0.0007381800000000001 3.3 0.00073828 0 0.0007382 0 0.0007383 3.3 0.00073822 3.3 0.00073832 0 0.00073824 0 0.00073834 3.3 0.00073826 3.3 0.00073836 0 0.00073828 0 0.00073838 3.3 0.0007383 3.3 0.0007384 0 0.00073832 0 0.0007384199999999999 3.3 0.0007383400000000001 3.3 0.00073844 0 0.0007383600000000001 0 0.00073846 3.3 0.0007383800000000001 3.3 0.00073848 0 0.0007384000000000001 0 0.0007385 3.3 0.00073842 3.3 0.00073852 0 0.00073844 0 0.00073854 3.3 0.00073846 3.3 0.00073856 0 0.00073848 0 0.00073858 3.3 0.0007385 3.3 0.0007386 0 0.00073852 0 0.0007386199999999999 3.3 0.00073854 3.3 0.0007386399999999999 0 0.0007385600000000001 0 0.00073866 3.3 0.0007385800000000001 3.3 0.00073868 0 0.0007386000000000001 0 0.0007387 3.3 0.00073862 3.3 0.00073872 0 0.00073864 0 0.00073874 3.3 0.00073866 3.3 0.00073876 0 0.00073868 0 0.00073878 3.3 0.0007387 3.3 0.0007388 0 0.00073872 0 0.00073882 3.3 0.00073874 3.3 0.0007388399999999999 0 0.0007387600000000001 0 0.00073886 3.3 0.0007387800000000001 3.3 0.00073888 0 0.0007388000000000001 0 0.0007389 3.3 0.0007388200000000001 3.3 0.00073892 0 0.00073884 0 0.00073894 3.3 0.00073886 3.3 0.00073896 0 0.00073888 0 0.00073898 3.3 0.0007389 3.3 0.000739 0 0.00073892 0 0.00073902 3.3 0.00073894 3.3 0.0007390399999999999 0 0.00073896 0 0.0007390599999999999 3.3 0.0007389800000000001 3.3 0.00073908 0 0.0007390000000000001 0 0.0007391 3.3 0.0007390200000000001 3.3 0.00073912 0 0.00073904 0 0.00073914 3.3 0.00073906 3.3 0.00073916 0 0.00073908 0 0.00073918 3.3 0.0007391 3.3 0.0007392 0 0.00073912 0 0.00073922 3.3 0.00073914 3.3 0.00073924 0 0.00073916 0 0.0007392599999999999 3.3 0.0007391800000000001 3.3 0.00073928 0 0.0007392000000000001 0 0.0007393 3.3 0.0007392200000000001 3.3 0.00073932 0 0.0007392400000000001 0 0.00073934 3.3 0.00073926 3.3 0.00073936 0 0.00073928 0 0.00073938 3.3 0.0007393 3.3 0.0007394 0 0.00073932 0 0.00073942 3.3 0.00073934 3.3 0.00073944 0 0.00073936 0 0.0007394599999999999 3.3 0.00073938 3.3 0.0007394799999999999 0 0.0007394000000000001 0 0.0007395 3.3 0.0007394200000000001 3.3 0.00073952 0 0.0007394400000000001 0 0.00073954 3.3 0.00073946 3.3 0.00073956 0 0.00073948 0 0.00073958 3.3 0.0007395 3.3 0.0007396 0 0.00073952 0 0.00073962 3.3 0.00073954 3.3 0.00073964 0 0.00073956 0 0.00073966 3.3 0.00073958 3.3 0.0007396799999999999 0 0.0007396000000000001 0 0.0007397 3.3 0.0007396200000000001 3.3 0.00073972 0 0.0007396400000000001 0 0.00073974 3.3 0.0007396600000000001 3.3 0.00073976 0 0.00073968 0 0.00073978 3.3 0.0007397 3.3 0.0007398 0 0.00073972 0 0.00073982 3.3 0.00073974 3.3 0.00073984 0 0.00073976 0 0.00073986 3.3 0.00073978 3.3 0.0007398799999999999 0 0.0007398 0 0.0007398999999999999 3.3 0.0007398200000000001 3.3 0.00073992 0 0.0007398400000000001 0 0.00073994 3.3 0.0007398600000000001 3.3 0.00073996 0 0.00073988 0 0.00073998 3.3 0.0007399 3.3 0.00074 0 0.00073992 0 0.00074002 3.3 0.00073994 3.3 0.00074004 0 0.00073996 0 0.00074006 3.3 0.00073998 3.3 0.00074008 0 0.00074 0 0.0007400999999999999 3.3 0.0007400200000000001 3.3 0.00074012 0 0.0007400400000000001 0 0.00074014 3.3 0.0007400600000000001 3.3 0.00074016 0 0.0007400800000000001 0 0.00074018 3.3 0.0007401 3.3 0.0007402 0 0.00074012 0 0.00074022 3.3 0.00074014 3.3 0.00074024 0 0.00074016 0 0.00074026 3.3 0.00074018 3.3 0.00074028 0 0.0007402 0 0.0007402999999999999 3.3 0.00074022 3.3 0.0007403199999999999 0 0.0007402400000000001 0 0.00074034 3.3 0.0007402600000000001 3.3 0.00074036 0 0.0007402800000000001 0 0.00074038 3.3 0.0007403 3.3 0.0007404 0 0.00074032 0 0.00074042 3.3 0.00074034 3.3 0.00074044 0 0.00074036 0 0.00074046 3.3 0.00074038 3.3 0.00074048 0 0.0007404 0 0.0007405 3.3 0.00074042 3.3 0.0007405199999999999 0 0.0007404400000000001 0 0.00074054 3.3 0.0007404600000000001 3.3 0.00074056 0 0.0007404800000000001 0 0.00074058 3.3 0.0007405000000000001 3.3 0.0007406 0 0.00074052 0 0.00074062 3.3 0.00074054 3.3 0.00074064 0 0.00074056 0 0.00074066 3.3 0.00074058 3.3 0.00074068 0 0.0007406 0 0.0007407 3.3 0.00074062 3.3 0.0007407199999999999 0 0.00074064 0 0.0007407399999999999 3.3 0.0007406600000000001 3.3 0.00074076 0 0.0007406800000000001 0 0.00074078 3.3 0.0007407000000000001 3.3 0.0007408 0 0.00074072 0 0.00074082 3.3 0.00074074 3.3 0.00074084 0 0.00074076 0 0.00074086 3.3 0.00074078 3.3 0.00074088 0 0.0007408 0 0.0007409 3.3 0.00074082 3.3 0.00074092 0 0.00074084 0 0.0007409399999999999 3.3 0.0007408600000000001 3.3 0.00074096 0 0.0007408800000000001 0 0.00074098 3.3 0.0007409000000000001 3.3 0.000741 0 0.0007409200000000001 0 0.00074102 3.3 0.00074094 3.3 0.00074104 0 0.00074096 0 0.00074106 3.3 0.00074098 3.3 0.00074108 0 0.000741 0 0.0007411 3.3 0.00074102 3.3 0.00074112 0 0.00074104 0 0.0007411399999999999 3.3 0.0007410600000000001 3.3 0.00074116 0 0.0007410800000000001 0 0.00074118 3.3 0.0007411000000000001 3.3 0.0007412 0 0.0007411200000000001 0 0.00074122 3.3 0.00074114 3.3 0.00074124 0 0.00074116 0 0.00074126 3.3 0.00074118 3.3 0.00074128 0 0.0007412 0 0.0007413 3.3 0.00074122 3.3 0.00074132 0 0.00074124 0 0.00074134 3.3 0.00074126 3.3 0.0007413599999999999 0 0.0007412800000000001 0 0.00074138 3.3 0.0007413000000000001 3.3 0.0007414 0 0.0007413200000000001 0 0.00074142 3.3 0.0007413400000000001 3.3 0.00074144 0 0.00074136 0 0.00074146 3.3 0.00074138 3.3 0.00074148 0 0.0007414 0 0.0007415 3.3 0.00074142 3.3 0.00074152 0 0.00074144 0 0.00074154 3.3 0.00074146 3.3 0.0007415599999999999 0 0.0007414800000000001 0 0.00074158 3.3 0.0007415000000000001 3.3 0.0007416 0 0.0007415200000000001 0 0.00074162 3.3 0.0007415400000000001 3.3 0.00074164 0 0.00074156 0 0.00074166 3.3 0.00074158 3.3 0.00074168 0 0.0007416 0 0.0007417 3.3 0.00074162 3.3 0.00074172 0 0.00074164 0 0.00074174 3.3 0.00074166 3.3 0.0007417599999999999 0 0.00074168 0 0.0007417799999999999 3.3 0.0007417000000000001 3.3 0.0007418 0 0.0007417200000000001 0 0.00074182 3.3 0.0007417400000000001 3.3 0.00074184 0 0.00074176 0 0.00074186 3.3 0.00074178 3.3 0.00074188 0 0.0007418 0 0.0007419 3.3 0.00074182 3.3 0.00074192 0 0.00074184 0 0.00074194 3.3 0.00074186 3.3 0.00074196 0 0.00074188 0 0.0007419799999999999 3.3 0.0007419000000000001 3.3 0.000742 0 0.0007419200000000001 0 0.00074202 3.3 0.0007419400000000001 3.3 0.00074204 0 0.0007419600000000001 0 0.00074206 3.3 0.00074198 3.3 0.00074208 0 0.000742 0 0.0007421 3.3 0.00074202 3.3 0.00074212 0 0.00074204 0 0.00074214 3.3 0.00074206 3.3 0.00074216 0 0.00074208 0 0.0007421799999999999 3.3 0.0007421 3.3 0.0007421999999999999 0 0.0007421200000000001 0 0.00074222 3.3 0.0007421400000000001 3.3 0.00074224 0 0.0007421600000000001 0 0.00074226 3.3 0.00074218 3.3 0.00074228 0 0.0007422 0 0.0007423 3.3 0.00074222 3.3 0.00074232 0 0.00074224 0 0.00074234 3.3 0.00074226 3.3 0.00074236 0 0.00074228 0 0.00074238 3.3 0.0007423 3.3 0.0007423999999999999 0 0.0007423200000000001 0 0.00074242 3.3 0.0007423400000000001 3.3 0.00074244 0 0.0007423600000000001 0 0.00074246 3.3 0.0007423800000000001 3.3 0.00074248 0 0.0007424 0 0.0007425 3.3 0.00074242 3.3 0.00074252 0 0.00074244 0 0.00074254 3.3 0.00074246 3.3 0.00074256 0 0.00074248 0 0.00074258 3.3 0.0007425 3.3 0.0007425999999999999 0 0.00074252 0 0.0007426199999999999 3.3 0.0007425400000000001 3.3 0.00074264 0 0.0007425600000000001 0 0.00074266 3.3 0.0007425800000000001 3.3 0.00074268 0 0.0007426 0 0.0007427 3.3 0.00074262 3.3 0.00074272 0 0.00074264 0 0.00074274 3.3 0.00074266 3.3 0.00074276 0 0.00074268 0 0.00074278 3.3 0.0007427 3.3 0.0007428 0 0.00074272 0 0.0007428199999999999 3.3 0.0007427400000000001 3.3 0.00074284 0 0.0007427600000000001 0 0.00074286 3.3 0.0007427800000000001 3.3 0.00074288 0 0.0007428000000000001 0 0.0007429 3.3 0.00074282 3.3 0.00074292 0 0.00074284 0 0.00074294 3.3 0.00074286 3.3 0.00074296 0 0.00074288 0 0.00074298 3.3 0.0007429 3.3 0.000743 0 0.00074292 0 0.0007430199999999999 3.3 0.00074294 3.3 0.0007430399999999999 0 0.0007429600000000001 0 0.00074306 3.3 0.0007429800000000001 3.3 0.00074308 0 0.0007430000000000001 0 0.0007431 3.3 0.00074302 3.3 0.00074312 0 0.00074304 0 0.00074314 3.3 0.00074306 3.3 0.00074316 0 0.00074308 0 0.00074318 3.3 0.0007431 3.3 0.0007432 0 0.00074312 0 0.00074322 3.3 0.00074314 3.3 0.0007432399999999999 0 0.0007431600000000001 0 0.00074326 3.3 0.0007431800000000001 3.3 0.00074328 0 0.0007432000000000001 0 0.0007433 3.3 0.0007432200000000001 3.3 0.00074332 0 0.00074324 0 0.00074334 3.3 0.00074326 3.3 0.00074336 0 0.00074328 0 0.00074338 3.3 0.0007433 3.3 0.0007434 0 0.00074332 0 0.00074342 3.3 0.00074334 3.3 0.0007434399999999999 0 0.00074336 0 0.0007434599999999999 3.3 0.0007433800000000001 3.3 0.00074348 0 0.0007434000000000001 0 0.0007435 3.3 0.0007434200000000001 3.3 0.00074352 0 0.00074344 0 0.00074354 3.3 0.00074346 3.3 0.00074356 0 0.00074348 0 0.00074358 3.3 0.0007435 3.3 0.0007436 0 0.00074352 0 0.00074362 3.3 0.00074354 3.3 0.00074364 0 0.00074356 0 0.0007436599999999999 3.3 0.0007435800000000001 3.3 0.00074368 0 0.0007436000000000001 0 0.0007437 3.3 0.0007436200000000001 3.3 0.00074372 0 0.0007436400000000001 0 0.00074374 3.3 0.00074366 3.3 0.00074376 0 0.00074368 0 0.00074378 3.3 0.0007437 3.3 0.0007438 0 0.00074372 0 0.00074382 3.3 0.00074374 3.3 0.00074384 0 0.00074376 0 0.0007438599999999999 3.3 0.00074378 3.3 0.0007438799999999999 0 0.0007438000000000001 0 0.0007439 3.3 0.0007438200000000001 3.3 0.00074392 0 0.0007438400000000001 0 0.00074394 3.3 0.00074386 3.3 0.00074396 0 0.00074388 0 0.00074398 3.3 0.0007439 3.3 0.000744 0 0.00074392 0 0.00074402 3.3 0.00074394 3.3 0.00074404 0 0.00074396 0 0.00074406 3.3 0.00074398 3.3 0.0007440799999999999 0 0.0007440000000000001 0 0.0007441 3.3 0.0007440200000000001 3.3 0.00074412 0 0.0007440400000000001 0 0.00074414 3.3 0.0007440600000000001 3.3 0.00074416 0 0.00074408 0 0.00074418 3.3 0.0007441 3.3 0.0007442 0 0.00074412 0 0.00074422 3.3 0.00074414 3.3 0.00074424 0 0.00074416 0 0.00074426 3.3 0.00074418 3.3 0.0007442799999999999 0 0.0007442 0 0.0007442999999999999 3.3 0.0007442200000000001 3.3 0.00074432 0 0.0007442400000000001 0 0.00074434 3.3 0.0007442600000000001 3.3 0.00074436 0 0.00074428 0 0.00074438 3.3 0.0007443 3.3 0.0007444 0 0.00074432 0 0.00074442 3.3 0.00074434 3.3 0.00074444 0 0.00074436 0 0.00074446 3.3 0.00074438 3.3 0.00074448 0 0.0007444 0 0.0007444999999999999 3.3 0.0007444200000000001 3.3 0.00074452 0 0.0007444400000000001 0 0.00074454 3.3 0.0007444600000000001 3.3 0.00074456 0 0.0007444800000000001 0 0.00074458 3.3 0.0007445 3.3 0.0007446 0 0.00074452 0 0.00074462 3.3 0.00074454 3.3 0.00074464 0 0.00074456 0 0.00074466 3.3 0.00074458 3.3 0.00074468 0 0.0007446 0 0.0007446999999999999 3.3 0.0007446200000000001 3.3 0.00074472 0 0.0007446400000000001 0 0.00074474 3.3 0.0007446600000000001 3.3 0.00074476 0 0.0007446800000000001 0 0.00074478 3.3 0.0007447 3.3 0.0007448 0 0.00074472 0 0.00074482 3.3 0.00074474 3.3 0.00074484 0 0.00074476 0 0.00074486 3.3 0.00074478 3.3 0.00074488 0 0.0007448 0 0.0007449 3.3 0.00074482 3.3 0.0007449199999999999 0 0.0007448400000000001 0 0.00074494 3.3 0.0007448600000000001 3.3 0.00074496 0 0.0007448800000000001 0 0.00074498 3.3 0.0007449000000000001 3.3 0.000745 0 0.00074492 0 0.00074502 3.3 0.00074494 3.3 0.00074504 0 0.00074496 0 0.00074506 3.3 0.00074498 3.3 0.00074508 0 0.000745 0 0.0007451 3.3 0.00074502 3.3 0.0007451199999999999 0 0.0007450400000000001 0 0.00074514 3.3 0.0007450600000000001 3.3 0.00074516 0 0.0007450800000000001 0 0.00074518 3.3 0.0007451000000000001 3.3 0.0007452 0 0.00074512 0 0.00074522 3.3 0.00074514 3.3 0.00074524 0 0.00074516 0 0.00074526 3.3 0.00074518 3.3 0.00074528 0 0.0007452 0 0.0007453 3.3 0.00074522 3.3 0.0007453199999999999 0 0.00074524 0 0.0007453399999999999 3.3 0.0007452600000000001 3.3 0.00074536 0 0.0007452800000000001 0 0.00074538 3.3 0.0007453000000000001 3.3 0.0007454 0 0.00074532 0 0.00074542 3.3 0.00074534 3.3 0.00074544 0 0.00074536 0 0.00074546 3.3 0.00074538 3.3 0.00074548 0 0.0007454 0 0.0007455 3.3 0.00074542 3.3 0.00074552 0 0.00074544 0 0.0007455399999999999 3.3 0.0007454600000000001 3.3 0.00074556 0 0.0007454800000000001 0 0.00074558 3.3 0.0007455000000000001 3.3 0.0007456 0 0.0007455200000000001 0 0.00074562 3.3 0.00074554 3.3 0.00074564 0 0.00074556 0 0.00074566 3.3 0.00074558 3.3 0.00074568 0 0.0007456 0 0.0007457 3.3 0.00074562 3.3 0.00074572 0 0.00074564 0 0.0007457399999999999 3.3 0.00074566 3.3 0.0007457599999999999 0 0.0007456800000000001 0 0.00074578 3.3 0.0007457000000000001 3.3 0.0007458 0 0.0007457200000000001 0 0.00074582 3.3 0.00074574 3.3 0.00074584 0 0.00074576 0 0.00074586 3.3 0.00074578 3.3 0.00074588 0 0.0007458 0 0.0007459 3.3 0.00074582 3.3 0.00074592 0 0.00074584 0 0.00074594 3.3 0.00074586 3.3 0.0007459599999999999 0 0.0007458800000000001 0 0.00074598 3.3 0.0007459000000000001 3.3 0.000746 0 0.0007459200000000001 0 0.00074602 3.3 0.0007459400000000001 3.3 0.00074604 0 0.00074596 0 0.00074606 3.3 0.00074598 3.3 0.00074608 0 0.000746 0 0.0007461 3.3 0.00074602 3.3 0.00074612 0 0.00074604 0 0.00074614 3.3 0.00074606 3.3 0.0007461599999999999 0 0.00074608 0 0.0007461799999999999 3.3 0.0007461000000000001 3.3 0.0007462 0 0.0007461200000000001 0 0.00074622 3.3 0.0007461400000000001 3.3 0.00074624 0 0.00074616 0 0.00074626 3.3 0.00074618 3.3 0.00074628 0 0.0007462 0 0.0007463 3.3 0.00074622 3.3 0.00074632 0 0.00074624 0 0.00074634 3.3 0.00074626 3.3 0.00074636 0 0.00074628 0 0.0007463799999999999 3.3 0.0007463000000000001 3.3 0.0007464 0 0.0007463200000000001 0 0.00074642 3.3 0.0007463400000000001 3.3 0.00074644 0 0.0007463600000000001 0 0.00074646 3.3 0.00074638 3.3 0.00074648 0 0.0007464 0 0.0007465 3.3 0.00074642 3.3 0.00074652 0 0.00074644 0 0.00074654 3.3 0.00074646 3.3 0.00074656 0 0.00074648 0 0.0007465799999999999 3.3 0.0007465 3.3 0.0007465999999999999 0 0.0007465200000000001 0 0.00074662 3.3 0.0007465400000000001 3.3 0.00074664 0 0.0007465600000000001 0 0.00074666 3.3 0.00074658 3.3 0.00074668 0 0.0007466 0 0.0007467 3.3 0.00074662 3.3 0.00074672 0 0.00074664 0 0.00074674 3.3 0.00074666 3.3 0.00074676 0 0.00074668 0 0.00074678 3.3 0.0007467 3.3 0.0007467999999999999 0 0.0007467200000000001 0 0.00074682 3.3 0.0007467400000000001 3.3 0.00074684 0 0.0007467600000000001 0 0.00074686 3.3 0.0007467800000000001 3.3 0.00074688 0 0.0007468 0 0.0007469 3.3 0.00074682 3.3 0.00074692 0 0.00074684 0 0.00074694 3.3 0.00074686 3.3 0.00074696 0 0.00074688 0 0.00074698 3.3 0.0007469 3.3 0.0007469999999999999 0 0.00074692 0 0.0007470199999999999 3.3 0.0007469400000000001 3.3 0.00074704 0 0.0007469600000000001 0 0.00074706 3.3 0.0007469800000000001 3.3 0.00074708 0 0.000747 0 0.0007471 3.3 0.00074702 3.3 0.00074712 0 0.00074704 0 0.00074714 3.3 0.00074706 3.3 0.00074716 0 0.00074708 0 0.00074718 3.3 0.0007471 3.3 0.0007472 0 0.00074712 0 0.0007472199999999999 3.3 0.0007471400000000001 3.3 0.00074724 0 0.0007471600000000001 0 0.00074726 3.3 0.0007471800000000001 3.3 0.00074728 0 0.0007472000000000001 0 0.0007473 3.3 0.00074722 3.3 0.00074732 0 0.00074724 0 0.00074734 3.3 0.00074726 3.3 0.00074736 0 0.00074728 0 0.00074738 3.3 0.0007473 3.3 0.0007474 0 0.00074732 0 0.0007474199999999999 3.3 0.00074734 3.3 0.0007474399999999999 0 0.0007473600000000001 0 0.00074746 3.3 0.0007473800000000001 3.3 0.00074748 0 0.0007474000000000001 0 0.0007475 3.3 0.00074742 3.3 0.00074752 0 0.00074744 0 0.00074754 3.3 0.00074746 3.3 0.00074756 0 0.00074748 0 0.00074758 3.3 0.0007475 3.3 0.0007476 0 0.00074752 0 0.00074762 3.3 0.00074754 3.3 0.0007476399999999999 0 0.0007475600000000001 0 0.00074766 3.3 0.0007475800000000001 3.3 0.00074768 0 0.0007476000000000001 0 0.0007477 3.3 0.0007476200000000001 3.3 0.00074772 0 0.00074764 0 0.00074774 3.3 0.00074766 3.3 0.00074776 0 0.00074768 0 0.00074778 3.3 0.0007477 3.3 0.0007478 0 0.00074772 0 0.00074782 3.3 0.00074774 3.3 0.0007478399999999999 0 0.00074776 0 0.0007478599999999999 3.3 0.0007477800000000001 3.3 0.00074788 0 0.0007478000000000001 0 0.0007479 3.3 0.0007478200000000001 3.3 0.00074792 0 0.00074784 0 0.00074794 3.3 0.00074786 3.3 0.00074796 0 0.00074788 0 0.00074798 3.3 0.0007479 3.3 0.000748 0 0.00074792 0 0.00074802 3.3 0.00074794 3.3 0.00074804 0 0.00074796 0 0.0007480599999999999 3.3 0.0007479800000000001 3.3 0.00074808 0 0.0007480000000000001 0 0.0007481 3.3 0.0007480200000000001 3.3 0.00074812 0 0.0007480400000000001 0 0.00074814 3.3 0.00074806 3.3 0.00074816 0 0.00074808 0 0.00074818 3.3 0.0007481 3.3 0.0007482 0 0.00074812 0 0.00074822 3.3 0.00074814 3.3 0.00074824 0 0.00074816 0 0.0007482599999999999 3.3 0.0007481800000000001 3.3 0.00074828 0 0.0007482000000000001 0 0.0007483 3.3 0.0007482200000000001 3.3 0.00074832 0 0.0007482400000000001 0 0.00074834 3.3 0.00074826 3.3 0.00074836 0 0.00074828 0 0.00074838 3.3 0.0007483 3.3 0.0007484 0 0.00074832 0 0.00074842 3.3 0.00074834 3.3 0.00074844 0 0.00074836 0 0.0007484599999999999 3.3 0.00074838 3.3 0.0007484799999999999 0 0.0007484000000000001 0 0.0007485 3.3 0.0007484200000000001 3.3 0.00074852 0 0.0007484400000000001 0 0.00074854 3.3 0.00074846 3.3 0.00074856 0 0.00074848 0 0.00074858 3.3 0.0007485 3.3 0.0007486 0 0.00074852 0 0.00074862 3.3 0.00074854 3.3 0.00074864 0 0.00074856 0 0.00074866 3.3 0.00074858 3.3 0.0007486799999999999 0 0.0007486000000000001 0 0.0007487 3.3 0.0007486200000000001 3.3 0.00074872 0 0.0007486400000000001 0 0.00074874 3.3 0.0007486600000000001 3.3 0.00074876 0 0.00074868 0 0.00074878 3.3 0.0007487 3.3 0.0007488 0 0.00074872 0 0.00074882 3.3 0.00074874 3.3 0.00074884 0 0.00074876 0 0.00074886 3.3 0.00074878 3.3 0.0007488799999999999 0 0.0007488 0 0.0007488999999999999 3.3 0.0007488200000000001 3.3 0.00074892 0 0.0007488400000000001 0 0.00074894 3.3 0.0007488600000000001 3.3 0.00074896 0 0.00074888 0 0.00074898 3.3 0.0007489 3.3 0.000749 0 0.00074892 0 0.00074902 3.3 0.00074894 3.3 0.00074904 0 0.00074896 0 0.00074906 3.3 0.00074898 3.3 0.00074908 0 0.000749 0 0.0007490999999999999 3.3 0.0007490200000000001 3.3 0.00074912 0 0.0007490400000000001 0 0.00074914 3.3 0.0007490600000000001 3.3 0.00074916 0 0.0007490800000000001 0 0.00074918 3.3 0.0007491 3.3 0.0007492 0 0.00074912 0 0.00074922 3.3 0.00074914 3.3 0.00074924 0 0.00074916 0 0.00074926 3.3 0.00074918 3.3 0.00074928 0 0.0007492 0 0.0007492999999999999 3.3 0.00074922 3.3 0.0007493199999999999 0 0.0007492400000000001 0 0.00074934 3.3 0.0007492600000000001 3.3 0.00074936 0 0.0007492800000000001 0 0.00074938 3.3 0.0007493 3.3 0.0007494 0 0.00074932 0 0.00074942 3.3 0.00074934 3.3 0.00074944 0 0.00074936 0 0.00074946 3.3 0.00074938 3.3 0.00074948 0 0.0007494 0 0.0007495 3.3 0.00074942 3.3 0.0007495199999999999 0 0.0007494400000000001 0 0.00074954 3.3 0.0007494600000000001 3.3 0.00074956 0 0.0007494800000000001 0 0.00074958 3.3 0.0007495000000000001 3.3 0.0007496 0 0.00074952 0 0.00074962 3.3 0.00074954 3.3 0.00074964 0 0.00074956 0 0.00074966 3.3 0.00074958 3.3 0.00074968 0 0.0007496 0 0.0007497 3.3 0.00074962 3.3 0.0007497199999999999 0 0.00074964 0 0.0007497399999999999 3.3 0.0007496600000000001 3.3 0.00074976 0 0.0007496800000000001 0 0.00074978 3.3 0.0007497000000000001 3.3 0.0007498 0 0.00074972 0 0.00074982 3.3 0.00074974 3.3 0.00074984 0 0.00074976 0 0.00074986 3.3 0.00074978 3.3 0.00074988 0 0.0007498 0 0.0007499 3.3 0.00074982 3.3 0.00074992 0 0.00074984 0 0.0007499399999999999 3.3 0.0007498600000000001 3.3 0.00074996 0 0.0007498800000000001 0 0.00074998 3.3 0.0007499000000000001 3.3 0.00075 0 0.0007499200000000001 0 0.00075002 3.3 0.00074994 3.3 0.00075004 0 0.00074996 0 0.00075006 3.3 0.00074998 3.3 0.00075008 0 0.00075 0 0.0007501 3.3 0.00075002 3.3 0.00075012 0 0.00075004 0 0.0007501399999999999 3.3 0.00075006 3.3 0.0007501599999999999 0 0.0007500800000000001 0 0.00075018 3.3 0.0007501000000000001 3.3 0.0007502 0 0.0007501200000000001 0 0.00075022 3.3 0.00075014 3.3 0.00075024 0 0.00075016 0 0.00075026 3.3 0.00075018 3.3 0.00075028 0 0.0007502 0 0.0007503 3.3 0.00075022 3.3 0.00075032 0 0.00075024 0 0.00075034 3.3 0.00075026 3.3 0.0007503599999999999 0 0.0007502800000000001 0 0.00075038 3.3 0.0007503000000000001 3.3 0.0007504 0 0.0007503200000000001 0 0.00075042 3.3 0.0007503400000000001 3.3 0.00075044 0 0.00075036 0 0.00075046 3.3 0.00075038 3.3 0.00075048 0 0.0007504 0 0.0007505 3.3 0.00075042 3.3 0.00075052 0 0.00075044 0 0.00075054 3.3 0.00075046 3.3 0.0007505599999999999 0 0.00075048 0 0.0007505799999999999 3.3 0.0007505000000000001 3.3 0.0007506 0 0.0007505200000000001 0 0.00075062 3.3 0.0007505400000000001 3.3 0.00075064 0 0.00075056 0 0.00075066 3.3 0.00075058 3.3 0.00075068 0 0.0007506 0 0.0007507 3.3 0.00075062 3.3 0.00075072 0 0.00075064 0 0.00075074 3.3 0.00075066 3.3 0.00075076 0 0.00075068 0 0.0007507799999999999 3.3 0.0007507000000000001 3.3 0.0007508 0 0.0007507200000000001 0 0.00075082 3.3 0.0007507400000000001 3.3 0.00075084 0 0.0007507600000000001 0 0.00075086 3.3 0.00075078 3.3 0.00075088 0 0.0007508 0 0.0007509 3.3 0.00075082 3.3 0.00075092 0 0.00075084 0 0.00075094 3.3 0.00075086 3.3 0.00075096 0 0.00075088 0 0.0007509799999999999 3.3 0.0007509 3.3 0.0007509999999999999 0 0.0007509200000000001 0 0.00075102 3.3 0.0007509400000000001 3.3 0.00075104 0 0.0007509600000000001 0 0.00075106 3.3 0.00075098 3.3 0.00075108 0 0.000751 0 0.0007511 3.3 0.00075102 3.3 0.00075112 0 0.00075104 0 0.00075114 3.3 0.00075106 3.3 0.00075116 0 0.00075108 0 0.00075118 3.3 0.0007511 3.3 0.0007511999999999999 0 0.0007511200000000001 0 0.00075122 3.3 0.0007511400000000001 3.3 0.00075124 0 0.0007511600000000001 0 0.00075126 3.3 0.0007511800000000001 3.3 0.00075128 0 0.0007512 0 0.0007513 3.3 0.00075122 3.3 0.00075132 0 0.00075124 0 0.00075134 3.3 0.00075126 3.3 0.00075136 0 0.00075128 0 0.00075138 3.3 0.0007513 3.3 0.0007513999999999999 0 0.00075132 0 0.0007514199999999999 3.3 0.0007513400000000001 3.3 0.00075144 0 0.0007513600000000001 0 0.00075146 3.3 0.0007513800000000001 3.3 0.00075148 0 0.0007514 0 0.0007515 3.3 0.00075142 3.3 0.00075152 0 0.00075144 0 0.00075154 3.3 0.00075146 3.3 0.00075156 0 0.00075148 0 0.00075158 3.3 0.0007515 3.3 0.0007516 0 0.00075152 0 0.0007516199999999999 3.3 0.0007515400000000001 3.3 0.00075164 0 0.0007515600000000001 0 0.00075166 3.3 0.0007515800000000001 3.3 0.00075168 0 0.0007516000000000001 0 0.0007517 3.3 0.00075162 3.3 0.00075172 0 0.00075164 0 0.00075174 3.3 0.00075166 3.3 0.00075176 0 0.00075168 0 0.00075178 3.3 0.0007517 3.3 0.0007518 0 0.00075172 0 0.0007518199999999999 3.3 0.0007517400000000001 3.3 0.00075184 0 0.0007517600000000001 0 0.00075186 3.3 0.0007517800000000001 3.3 0.00075188 0 0.0007518000000000001 0 0.0007519 3.3 0.00075182 3.3 0.00075192 0 0.00075184 0 0.00075194 3.3 0.00075186 3.3 0.00075196 0 0.00075188 0 0.00075198 3.3 0.0007519 3.3 0.000752 0 0.00075192 0 0.0007520199999999999 3.3 0.00075194 3.3 0.0007520399999999999 0 0.0007519600000000001 0 0.00075206 3.3 0.0007519800000000001 3.3 0.00075208 0 0.0007520000000000001 0 0.0007521 3.3 0.00075202 3.3 0.00075212 0 0.00075204 0 0.00075214 3.3 0.00075206 3.3 0.00075216 0 0.00075208 0 0.00075218 3.3 0.0007521 3.3 0.0007522 0 0.00075212 0 0.00075222 3.3 0.00075214 3.3 0.0007522399999999999 0 0.0007521600000000001 0 0.00075226 3.3 0.0007521800000000001 3.3 0.00075228 0 0.0007522000000000001 0 0.0007523 3.3 0.0007522200000000001 3.3 0.00075232 0 0.00075224 0 0.00075234 3.3 0.00075226 3.3 0.00075236 0 0.00075228 0 0.00075238 3.3 0.0007523 3.3 0.0007524 0 0.00075232 0 0.00075242 3.3 0.00075234 3.3 0.0007524399999999999 0 0.00075236 0 0.0007524599999999999 3.3 0.0007523800000000001 3.3 0.00075248 0 0.0007524000000000001 0 0.0007525 3.3 0.0007524200000000001 3.3 0.00075252 0 0.00075244 0 0.00075254 3.3 0.00075246 3.3 0.00075256 0 0.00075248 0 0.00075258 3.3 0.0007525 3.3 0.0007526 0 0.00075252 0 0.00075262 3.3 0.00075254 3.3 0.00075264 0 0.00075256 0 0.0007526599999999999 3.3 0.0007525800000000001 3.3 0.00075268 0 0.0007526000000000001 0 0.0007527 3.3 0.0007526200000000001 3.3 0.00075272 0 0.0007526400000000001 0 0.00075274 3.3 0.00075266 3.3 0.00075276 0 0.00075268 0 0.00075278 3.3 0.0007527 3.3 0.0007528 0 0.00075272 0 0.00075282 3.3 0.00075274 3.3 0.00075284 0 0.00075276 0 0.0007528599999999999 3.3 0.00075278 3.3 0.0007528799999999999 0 0.0007528000000000001 0 0.0007529 3.3 0.0007528200000000001 3.3 0.00075292 0 0.0007528400000000001 0 0.00075294 3.3 0.00075286 3.3 0.00075296 0 0.00075288 0 0.00075298 3.3 0.0007529 3.3 0.000753 0 0.00075292 0 0.00075302 3.3 0.00075294 3.3 0.00075304 0 0.00075296 0 0.00075306 3.3 0.00075298 3.3 0.0007530799999999999 0 0.0007530000000000001 0 0.0007531 3.3 0.0007530200000000001 3.3 0.00075312 0 0.0007530400000000001 0 0.00075314 3.3 0.0007530600000000001 3.3 0.00075316 0 0.00075308 0 0.00075318 3.3 0.0007531 3.3 0.0007532 0 0.00075312 0 0.00075322 3.3 0.00075314 3.3 0.00075324 0 0.00075316 0 0.00075326 3.3 0.00075318 3.3 0.0007532799999999999 0 0.0007532 0 0.0007532999999999999 3.3 0.0007532200000000001 3.3 0.00075332 0 0.0007532400000000001 0 0.00075334 3.3 0.0007532600000000001 3.3 0.00075336 0 0.00075328 0 0.00075338 3.3 0.0007533 3.3 0.0007534 0 0.00075332 0 0.00075342 3.3 0.00075334 3.3 0.00075344 0 0.00075336 0 0.00075346 3.3 0.00075338 3.3 0.00075348 0 0.0007534 0 0.0007534999999999999 3.3 0.0007534200000000001 3.3 0.00075352 0 0.0007534400000000001 0 0.00075354 3.3 0.0007534600000000001 3.3 0.00075356 0 0.0007534800000000001 0 0.00075358 3.3 0.0007535 3.3 0.0007536 0 0.00075352 0 0.00075362 3.3 0.00075354 3.3 0.00075364 0 0.00075356 0 0.00075366 3.3 0.00075358 3.3 0.00075368 0 0.0007536 0 0.0007536999999999999 3.3 0.00075362 3.3 0.0007537199999999999 0 0.0007536400000000001 0 0.00075374 3.3 0.0007536600000000001 3.3 0.00075376 0 0.0007536800000000001 0 0.00075378 3.3 0.0007537 3.3 0.0007538 0 0.00075372 0 0.00075382 3.3 0.00075374 3.3 0.00075384 0 0.00075376 0 0.00075386 3.3 0.00075378 3.3 0.00075388 0 0.0007538 0 0.0007539 3.3 0.00075382 3.3 0.0007539199999999999 0 0.0007538400000000001 0 0.00075394 3.3 0.0007538600000000001 3.3 0.00075396 0 0.0007538800000000001 0 0.00075398 3.3 0.0007539000000000001 3.3 0.000754 0 0.00075392 0 0.00075402 3.3 0.00075394 3.3 0.00075404 0 0.00075396 0 0.00075406 3.3 0.00075398 3.3 0.00075408 0 0.000754 0 0.0007541 3.3 0.00075402 3.3 0.0007541199999999999 0 0.00075404 0 0.0007541399999999999 3.3 0.0007540600000000001 3.3 0.00075416 0 0.0007540800000000001 0 0.00075418 3.3 0.0007541000000000001 3.3 0.0007542 0 0.00075412 0 0.00075422 3.3 0.00075414 3.3 0.00075424 0 0.00075416 0 0.00075426 3.3 0.00075418 3.3 0.00075428 0 0.0007542 0 0.0007543 3.3 0.00075422 3.3 0.00075432 0 0.00075424 0 0.0007543399999999999 3.3 0.0007542600000000001 3.3 0.00075436 0 0.0007542800000000001 0 0.00075438 3.3 0.0007543000000000001 3.3 0.0007544 0 0.0007543200000000001 0 0.00075442 3.3 0.00075434 3.3 0.00075444 0 0.00075436 0 0.00075446 3.3 0.00075438 3.3 0.00075448 0 0.0007544 0 0.0007545 3.3 0.00075442 3.3 0.00075452 0 0.00075444 0 0.0007545399999999999 3.3 0.00075446 3.3 0.0007545599999999999 0 0.0007544800000000001 0 0.00075458 3.3 0.0007545000000000001 3.3 0.0007546 0 0.0007545200000000001 0 0.00075462 3.3 0.00075454 3.3 0.00075464 0 0.00075456 0 0.00075466 3.3 0.00075458 3.3 0.00075468 0 0.0007546 0 0.0007547 3.3 0.00075462 3.3 0.00075472 0 0.00075464 0 0.00075474 3.3 0.00075466 3.3 0.0007547599999999999 0 0.0007546800000000001 0 0.00075478 3.3 0.0007547000000000001 3.3 0.0007548 0 0.0007547200000000001 0 0.00075482 3.3 0.0007547400000000001 3.3 0.00075484 0 0.00075476 0 0.00075486 3.3 0.00075478 3.3 0.00075488 0 0.0007548 0 0.0007549 3.3 0.00075482 3.3 0.00075492 0 0.00075484 0 0.00075494 3.3 0.00075486 3.3 0.0007549599999999999 0 0.00075488 0 0.0007549799999999999 3.3 0.0007549000000000001 3.3 0.000755 0 0.0007549200000000001 0 0.00075502 3.3 0.0007549400000000001 3.3 0.00075504 0 0.00075496 0 0.00075506 3.3 0.00075498 3.3 0.00075508 0 0.000755 0 0.0007551 3.3 0.00075502 3.3 0.00075512 0 0.00075504 0 0.00075514 3.3 0.00075506 3.3 0.00075516 0 0.00075508 0 0.0007551799999999999 3.3 0.0007551000000000001 3.3 0.0007552 0 0.0007551200000000001 0 0.00075522 3.3 0.0007551400000000001 3.3 0.00075524 0 0.0007551600000000001 0 0.00075526 3.3 0.00075518 3.3 0.00075528 0 0.0007552 0 0.0007553 3.3 0.00075522 3.3 0.00075532 0 0.00075524 0 0.00075534 3.3 0.00075526 3.3 0.00075536 0 0.00075528 0 0.0007553799999999999 3.3 0.0007553000000000001 3.3 0.0007554 0 0.0007553200000000001 0 0.00075542 3.3 0.0007553400000000001 3.3 0.00075544 0 0.0007553600000000001 0 0.00075546 3.3 0.00075538 3.3 0.00075548 0 0.0007554 0 0.0007555 3.3 0.00075542 3.3 0.00075552 0 0.00075544 0 0.00075554 3.3 0.00075546 3.3 0.00075556 0 0.00075548 0 0.0007555799999999999 3.3 0.0007555 3.3 0.0007555999999999999 0 0.0007555200000000001 0 0.00075562 3.3 0.0007555400000000001 3.3 0.00075564 0 0.0007555600000000001 0 0.00075566 3.3 0.00075558 3.3 0.00075568 0 0.0007556 0 0.0007557 3.3 0.00075562 3.3 0.00075572 0 0.00075564 0 0.00075574 3.3 0.00075566 3.3 0.00075576 0 0.00075568 0 0.00075578 3.3 0.0007557 3.3 0.0007557999999999999 0 0.0007557200000000001 0 0.00075582 3.3 0.0007557400000000001 3.3 0.00075584 0 0.0007557600000000001 0 0.00075586 3.3 0.0007557800000000001 3.3 0.00075588 0 0.0007558 0 0.0007559 3.3 0.00075582 3.3 0.00075592 0 0.00075584 0 0.00075594 3.3 0.00075586 3.3 0.00075596 0 0.00075588 0 0.00075598 3.3 0.0007559 3.3 0.0007559999999999999 0 0.00075592 0 0.0007560199999999999 3.3 0.0007559400000000001 3.3 0.00075604 0 0.0007559600000000001 0 0.00075606 3.3 0.0007559800000000001 3.3 0.00075608 0 0.000756 0 0.0007561 3.3 0.00075602 3.3 0.00075612 0 0.00075604 0 0.00075614 3.3 0.00075606 3.3 0.00075616 0 0.00075608 0 0.00075618 3.3 0.0007561 3.3 0.0007562 0 0.00075612 0 0.0007562199999999999 3.3 0.0007561400000000001 3.3 0.00075624 0 0.0007561600000000001 0 0.00075626 3.3 0.0007561800000000001 3.3 0.00075628 0 0.0007562000000000001 0 0.0007563 3.3 0.00075622 3.3 0.00075632 0 0.00075624 0 0.00075634 3.3 0.00075626 3.3 0.00075636 0 0.00075628 0 0.00075638 3.3 0.0007563 3.3 0.0007564 0 0.00075632 0 0.0007564199999999999 3.3 0.00075634 3.3 0.0007564399999999999 0 0.0007563600000000001 0 0.00075646 3.3 0.0007563800000000001 3.3 0.00075648 0 0.0007564000000000001 0 0.0007565 3.3 0.00075642 3.3 0.00075652 0 0.00075644 0 0.00075654 3.3 0.00075646 3.3 0.00075656 0 0.00075648 0 0.00075658 3.3 0.0007565 3.3 0.0007566 0 0.00075652 0 0.00075662 3.3 0.00075654 3.3 0.0007566399999999999 0 0.0007565600000000001 0 0.00075666 3.3 0.0007565800000000001 3.3 0.00075668 0 0.0007566000000000001 0 0.0007567 3.3 0.0007566200000000001 3.3 0.00075672 0 0.00075664 0 0.00075674 3.3 0.00075666 3.3 0.00075676 0 0.00075668 0 0.00075678 3.3 0.0007567 3.3 0.0007568 0 0.00075672 0 0.00075682 3.3 0.00075674 3.3 0.0007568399999999999 0 0.00075676 0 0.0007568599999999999 3.3 0.0007567800000000001 3.3 0.00075688 0 0.0007568000000000001 0 0.0007569 3.3 0.0007568200000000001 3.3 0.00075692 0 0.00075684 0 0.00075694 3.3 0.00075686 3.3 0.00075696 0 0.00075688 0 0.00075698 3.3 0.0007569 3.3 0.000757 0 0.00075692 0 0.00075702 3.3 0.00075694 3.3 0.00075704 0 0.00075696 0 0.0007570599999999999 3.3 0.0007569800000000001 3.3 0.00075708 0 0.0007570000000000001 0 0.0007571 3.3 0.0007570200000000001 3.3 0.00075712 0 0.0007570400000000001 0 0.00075714 3.3 0.00075706 3.3 0.00075716 0 0.00075708 0 0.00075718 3.3 0.0007571 3.3 0.0007572 0 0.00075712 0 0.00075722 3.3 0.00075714 3.3 0.00075724 0 0.00075716 0 0.0007572599999999999 3.3 0.00075718 3.3 0.0007572799999999999 0 0.0007572000000000001 0 0.0007573 3.3 0.0007572200000000001 3.3 0.00075732 0 0.0007572400000000001 0 0.00075734 3.3 0.00075726 3.3 0.00075736 0 0.00075728 0 0.00075738 3.3 0.0007573 3.3 0.0007574 0 0.00075732 0 0.00075742 3.3 0.00075734 3.3 0.00075744 0 0.00075736 0 0.00075746 3.3 0.00075738 3.3 0.0007574799999999999 0 0.0007574000000000001 0 0.0007575 3.3 0.0007574200000000001 3.3 0.00075752 0 0.0007574400000000001 0 0.00075754 3.3 0.0007574600000000001 3.3 0.00075756 0 0.00075748 0 0.00075758 3.3 0.0007575 3.3 0.0007576 0 0.00075752 0 0.00075762 3.3 0.00075754 3.3 0.00075764 0 0.00075756 0 0.00075766 3.3 0.00075758 3.3 0.0007576799999999999 0 0.0007576 0 0.0007576999999999999 3.3 0.0007576200000000001 3.3 0.00075772 0 0.0007576400000000001 0 0.00075774 3.3 0.0007576600000000001 3.3 0.00075776 0 0.00075768 0 0.00075778 3.3 0.0007577 3.3 0.0007578 0 0.00075772 0 0.00075782 3.3 0.00075774 3.3 0.00075784 0 0.00075776 0 0.00075786 3.3 0.00075778 3.3 0.00075788 0 0.0007578 0 0.0007578999999999999 3.3 0.0007578200000000001 3.3 0.00075792 0 0.0007578400000000001 0 0.00075794 3.3 0.0007578600000000001 3.3 0.00075796 0 0.0007578800000000001 0 0.00075798 3.3 0.0007579 3.3 0.000758 0 0.00075792 0 0.00075802 3.3 0.00075794 3.3 0.00075804 0 0.00075796 0 0.00075806 3.3 0.00075798 3.3 0.00075808 0 0.000758 0 0.0007580999999999999 3.3 0.00075802 3.3 0.0007581199999999999 0 0.0007580400000000001 0 0.00075814 3.3 0.0007580600000000001 3.3 0.00075816 0 0.0007580800000000001 0 0.00075818 3.3 0.0007581 3.3 0.0007582 0 0.00075812 0 0.00075822 3.3 0.00075814 3.3 0.00075824 0 0.00075816 0 0.00075826 3.3 0.00075818 3.3 0.00075828 0 0.0007582 0 0.0007583 3.3 0.00075822 3.3 0.0007583199999999999 0 0.0007582400000000001 0 0.00075834 3.3 0.0007582600000000001 3.3 0.00075836 0 0.0007582800000000001 0 0.00075838 3.3 0.0007583000000000001 3.3 0.0007584 0 0.00075832 0 0.00075842 3.3 0.00075834 3.3 0.00075844 0 0.00075836 0 0.00075846 3.3 0.00075838 3.3 0.00075848 0 0.0007584 0 0.0007585 3.3 0.00075842 3.3 0.0007585199999999999 0 0.0007584400000000001 0 0.00075854 3.3 0.0007584600000000001 3.3 0.00075856 0 0.0007584800000000001 0 0.00075858 3.3 0.0007585000000000001 3.3 0.0007586 0 0.00075852 0 0.00075862 3.3 0.00075854 3.3 0.00075864 0 0.00075856 0 0.00075866 3.3 0.00075858 3.3 0.00075868 0 0.0007586 0 0.0007587 3.3 0.00075862 3.3 0.0007587199999999999 0 0.00075864 0 0.0007587399999999999 3.3 0.0007586600000000001 3.3 0.00075876 0 0.0007586800000000001 0 0.00075878 3.3 0.0007587000000000001 3.3 0.0007588 0 0.00075872 0 0.00075882 3.3 0.00075874 3.3 0.00075884 0 0.00075876 0 0.00075886 3.3 0.00075878 3.3 0.00075888 0 0.0007588 0 0.0007589 3.3 0.00075882 3.3 0.00075892 0 0.00075884 0 0.0007589399999999999 3.3 0.0007588600000000001 3.3 0.00075896 0 0.0007588800000000001 0 0.00075898 3.3 0.0007589000000000001 3.3 0.000759 0 0.0007589200000000001 0 0.00075902 3.3 0.00075894 3.3 0.00075904 0 0.00075896 0 0.00075906 3.3 0.00075898 3.3 0.00075908 0 0.000759 0 0.0007591 3.3 0.00075902 3.3 0.00075912 0 0.00075904 0 0.0007591399999999999 3.3 0.00075906 3.3 0.0007591599999999999 0 0.0007590800000000001 0 0.00075918 3.3 0.0007591000000000001 3.3 0.0007592 0 0.0007591200000000001 0 0.00075922 3.3 0.00075914 3.3 0.00075924 0 0.00075916 0 0.00075926 3.3 0.00075918 3.3 0.00075928 0 0.0007592 0 0.0007593 3.3 0.00075922 3.3 0.00075932 0 0.00075924 0 0.00075934 3.3 0.00075926 3.3 0.0007593599999999999 0 0.0007592800000000001 0 0.00075938 3.3 0.0007593000000000001 3.3 0.0007594 0 0.0007593200000000001 0 0.00075942 3.3 0.0007593400000000001 3.3 0.00075944 0 0.00075936 0 0.00075946 3.3 0.00075938 3.3 0.00075948 0 0.0007594 0 0.0007595 3.3 0.00075942 3.3 0.00075952 0 0.00075944 0 0.00075954 3.3 0.00075946 3.3 0.0007595599999999999 0 0.00075948 0 0.0007595799999999999 3.3 0.0007595000000000001 3.3 0.0007596 0 0.0007595200000000001 0 0.00075962 3.3 0.0007595400000000001 3.3 0.00075964 0 0.00075956 0 0.00075966 3.3 0.00075958 3.3 0.00075968 0 0.0007596 0 0.0007597 3.3 0.00075962 3.3 0.00075972 0 0.00075964 0 0.00075974 3.3 0.00075966 3.3 0.00075976 0 0.00075968 0 0.0007597799999999999 3.3 0.0007597000000000001 3.3 0.0007598 0 0.0007597200000000001 0 0.00075982 3.3 0.0007597400000000001 3.3 0.00075984 0 0.0007597600000000001 0 0.00075986 3.3 0.00075978 3.3 0.00075988 0 0.0007598 0 0.0007599 3.3 0.00075982 3.3 0.00075992 0 0.00075984 0 0.00075994 3.3 0.00075986 3.3 0.00075996 0 0.00075988 0 0.0007599799999999999 3.3 0.0007599 3.3 0.0007599999999999999 0 0.0007599200000000001 0 0.00076002 3.3 0.0007599400000000001 3.3 0.00076004 0 0.0007599600000000001 0 0.00076006 3.3 0.00075998 3.3 0.00076008 0 0.00076 0 0.0007601 3.3 0.00076002 3.3 0.00076012 0 0.00076004 0 0.00076014 3.3 0.00076006 3.3 0.00076016 0 0.00076008 0 0.00076018 3.3 0.0007601 3.3 0.0007601999999999999 0 0.0007601200000000001 0 0.00076022 3.3 0.0007601400000000001 3.3 0.00076024 0 0.0007601600000000001 0 0.00076026 3.3 0.0007601800000000001 3.3 0.00076028 0 0.0007602 0 0.0007603 3.3 0.00076022 3.3 0.00076032 0 0.00076024 0 0.00076034 3.3 0.00076026 3.3 0.00076036 0 0.00076028 0 0.00076038 3.3 0.0007603 3.3 0.0007603999999999999 0 0.00076032 0 0.0007604199999999999 3.3 0.0007603400000000001 3.3 0.00076044 0 0.0007603600000000001 0 0.00076046 3.3 0.0007603800000000001 3.3 0.00076048 0 0.0007604 0 0.0007605 3.3 0.00076042 3.3 0.00076052 0 0.00076044 0 0.00076054 3.3 0.00076046 3.3 0.00076056 0 0.00076048 0 0.00076058 3.3 0.0007605 3.3 0.0007606 0 0.00076052 0 0.0007606199999999999 3.3 0.0007605400000000001 3.3 0.00076064 0 0.0007605600000000001 0 0.00076066 3.3 0.0007605800000000001 3.3 0.00076068 0 0.0007606000000000001 0 0.0007607 3.3 0.00076062 3.3 0.00076072 0 0.00076064 0 0.00076074 3.3 0.00076066 3.3 0.00076076 0 0.00076068 0 0.00076078 3.3 0.0007607 3.3 0.0007608 0 0.00076072 0 0.0007608199999999999 3.3 0.00076074 3.3 0.0007608399999999999 0 0.0007607600000000001 0 0.00076086 3.3 0.0007607800000000001 3.3 0.00076088 0 0.0007608000000000001 0 0.0007609 3.3 0.00076082 3.3 0.00076092 0 0.00076084 0 0.00076094 3.3 0.00076086 3.3 0.00076096 0 0.00076088 0 0.00076098 3.3 0.0007609 3.3 0.000761 0 0.00076092 0 0.00076102 3.3 0.00076094 3.3 0.0007610399999999999 0 0.0007609600000000001 0 0.00076106 3.3 0.0007609800000000001 3.3 0.00076108 0 0.0007610000000000001 0 0.0007611 3.3 0.0007610200000000001 3.3 0.00076112 0 0.00076104 0 0.00076114 3.3 0.00076106 3.3 0.00076116 0 0.00076108 0 0.00076118 3.3 0.0007611 3.3 0.0007612 0 0.00076112 0 0.00076122 3.3 0.00076114 3.3 0.0007612399999999999 0 0.00076116 0 0.0007612599999999999 3.3 0.0007611800000000001 3.3 0.00076128 0 0.0007612000000000001 0 0.0007613 3.3 0.0007612200000000001 3.3 0.00076132 0 0.00076124 0 0.00076134 3.3 0.00076126 3.3 0.00076136 0 0.00076128 0 0.00076138 3.3 0.0007613 3.3 0.0007614 0 0.00076132 0 0.00076142 3.3 0.00076134 3.3 0.00076144 0 0.00076136 0 0.0007614599999999999 3.3 0.0007613800000000001 3.3 0.00076148 0 0.0007614000000000001 0 0.0007615 3.3 0.0007614200000000001 3.3 0.00076152 0 0.0007614400000000001 0 0.00076154 3.3 0.00076146 3.3 0.00076156 0 0.00076148 0 0.00076158 3.3 0.0007615 3.3 0.0007616 0 0.00076152 0 0.00076162 3.3 0.00076154 3.3 0.00076164 0 0.00076156 0 0.0007616599999999999 3.3 0.00076158 3.3 0.0007616799999999999 0 0.0007616000000000001 0 0.0007617 3.3 0.0007616200000000001 3.3 0.00076172 0 0.0007616400000000001 0 0.00076174 3.3 0.00076166 3.3 0.00076176 0 0.00076168 0 0.00076178 3.3 0.0007617 3.3 0.0007618 0 0.00076172 0 0.00076182 3.3 0.00076174 3.3 0.00076184 0 0.00076176 0 0.00076186 3.3 0.00076178 3.3 0.0007618799999999999 0 0.0007618000000000001 0 0.0007619 3.3 0.0007618200000000001 3.3 0.00076192 0 0.0007618400000000001 0 0.00076194 3.3 0.0007618600000000001 3.3 0.00076196 0 0.00076188 0 0.00076198 3.3 0.0007619 3.3 0.000762 0 0.00076192 0 0.00076202 3.3 0.00076194 3.3 0.00076204 0 0.00076196 0 0.00076206 3.3 0.00076198 3.3 0.0007620799999999999 0 0.0007620000000000001 0 0.0007621 3.3 0.0007620200000000001 3.3 0.00076212 0 0.0007620400000000001 0 0.00076214 3.3 0.0007620600000000001 3.3 0.00076216 0 0.00076208 0 0.00076218 3.3 0.0007621 3.3 0.0007622 0 0.00076212 0 0.00076222 3.3 0.00076214 3.3 0.00076224 0 0.00076216 0 0.00076226 3.3 0.00076218 3.3 0.0007622799999999999 0 0.0007622 0 0.0007622999999999999 3.3 0.0007622200000000001 3.3 0.00076232 0 0.0007622400000000001 0 0.00076234 3.3 0.0007622600000000001 3.3 0.00076236 0 0.00076228 0 0.00076238 3.3 0.0007623 3.3 0.0007624 0 0.00076232 0 0.00076242 3.3 0.00076234 3.3 0.00076244 0 0.00076236 0 0.00076246 3.3 0.00076238 3.3 0.00076248 0 0.0007624 0 0.0007624999999999999 3.3 0.0007624200000000001 3.3 0.00076252 0 0.0007624400000000001 0 0.00076254 3.3 0.0007624600000000001 3.3 0.00076256 0 0.0007624800000000001 0 0.00076258 3.3 0.0007625 3.3 0.0007626 0 0.00076252 0 0.00076262 3.3 0.00076254 3.3 0.00076264 0 0.00076256 0 0.00076266 3.3 0.00076258 3.3 0.00076268 0 0.0007626 0 0.0007626999999999999 3.3 0.00076262 3.3 0.0007627199999999999 0 0.0007626400000000001 0 0.00076274 3.3 0.0007626600000000001 3.3 0.00076276 0 0.0007626800000000001 0 0.00076278 3.3 0.0007627 3.3 0.0007628 0 0.00076272 0 0.00076282 3.3 0.00076274 3.3 0.00076284 0 0.00076276 0 0.00076286 3.3 0.00076278 3.3 0.00076288 0 0.0007628 0 0.0007629 3.3 0.00076282 3.3 0.0007629199999999999 0 0.0007628400000000001 0 0.00076294 3.3 0.0007628600000000001 3.3 0.00076296 0 0.0007628800000000001 0 0.00076298 3.3 0.0007629000000000001 3.3 0.000763 0 0.00076292 0 0.00076302 3.3 0.00076294 3.3 0.00076304 0 0.00076296 0 0.00076306 3.3 0.00076298 3.3 0.00076308 0 0.000763 0 0.0007631 3.3 0.00076302 3.3 0.0007631199999999999 0 0.00076304 0 0.0007631399999999999 3.3 0.0007630600000000001 3.3 0.00076316 0 0.0007630800000000001 0 0.00076318 3.3 0.0007631000000000001 3.3 0.0007632 0 0.00076312 0 0.00076322 3.3 0.00076314 3.3 0.00076324 0 0.00076316 0 0.00076326 3.3 0.00076318 3.3 0.00076328 0 0.0007632 0 0.0007633 3.3 0.00076322 3.3 0.00076332 0 0.00076324 0 0.0007633399999999999 3.3 0.0007632600000000001 3.3 0.00076336 0 0.0007632800000000001 0 0.00076338 3.3 0.0007633000000000001 3.3 0.0007634 0 0.0007633200000000001 0 0.00076342 3.3 0.00076334 3.3 0.00076344 0 0.00076336 0 0.00076346 3.3 0.00076338 3.3 0.00076348 0 0.0007634 0 0.0007635 3.3 0.00076342 3.3 0.00076352 0 0.00076344 0 0.0007635399999999999 3.3 0.00076346 3.3 0.0007635599999999999 0 0.0007634800000000001 0 0.00076358 3.3 0.0007635000000000001 3.3 0.0007636 0 0.0007635200000000001 0 0.00076362 3.3 0.00076354 3.3 0.00076364 0 0.00076356 0 0.00076366 3.3 0.00076358 3.3 0.00076368 0 0.0007636 0 0.0007637 3.3 0.00076362 3.3 0.00076372 0 0.00076364 0 0.00076374 3.3 0.00076366 3.3 0.0007637599999999999 0 0.0007636800000000001 0 0.00076378 3.3 0.0007637000000000001 3.3 0.0007638 0 0.0007637200000000001 0 0.00076382 3.3 0.0007637400000000001 3.3 0.00076384 0 0.00076376 0 0.00076386 3.3 0.00076378 3.3 0.00076388 0 0.0007638 0 0.0007639 3.3 0.00076382 3.3 0.00076392 0 0.00076384 0 0.00076394 3.3 0.00076386 3.3 0.0007639599999999999 0 0.00076388 0 0.0007639799999999999 3.3 0.0007639000000000001 3.3 0.000764 0 0.0007639200000000001 0 0.00076402 3.3 0.0007639400000000001 3.3 0.00076404 0 0.00076396 0 0.00076406 3.3 0.00076398 3.3 0.00076408 0 0.000764 0 0.0007641 3.3 0.00076402 3.3 0.00076412 0 0.00076404 0 0.00076414 3.3 0.00076406 3.3 0.00076416 0 0.00076408 0 0.0007641799999999999 3.3 0.0007641000000000001 3.3 0.0007642 0 0.0007641200000000001 0 0.00076422 3.3 0.0007641400000000001 3.3 0.00076424 0 0.0007641600000000001 0 0.00076426 3.3 0.00076418 3.3 0.00076428 0 0.0007642 0 0.0007643 3.3 0.00076422 3.3 0.00076432 0 0.00076424 0 0.00076434 3.3 0.00076426 3.3 0.00076436 0 0.00076428 0 0.0007643799999999999 3.3 0.0007643 3.3 0.0007643999999999999 0 0.0007643200000000001 0 0.00076442 3.3 0.0007643400000000001 3.3 0.00076444 0 0.0007643600000000001 0 0.00076446 3.3 0.00076438 3.3 0.00076448 0 0.0007644 0 0.0007645 3.3 0.00076442 3.3 0.00076452 0 0.00076444 0 0.00076454 3.3 0.00076446 3.3 0.00076456 0 0.00076448 0 0.00076458 3.3 0.0007645 3.3 0.0007645999999999999 0 0.0007645200000000001 0 0.00076462 3.3 0.0007645400000000001 3.3 0.00076464 0 0.0007645600000000001 0 0.00076466 3.3 0.0007645800000000001 3.3 0.00076468 0 0.0007646 0 0.0007647 3.3 0.00076462 3.3 0.00076472 0 0.00076464 0 0.00076474 3.3 0.00076466 3.3 0.00076476 0 0.00076468 0 0.00076478 3.3 0.0007647 3.3 0.0007647999999999999 0 0.00076472 0 0.0007648199999999999 3.3 0.0007647400000000001 3.3 0.00076484 0 0.0007647600000000001 0 0.00076486 3.3 0.0007647800000000001 3.3 0.00076488 0 0.0007648 0 0.0007649 3.3 0.00076482 3.3 0.00076492 0 0.00076484 0 0.00076494 3.3 0.00076486 3.3 0.00076496 0 0.00076488 0 0.00076498 3.3 0.0007649 3.3 0.000765 0 0.00076492 0 0.0007650199999999999 3.3 0.0007649400000000001 3.3 0.00076504 0 0.0007649600000000001 0 0.00076506 3.3 0.0007649800000000001 3.3 0.00076508 0 0.0007650000000000001 0 0.0007651 3.3 0.00076502 3.3 0.00076512 0 0.00076504 0 0.00076514 3.3 0.00076506 3.3 0.00076516 0 0.00076508 0 0.00076518 3.3 0.0007651 3.3 0.0007652 0 0.00076512 0 0.0007652199999999999 3.3 0.00076514 3.3 0.0007652399999999999 0 0.0007651600000000001 0 0.00076526 3.3 0.0007651800000000001 3.3 0.00076528 0 0.0007652000000000001 0 0.0007653 3.3 0.00076522 3.3 0.00076532 0 0.00076524 0 0.00076534 3.3 0.00076526 3.3 0.00076536 0 0.00076528 0 0.00076538 3.3 0.0007653 3.3 0.0007654 0 0.00076532 0 0.00076542 3.3 0.00076534 3.3 0.0007654399999999999 0 0.0007653600000000001 0 0.00076546 3.3 0.0007653800000000001 3.3 0.00076548 0 0.0007654000000000001 0 0.0007655 3.3 0.0007654200000000001 3.3 0.00076552 0 0.00076544 0 0.00076554 3.3 0.00076546 3.3 0.00076556 0 0.00076548 0 0.00076558 3.3 0.0007655 3.3 0.0007656 0 0.00076552 0 0.00076562 3.3 0.00076554 3.3 0.0007656399999999999 0 0.0007655600000000001 0 0.00076566 3.3 0.0007655800000000001 3.3 0.00076568 0 0.0007656000000000001 0 0.0007657 3.3 0.0007656200000000001 3.3 0.00076572 0 0.00076564 0 0.00076574 3.3 0.00076566 3.3 0.00076576 0 0.00076568 0 0.00076578 3.3 0.0007657 3.3 0.0007658 0 0.00076572 0 0.00076582 3.3 0.00076574 3.3 0.0007658399999999999 0 0.00076576 0 0.0007658599999999999 3.3 0.0007657800000000001 3.3 0.00076588 0 0.0007658000000000001 0 0.0007659 3.3 0.0007658200000000001 3.3 0.00076592 0 0.00076584 0 0.00076594 3.3 0.00076586 3.3 0.00076596 0 0.00076588 0 0.00076598 3.3 0.0007659 3.3 0.000766 0 0.00076592 0 0.00076602 3.3 0.00076594 3.3 0.00076604 0 0.00076596 0 0.0007660599999999999 3.3 0.0007659800000000001 3.3 0.00076608 0 0.0007660000000000001 0 0.0007661 3.3 0.0007660200000000001 3.3 0.00076612 0 0.0007660400000000001 0 0.00076614 3.3 0.00076606 3.3 0.00076616 0 0.00076608 0 0.00076618 3.3 0.0007661 3.3 0.0007662 0 0.00076612 0 0.00076622 3.3 0.00076614 3.3 0.00076624 0 0.00076616 0 0.0007662599999999999 3.3 0.00076618 3.3 0.0007662799999999999 0 0.0007662000000000001 0 0.0007663 3.3 0.0007662200000000001 3.3 0.00076632 0 0.0007662400000000001 0 0.00076634 3.3 0.00076626 3.3 0.00076636 0 0.00076628 0 0.00076638 3.3 0.0007663 3.3 0.0007664 0 0.00076632 0 0.00076642 3.3 0.00076634 3.3 0.00076644 0 0.00076636 0 0.00076646 3.3 0.00076638 3.3 0.0007664799999999999 0 0.0007664000000000001 0 0.0007665 3.3 0.0007664200000000001 3.3 0.00076652 0 0.0007664400000000001 0 0.00076654 3.3 0.0007664600000000001 3.3 0.00076656 0 0.00076648 0 0.00076658 3.3 0.0007665 3.3 0.0007666 0 0.00076652 0 0.00076662 3.3 0.00076654 3.3 0.00076664 0 0.00076656 0 0.00076666 3.3 0.00076658 3.3 0.0007666799999999999 0 0.0007666 0 0.0007666999999999999 3.3 0.0007666200000000001 3.3 0.00076672 0 0.0007666400000000001 0 0.00076674 3.3 0.0007666600000000001 3.3 0.00076676 0 0.00076668 0 0.00076678 3.3 0.0007667 3.3 0.0007668 0 0.00076672 0 0.00076682 3.3 0.00076674 3.3 0.00076684 0 0.00076676 0 0.00076686 3.3 0.00076678 3.3 0.00076688 0 0.0007668 0 0.0007668999999999999 3.3 0.0007668200000000001 3.3 0.00076692 0 0.0007668400000000001 0 0.00076694 3.3 0.0007668600000000001 3.3 0.00076696 0 0.0007668800000000001 0 0.00076698 3.3 0.0007669 3.3 0.000767 0 0.00076692 0 0.00076702 3.3 0.00076694 3.3 0.00076704 0 0.00076696 0 0.00076706 3.3 0.00076698 3.3 0.00076708 0 0.000767 0 0.0007670999999999999 3.3 0.00076702 3.3 0.0007671199999999999 0 0.0007670400000000001 0 0.00076714 3.3 0.0007670600000000001 3.3 0.00076716 0 0.0007670800000000001 0 0.00076718 3.3 0.0007671 3.3 0.0007672 0 0.00076712 0 0.00076722 3.3 0.00076714 3.3 0.00076724 0 0.00076716 0 0.00076726 3.3 0.00076718 3.3 0.00076728 0 0.0007672 0 0.0007673 3.3 0.00076722 3.3 0.0007673199999999999 0 0.0007672400000000001 0 0.00076734 3.3 0.0007672600000000001 3.3 0.00076736 0 0.0007672800000000001 0 0.00076738 3.3 0.0007673000000000001 3.3 0.0007674 0 0.00076732 0 0.00076742 3.3 0.00076734 3.3 0.00076744 0 0.00076736 0 0.00076746 3.3 0.00076738 3.3 0.00076748 0 0.0007674 0 0.0007675 3.3 0.00076742 3.3 0.0007675199999999999 0 0.00076744 0 0.0007675399999999999 3.3 0.0007674600000000001 3.3 0.00076756 0 0.0007674800000000001 0 0.00076758 3.3 0.0007675000000000001 3.3 0.0007676 0 0.00076752 0 0.00076762 3.3 0.00076754 3.3 0.00076764 0 0.00076756 0 0.00076766 3.3 0.00076758 3.3 0.00076768 0 0.0007676 0 0.0007677 3.3 0.00076762 3.3 0.00076772 0 0.00076764 0 0.0007677399999999999 3.3 0.0007676600000000001 3.3 0.00076776 0 0.0007676800000000001 0 0.00076778 3.3 0.0007677000000000001 3.3 0.0007678 0 0.0007677200000000001 0 0.00076782 3.3 0.00076774 3.3 0.00076784 0 0.00076776 0 0.00076786 3.3 0.00076778 3.3 0.00076788 0 0.0007678 0 0.0007679 3.3 0.00076782 3.3 0.00076792 0 0.00076784 0 0.0007679399999999999 3.3 0.00076786 3.3 0.0007679599999999999 0 0.0007678800000000001 0 0.00076798 3.3 0.0007679000000000001 3.3 0.000768 0 0.0007679200000000001 0 0.00076802 3.3 0.00076794 3.3 0.00076804 0 0.00076796 0 0.00076806 3.3 0.00076798 3.3 0.00076808 0 0.000768 0 0.0007681 3.3 0.00076802 3.3 0.00076812 0 0.00076804 0 0.00076814 3.3 0.00076806 3.3 0.0007681599999999999 0 0.0007680800000000001 0 0.00076818 3.3 0.0007681000000000001 3.3 0.0007682 0 0.0007681200000000001 0 0.00076822 3.3 0.0007681400000000001 3.3 0.00076824 0 0.00076816 0 0.00076826 3.3 0.00076818 3.3 0.00076828 0 0.0007682 0 0.0007683 3.3 0.00076822 3.3 0.00076832 0 0.00076824 0 0.00076834 3.3 0.00076826 3.3 0.0007683599999999999 0 0.00076828 0 0.0007683799999999999 3.3 0.0007683000000000001 3.3 0.0007684 0 0.0007683200000000001 0 0.00076842 3.3 0.0007683400000000001 3.3 0.00076844 0 0.00076836 0 0.00076846 3.3 0.00076838 3.3 0.00076848 0 0.0007684 0 0.0007685 3.3 0.00076842 3.3 0.00076852 0 0.00076844 0 0.00076854 3.3 0.00076846 3.3 0.00076856 0 0.00076848 0 0.0007685799999999999 3.3 0.0007685000000000001 3.3 0.0007686 0 0.0007685200000000001 0 0.00076862 3.3 0.0007685400000000001 3.3 0.00076864 0 0.0007685600000000001 0 0.00076866 3.3 0.00076858 3.3 0.00076868 0 0.0007686 0 0.0007687 3.3 0.00076862 3.3 0.00076872 0 0.00076864 0 0.00076874 3.3 0.00076866 3.3 0.00076876 0 0.00076868 0 0.0007687799999999999 3.3 0.0007687 3.3 0.0007687999999999999 0 0.0007687200000000001 0 0.00076882 3.3 0.0007687400000000001 3.3 0.00076884 0 0.0007687600000000001 0 0.00076886 3.3 0.00076878 3.3 0.00076888 0 0.0007688 0 0.0007689 3.3 0.00076882 3.3 0.00076892 0 0.00076884 0 0.00076894 3.3 0.00076886 3.3 0.00076896 0 0.00076888 0 0.0007689799999999999 3.3 0.0007689 3.3 0.0007689999999999999 0 0.0007689200000000001 0 0.00076902 3.3 0.0007689400000000001 3.3 0.00076904 0 0.0007689600000000001 0 0.00076906 3.3 0.00076898 3.3 0.00076908 0 0.000769 0 0.0007691 3.3 0.00076902 3.3 0.00076912 0 0.00076904 0 0.00076914 3.3 0.00076906 3.3 0.00076916 0 0.00076908 0 0.00076918 3.3 0.0007691 3.3 0.0007691999999999999 0 0.0007691200000000001 0 0.00076922 3.3 0.0007691400000000001 3.3 0.00076924 0 0.0007691600000000001 0 0.00076926 3.3 0.0007691800000000001 3.3 0.00076928 0 0.0007692 0 0.0007693 3.3 0.00076922 3.3 0.00076932 0 0.00076924 0 0.00076934 3.3 0.00076926 3.3 0.00076936 0 0.00076928 0 0.00076938 3.3 0.0007693 3.3 0.0007693999999999999 0 0.00076932 0 0.0007694199999999999 3.3 0.0007693400000000001 3.3 0.00076944 0 0.0007693600000000001 0 0.00076946 3.3 0.0007693800000000001 3.3 0.00076948 0 0.0007694 0 0.0007695 3.3 0.00076942 3.3 0.00076952 0 0.00076944 0 0.00076954 3.3 0.00076946 3.3 0.00076956 0 0.00076948 0 0.00076958 3.3 0.0007695 3.3 0.0007696 0 0.00076952 0 0.0007696199999999999 3.3 0.0007695400000000001 3.3 0.00076964 0 0.0007695600000000001 0 0.00076966 3.3 0.0007695800000000001 3.3 0.00076968 0 0.0007696000000000001 0 0.0007697 3.3 0.00076962 3.3 0.00076972 0 0.00076964 0 0.00076974 3.3 0.00076966 3.3 0.00076976 0 0.00076968 0 0.00076978 3.3 0.0007697 3.3 0.0007698 0 0.00076972 0 0.0007698199999999999 3.3 0.00076974 3.3 0.0007698399999999999 0 0.0007697600000000001 0 0.00076986 3.3 0.0007697800000000001 3.3 0.00076988 0 0.0007698000000000001 0 0.0007699 3.3 0.00076982 3.3 0.00076992 0 0.00076984 0 0.00076994 3.3 0.00076986 3.3 0.00076996 0 0.00076988 0 0.00076998 3.3 0.0007699 3.3 0.00077 0 0.00076992 0 0.00077002 3.3 0.00076994 3.3 0.0007700399999999999 0 0.0007699600000000001 0 0.00077006 3.3 0.0007699800000000001 3.3 0.00077008 0 0.0007700000000000001 0 0.0007701 3.3 0.0007700200000000001 3.3 0.00077012 0 0.00077004 0 0.00077014 3.3 0.00077006 3.3 0.00077016 0 0.00077008 0 0.00077018 3.3 0.0007701 3.3 0.0007702 0 0.00077012 0 0.00077022 3.3 0.00077014 3.3 0.0007702399999999999 0 0.00077016 0 0.0007702599999999999 3.3 0.0007701800000000001 3.3 0.00077028 0 0.0007702000000000001 0 0.0007703 3.3 0.0007702200000000001 3.3 0.00077032 0 0.00077024 0 0.00077034 3.3 0.00077026 3.3 0.00077036 0 0.00077028 0 0.00077038 3.3 0.0007703 3.3 0.0007704 0 0.00077032 0 0.00077042 3.3 0.00077034 3.3 0.00077044 0 0.00077036 0 0.0007704599999999999 3.3 0.0007703800000000001 3.3 0.00077048 0 0.0007704000000000001 0 0.0007705 3.3 0.0007704200000000001 3.3 0.00077052 0 0.0007704400000000001 0 0.00077054 3.3 0.00077046 3.3 0.00077056 0 0.00077048 0 0.00077058 3.3 0.0007705 3.3 0.0007706 0 0.00077052 0 0.00077062 3.3 0.00077054 3.3 0.00077064 0 0.00077056 0 0.0007706599999999999 3.3 0.00077058 3.3 0.0007706799999999999 0 0.0007706000000000001 0 0.0007707 3.3 0.0007706200000000001 3.3 0.00077072 0 0.0007706400000000001 0 0.00077074 3.3 0.00077066 3.3 0.00077076 0 0.00077068 0 0.00077078 3.3 0.0007707 3.3 0.0007708 0 0.00077072 0 0.00077082 3.3 0.00077074 3.3 0.00077084 0 0.00077076 0 0.00077086 3.3 0.00077078 3.3 0.0007708799999999999 0 0.0007708000000000001 0 0.0007709 3.3 0.0007708200000000001 3.3 0.00077092 0 0.0007708400000000001 0 0.00077094 3.3 0.0007708600000000001 3.3 0.00077096 0 0.00077088 0 0.00077098 3.3 0.0007709 3.3 0.000771 0 0.00077092 0 0.00077102 3.3 0.00077094 3.3 0.00077104 0 0.00077096 0 0.00077106 3.3 0.00077098 3.3 0.0007710799999999999 0 0.000771 0 0.0007710999999999999 3.3 0.0007710200000000001 3.3 0.00077112 0 0.0007710400000000001 0 0.00077114 3.3 0.0007710600000000001 3.3 0.00077116 0 0.00077108 0 0.00077118 3.3 0.0007711 3.3 0.0007712 0 0.00077112 0 0.00077122 3.3 0.00077114 3.3 0.00077124 0 0.00077116 0 0.00077126 3.3 0.00077118 3.3 0.00077128 0 0.0007712 0 0.0007712999999999999 3.3 0.0007712200000000001 3.3 0.00077132 0 0.0007712400000000001 0 0.00077134 3.3 0.0007712600000000001 3.3 0.00077136 0 0.0007712800000000001 0 0.00077138 3.3 0.0007713 3.3 0.0007714 0 0.00077132 0 0.00077142 3.3 0.00077134 3.3 0.00077144 0 0.00077136 0 0.00077146 3.3 0.00077138 3.3 0.00077148 0 0.0007714 0 0.0007714999999999999 3.3 0.00077142 3.3 0.0007715199999999999 0 0.0007714400000000001 0 0.00077154 3.3 0.0007714600000000001 3.3 0.00077156 0 0.0007714800000000001 0 0.00077158 3.3 0.0007715 3.3 0.0007716 0 0.00077152 0 0.00077162 3.3 0.00077154 3.3 0.00077164 0 0.00077156 0 0.00077166 3.3 0.00077158 3.3 0.00077168 0 0.0007716 0 0.0007717 3.3 0.00077162 3.3 0.0007717199999999999 0 0.0007716400000000001 0 0.00077174 3.3 0.0007716600000000001 3.3 0.00077176 0 0.0007716800000000001 0 0.00077178 3.3 0.0007717000000000001 3.3 0.0007718 0 0.00077172 0 0.00077182 3.3 0.00077174 3.3 0.00077184 0 0.00077176 0 0.00077186 3.3 0.00077178 3.3 0.00077188 0 0.0007718 0 0.0007719 3.3 0.00077182 3.3 0.0007719199999999999 0 0.00077184 0 0.0007719399999999999 3.3 0.0007718600000000001 3.3 0.00077196 0 0.0007718800000000001 0 0.00077198 3.3 0.0007719000000000001 3.3 0.000772 0 0.00077192 0 0.00077202 3.3 0.00077194 3.3 0.00077204 0 0.00077196 0 0.00077206 3.3 0.00077198 3.3 0.00077208 0 0.000772 0 0.0007721 3.3 0.00077202 3.3 0.00077212 0 0.00077204 0 0.0007721399999999999 3.3 0.0007720600000000001 3.3 0.00077216 0 0.0007720800000000001 0 0.00077218 3.3 0.0007721000000000001 3.3 0.0007722 0 0.0007721200000000001 0 0.00077222 3.3 0.00077214 3.3 0.00077224 0 0.00077216 0 0.00077226 3.3 0.00077218 3.3 0.00077228 0 0.0007722 0 0.0007723 3.3 0.00077222 3.3 0.00077232 0 0.00077224 0 0.0007723399999999999 3.3 0.00077226 3.3 0.0007723599999999999 0 0.0007722800000000001 0 0.00077238 3.3 0.0007723000000000001 3.3 0.0007724 0 0.0007723200000000001 0 0.00077242 3.3 0.00077234 3.3 0.00077244 0 0.00077236 0 0.00077246 3.3 0.00077238 3.3 0.00077248 0 0.0007724 0 0.0007725 3.3 0.00077242 3.3 0.00077252 0 0.00077244 0 0.0007725399999999999 3.3 0.00077246 3.3 0.0007725599999999999 0 0.0007724800000000001 0 0.00077258 3.3 0.0007725000000000001 3.3 0.0007726 0 0.0007725200000000001 0 0.00077262 3.3 0.00077254 3.3 0.00077264 0 0.00077256 0 0.00077266 3.3 0.00077258 3.3 0.00077268 0 0.0007726 0 0.0007727 3.3 0.00077262 3.3 0.00077272 0 0.00077264 0 0.00077274 3.3 0.00077266 3.3 0.0007727599999999999 0 0.0007726800000000001 0 0.00077278 3.3 0.0007727000000000001 3.3 0.0007728 0 0.0007727200000000001 0 0.00077282 3.3 0.0007727400000000001 3.3 0.00077284 0 0.00077276 0 0.00077286 3.3 0.00077278 3.3 0.00077288 0 0.0007728 0 0.0007729 3.3 0.00077282 3.3 0.00077292 0 0.00077284 0 0.00077294 3.3 0.00077286 3.3 0.0007729599999999999 0 0.00077288 0 0.0007729799999999999 3.3 0.0007729000000000001 3.3 0.000773 0 0.0007729200000000001 0 0.00077302 3.3 0.0007729400000000001 3.3 0.00077304 0 0.00077296 0 0.00077306 3.3 0.00077298 3.3 0.00077308 0 0.000773 0 0.0007731 3.3 0.00077302 3.3 0.00077312 0 0.00077304 0 0.00077314 3.3 0.00077306 3.3 0.00077316 0 0.00077308 0 0.0007731799999999999 3.3 0.0007731000000000001 3.3 0.0007732 0 0.0007731200000000001 0 0.00077322 3.3 0.0007731400000000001 3.3 0.00077324 0 0.0007731600000000001 0 0.00077326 3.3 0.00077318 3.3 0.00077328 0 0.0007732 0 0.0007733 3.3 0.00077322 3.3 0.00077332 0 0.00077324 0 0.00077334 3.3 0.00077326 3.3 0.00077336 0 0.00077328 0 0.0007733799999999999 3.3 0.0007733 3.3 0.0007733999999999999 0 0.0007733200000000001 0 0.00077342 3.3 0.0007733400000000001 3.3 0.00077344 0 0.0007733600000000001 0 0.00077346 3.3 0.00077338 3.3 0.00077348 0 0.0007734 0 0.0007735 3.3 0.00077342 3.3 0.00077352 0 0.00077344 0 0.00077354 3.3 0.00077346 3.3 0.00077356 0 0.00077348 0 0.00077358 3.3 0.0007735 3.3 0.0007735999999999999 0 0.0007735200000000001 0 0.00077362 3.3 0.0007735400000000001 3.3 0.00077364 0 0.0007735600000000001 0 0.00077366 3.3 0.0007735800000000001 3.3 0.00077368 0 0.0007736 0 0.0007737 3.3 0.00077362 3.3 0.00077372 0 0.00077364 0 0.00077374 3.3 0.00077366 3.3 0.00077376 0 0.00077368 0 0.00077378 3.3 0.0007737 3.3 0.0007737999999999999 0 0.00077372 0 0.0007738199999999999 3.3 0.0007737400000000001 3.3 0.00077384 0 0.0007737600000000001 0 0.00077386 3.3 0.0007737800000000001 3.3 0.00077388 0 0.0007738 0 0.0007739 3.3 0.00077382 3.3 0.00077392 0 0.00077384 0 0.00077394 3.3 0.00077386 3.3 0.00077396 0 0.00077388 0 0.00077398 3.3 0.0007739 3.3 0.000774 0 0.00077392 0 0.0007740199999999999 3.3 0.0007739400000000001 3.3 0.00077404 0 0.0007739600000000001 0 0.00077406 3.3 0.0007739800000000001 3.3 0.00077408 0 0.0007740000000000001 0 0.0007741 3.3 0.00077402 3.3 0.00077412 0 0.00077404 0 0.00077414 3.3 0.00077406 3.3 0.00077416 0 0.00077408 0 0.00077418 3.3 0.0007741 3.3 0.0007742 0 0.00077412 0 0.0007742199999999999 3.3 0.00077414 3.3 0.0007742399999999999 0 0.0007741600000000001 0 0.00077426 3.3 0.0007741800000000001 3.3 0.00077428 0 0.0007742000000000001 0 0.0007743 3.3 0.00077422 3.3 0.00077432 0 0.00077424 0 0.00077434 3.3 0.00077426 3.3 0.00077436 0 0.00077428 0 0.00077438 3.3 0.0007743 3.3 0.0007744 0 0.00077432 0 0.00077442 3.3 0.00077434 3.3 0.0007744399999999999 0 0.0007743600000000001 0 0.00077446 3.3 0.0007743800000000001 3.3 0.00077448 0 0.0007744000000000001 0 0.0007745 3.3 0.0007744200000000001 3.3 0.00077452 0 0.00077444 0 0.00077454 3.3 0.00077446 3.3 0.00077456 0 0.00077448 0 0.00077458 3.3 0.0007745 3.3 0.0007746 0 0.00077452 0 0.00077462 3.3 0.00077454 3.3 0.0007746399999999999 0 0.00077456 0 0.0007746599999999999 3.3 0.0007745800000000001 3.3 0.00077468 0 0.0007746000000000001 0 0.0007747 3.3 0.0007746200000000001 3.3 0.00077472 0 0.00077464 0 0.00077474 3.3 0.00077466 3.3 0.00077476 0 0.00077468 0 0.00077478 3.3 0.0007747 3.3 0.0007748 0 0.00077472 0 0.00077482 3.3 0.00077474 3.3 0.00077484 0 0.00077476 0 0.0007748599999999999 3.3 0.0007747800000000001 3.3 0.00077488 0 0.0007748000000000001 0 0.0007749 3.3 0.0007748200000000001 3.3 0.00077492 0 0.0007748400000000001 0 0.00077494 3.3 0.00077486 3.3 0.00077496 0 0.00077488 0 0.00077498 3.3 0.0007749 3.3 0.000775 0 0.00077492 0 0.00077502 3.3 0.00077494 3.3 0.00077504 0 0.00077496 0 0.0007750599999999999 3.3 0.00077498 3.3 0.0007750799999999999 0 0.0007750000000000001 0 0.0007751 3.3 0.0007750200000000001 3.3 0.00077512 0 0.0007750400000000001 0 0.00077514 3.3 0.00077506 3.3 0.00077516 0 0.00077508 0 0.00077518 3.3 0.0007751 3.3 0.0007752 0 0.00077512 0 0.00077522 3.3 0.00077514 3.3 0.00077524 0 0.00077516 0 0.00077526 3.3 0.00077518 3.3 0.0007752799999999999 0 0.0007752000000000001 0 0.0007753 3.3 0.0007752200000000001 3.3 0.00077532 0 0.0007752400000000001 0 0.00077534 3.3 0.0007752600000000001 3.3 0.00077536 0 0.00077528 0 0.00077538 3.3 0.0007753 3.3 0.0007754 0 0.00077532 0 0.00077542 3.3 0.00077534 3.3 0.00077544 0 0.00077536 0 0.00077546 3.3 0.00077538 3.3 0.0007754799999999999 0 0.0007754 0 0.0007754999999999999 3.3 0.0007754200000000001 3.3 0.00077552 0 0.0007754400000000001 0 0.00077554 3.3 0.0007754600000000001 3.3 0.00077556 0 0.00077548 0 0.00077558 3.3 0.0007755 3.3 0.0007756 0 0.00077552 0 0.00077562 3.3 0.00077554 3.3 0.00077564 0 0.00077556 0 0.00077566 3.3 0.00077558 3.3 0.00077568 0 0.0007756 0 0.0007756999999999999 3.3 0.0007756200000000001 3.3 0.00077572 0 0.0007756400000000001 0 0.00077574 3.3 0.0007756600000000001 3.3 0.00077576 0 0.0007756800000000001 0 0.00077578 3.3 0.0007757 3.3 0.0007758 0 0.00077572 0 0.00077582 3.3 0.00077574 3.3 0.00077584 0 0.00077576 0 0.00077586 3.3 0.00077578 3.3 0.00077588 0 0.0007758 0 0.0007758999999999999 3.3 0.0007758200000000001 3.3 0.00077592 0 0.0007758400000000001 0 0.00077594 3.3 0.0007758600000000001 3.3 0.00077596 0 0.0007758800000000001 0 0.00077598 3.3 0.0007759 3.3 0.000776 0 0.00077592 0 0.00077602 3.3 0.00077594 3.3 0.00077604 0 0.00077596 0 0.00077606 3.3 0.00077598 3.3 0.00077608 0 0.000776 0 0.0007760999999999999 3.3 0.00077602 3.3 0.0007761199999999999 0 0.0007760400000000001 0 0.00077614 3.3 0.0007760600000000001 3.3 0.00077616 0 0.0007760800000000001 0 0.00077618 3.3 0.0007761 3.3 0.0007762 0 0.00077612 0 0.00077622 3.3 0.00077614 3.3 0.00077624 0 0.00077616 0 0.00077626 3.3 0.00077618 3.3 0.00077628 0 0.0007762 0 0.0007763 3.3 0.00077622 3.3 0.0007763199999999999 0 0.0007762400000000001 0 0.00077634 3.3 0.0007762600000000001 3.3 0.00077636 0 0.0007762800000000001 0 0.00077638 3.3 0.0007763000000000001 3.3 0.0007764 0 0.00077632 0 0.00077642 3.3 0.00077634 3.3 0.00077644 0 0.00077636 0 0.00077646 3.3 0.00077638 3.3 0.00077648 0 0.0007764 0 0.0007765 3.3 0.00077642 3.3 0.0007765199999999999 0 0.00077644 0 0.0007765399999999999 3.3 0.0007764600000000001 3.3 0.00077656 0 0.0007764800000000001 0 0.00077658 3.3 0.0007765000000000001 3.3 0.0007766 0 0.00077652 0 0.00077662 3.3 0.00077654 3.3 0.00077664 0 0.00077656 0 0.00077666 3.3 0.00077658 3.3 0.00077668 0 0.0007766 0 0.0007767 3.3 0.00077662 3.3 0.00077672 0 0.00077664 0 0.0007767399999999999 3.3 0.0007766600000000001 3.3 0.00077676 0 0.0007766800000000001 0 0.00077678 3.3 0.0007767000000000001 3.3 0.0007768 0 0.0007767200000000001 0 0.00077682 3.3 0.00077674 3.3 0.00077684 0 0.00077676 0 0.00077686 3.3 0.00077678 3.3 0.00077688 0 0.0007768 0 0.0007769 3.3 0.00077682 3.3 0.00077692 0 0.00077684 0 0.0007769399999999999 3.3 0.00077686 3.3 0.0007769599999999999 0 0.0007768800000000001 0 0.00077698 3.3 0.0007769000000000001 3.3 0.000777 0 0.0007769200000000001 0 0.00077702 3.3 0.00077694 3.3 0.00077704 0 0.00077696 0 0.00077706 3.3 0.00077698 3.3 0.00077708 0 0.000777 0 0.0007771 3.3 0.00077702 3.3 0.00077712 0 0.00077704 0 0.00077714 3.3 0.00077706 3.3 0.0007771599999999999 0 0.0007770800000000001 0 0.00077718 3.3 0.0007771000000000001 3.3 0.0007772 0 0.0007771200000000001 0 0.00077722 3.3 0.0007771400000000001 3.3 0.00077724 0 0.00077716 0 0.00077726 3.3 0.00077718 3.3 0.00077728 0 0.0007772 0 0.0007773 3.3 0.00077722 3.3 0.00077732 0 0.00077724 0 0.00077734 3.3 0.00077726 3.3 0.0007773599999999999 0 0.00077728 0 0.0007773799999999999 3.3 0.0007773000000000001 3.3 0.0007774 0 0.0007773200000000001 0 0.00077742 3.3 0.0007773400000000001 3.3 0.00077744 0 0.00077736 0 0.00077746 3.3 0.00077738 3.3 0.00077748 0 0.0007774 0 0.0007775 3.3 0.00077742 3.3 0.00077752 0 0.00077744 0 0.00077754 3.3 0.00077746 3.3 0.00077756 0 0.00077748 0 0.0007775799999999999 3.3 0.0007775000000000001 3.3 0.0007776 0 0.0007775200000000001 0 0.00077762 3.3 0.0007775400000000001 3.3 0.00077764 0 0.0007775600000000001 0 0.00077766 3.3 0.00077758 3.3 0.00077768 0 0.0007776 0 0.0007777 3.3 0.00077762 3.3 0.00077772 0 0.00077764 0 0.00077774 3.3 0.00077766 3.3 0.00077776 0 0.00077768 0 0.0007777799999999999 3.3 0.0007777 3.3 0.0007777999999999999 0 0.0007777200000000001 0 0.00077782 3.3 0.0007777400000000001 3.3 0.00077784 0 0.0007777600000000001 0 0.00077786 3.3 0.00077778 3.3 0.00077788 0 0.0007778 0 0.0007779 3.3 0.00077782 3.3 0.00077792 0 0.00077784 0 0.00077794 3.3 0.00077786 3.3 0.00077796 0 0.00077788 0 0.00077798 3.3 0.0007779 3.3 0.0007779999999999999 0 0.0007779200000000001 0 0.00077802 3.3 0.0007779400000000001 3.3 0.00077804 0 0.0007779600000000001 0 0.00077806 3.3 0.0007779800000000001 3.3 0.00077808 0 0.000778 0 0.0007781 3.3 0.00077802 3.3 0.00077812 0 0.00077804 0 0.00077814 3.3 0.00077806 3.3 0.00077816 0 0.00077808 0 0.00077818 3.3 0.0007781 3.3 0.0007781999999999999 0 0.00077812 0 0.0007782199999999999 3.3 0.0007781400000000001 3.3 0.00077824 0 0.0007781600000000001 0 0.00077826 3.3 0.0007781800000000001 3.3 0.00077828 0 0.0007782 0 0.0007783 3.3 0.00077822 3.3 0.00077832 0 0.00077824 0 0.00077834 3.3 0.00077826 3.3 0.00077836 0 0.00077828 0 0.00077838 3.3 0.0007783 3.3 0.0007784 0 0.00077832 0 0.0007784199999999999 3.3 0.0007783400000000001 3.3 0.00077844 0 0.0007783600000000001 0 0.00077846 3.3 0.0007783800000000001 3.3 0.00077848 0 0.0007784000000000001 0 0.0007785 3.3 0.00077842 3.3 0.00077852 0 0.00077844 0 0.00077854 3.3 0.00077846 3.3 0.00077856 0 0.00077848 0 0.00077858 3.3 0.0007785 3.3 0.0007786 0 0.00077852 0 0.0007786199999999999 3.3 0.00077854 3.3 0.0007786399999999999 0 0.0007785600000000001 0 0.00077866 3.3 0.0007785800000000001 3.3 0.00077868 0 0.0007786000000000001 0 0.0007787 3.3 0.00077862 3.3 0.00077872 0 0.00077864 0 0.00077874 3.3 0.00077866 3.3 0.00077876 0 0.00077868 0 0.00077878 3.3 0.0007787 3.3 0.0007788 0 0.00077872 0 0.00077882 3.3 0.00077874 3.3 0.0007788399999999999 0 0.0007787600000000001 0 0.00077886 3.3 0.0007787800000000001 3.3 0.00077888 0 0.0007788000000000001 0 0.0007789 3.3 0.0007788200000000001 3.3 0.00077892 0 0.00077884 0 0.00077894 3.3 0.00077886 3.3 0.00077896 0 0.00077888 0 0.00077898 3.3 0.0007789 3.3 0.000779 0 0.00077892 0 0.00077902 3.3 0.00077894 3.3 0.0007790399999999999 0 0.00077896 0 0.0007790599999999999 3.3 0.0007789800000000001 3.3 0.00077908 0 0.0007790000000000001 0 0.0007791 3.3 0.0007790200000000001 3.3 0.00077912 0 0.00077904 0 0.00077914 3.3 0.00077906 3.3 0.00077916 0 0.00077908 0 0.00077918 3.3 0.0007791 3.3 0.0007792 0 0.00077912 0 0.00077922 3.3 0.00077914 3.3 0.0007792399999999999 0 0.00077916 0 0.0007792599999999999 3.3 0.0007791800000000001 3.3 0.00077928 0 0.0007792000000000001 0 0.0007793 3.3 0.0007792200000000001 3.3 0.00077932 0 0.00077924 0 0.00077934 3.3 0.00077926 3.3 0.00077936 0 0.00077928 0 0.00077938 3.3 0.0007793 3.3 0.0007794 0 0.00077932 0 0.00077942 3.3 0.00077934 3.3 0.00077944 0 0.00077936 0 0.0007794599999999999 3.3 0.0007793800000000001 3.3 0.00077948 0 0.0007794000000000001 0 0.0007795 3.3 0.0007794200000000001 3.3 0.00077952 0 0.0007794400000000001 0 0.00077954 3.3 0.00077946 3.3 0.00077956 0 0.00077948 0 0.00077958 3.3 0.0007795 3.3 0.0007796 0 0.00077952 0 0.00077962 3.3 0.00077954 3.3 0.00077964 0 0.00077956 0 0.0007796599999999999 3.3 0.00077958 3.3 0.0007796799999999999 0 0.0007796000000000001 0 0.0007797 3.3 0.0007796200000000001 3.3 0.00077972 0 0.0007796400000000001 0 0.00077974 3.3 0.00077966 3.3 0.00077976 0 0.00077968 0 0.00077978 3.3 0.0007797 3.3 0.0007798 0 0.00077972 0 0.00077982 3.3 0.00077974 3.3 0.00077984 0 0.00077976 0 0.00077986 3.3 0.00077978 3.3 0.0007798799999999999 0 0.0007798000000000001 0 0.0007799 3.3 0.0007798200000000001 3.3 0.00077992 0 0.0007798400000000001 0 0.00077994 3.3 0.0007798600000000001 3.3 0.00077996 0 0.00077988 0 0.00077998 3.3 0.0007799 3.3 0.00078 0 0.00077992 0 0.00078002 3.3 0.00077994 3.3 0.00078004 0 0.00077996 0 0.00078006 3.3 0.00077998 3.3 0.0007800799999999999 0 0.00078 0 0.0007800999999999999 3.3 0.0007800200000000001 3.3 0.00078012 0 0.0007800400000000001 0 0.00078014 3.3 0.0007800600000000001 3.3 0.00078016 0 0.00078008 0 0.00078018 3.3 0.0007801 3.3 0.0007802 0 0.00078012 0 0.00078022 3.3 0.00078014 3.3 0.00078024 0 0.00078016 0 0.00078026 3.3 0.00078018 3.3 0.00078028 0 0.0007802 0 0.0007802999999999999 3.3 0.0007802200000000001 3.3 0.00078032 0 0.0007802400000000001 0 0.00078034 3.3 0.0007802600000000001 3.3 0.00078036 0 0.0007802800000000001 0 0.00078038 3.3 0.0007803 3.3 0.0007804 0 0.00078032 0 0.00078042 3.3 0.00078034 3.3 0.00078044 0 0.00078036 0 0.00078046 3.3 0.00078038 3.3 0.00078048 0 0.0007804 0 0.0007804999999999999 3.3 0.00078042 3.3 0.0007805199999999999 0 0.0007804400000000001 0 0.00078054 3.3 0.0007804600000000001 3.3 0.00078056 0 0.0007804800000000001 0 0.00078058 3.3 0.0007805 3.3 0.0007806 0 0.00078052 0 0.00078062 3.3 0.00078054 3.3 0.00078064 0 0.00078056 0 0.00078066 3.3 0.00078058 3.3 0.00078068 0 0.0007806 0 0.0007807 3.3 0.00078062 3.3 0.0007807199999999999 0 0.0007806400000000001 0 0.00078074 3.3 0.0007806600000000001 3.3 0.00078076 0 0.0007806800000000001 0 0.00078078 3.3 0.0007807000000000001 3.3 0.0007808 0 0.00078072 0 0.00078082 3.3 0.00078074 3.3 0.00078084 0 0.00078076 0 0.00078086 3.3 0.00078078 3.3 0.00078088 0 0.0007808 0 0.0007809 3.3 0.00078082 3.3 0.0007809199999999999 0 0.00078084 0 0.0007809399999999999 3.3 0.0007808600000000001 3.3 0.00078096 0 0.0007808800000000001 0 0.00078098 3.3 0.0007809000000000001 3.3 0.000781 0 0.00078092 0 0.00078102 3.3 0.00078094 3.3 0.00078104 0 0.00078096 0 0.00078106 3.3 0.00078098 3.3 0.00078108 0 0.000781 0 0.0007811 3.3 0.00078102 3.3 0.00078112 0 0.00078104 0 0.0007811399999999999 3.3 0.0007810600000000001 3.3 0.00078116 0 0.0007810800000000001 0 0.00078118 3.3 0.0007811000000000001 3.3 0.0007812 0 0.0007811200000000001 0 0.00078122 3.3 0.00078114 3.3 0.00078124 0 0.00078116 0 0.00078126 3.3 0.00078118 3.3 0.00078128 0 0.0007812 0 0.0007813 3.3 0.00078122 3.3 0.00078132 0 0.00078124 0 0.0007813399999999999 3.3 0.00078126 3.3 0.0007813599999999999 0 0.0007812800000000001 0 0.00078138 3.3 0.0007813000000000001 3.3 0.0007814 0 0.0007813200000000001 0 0.00078142 3.3 0.00078134 3.3 0.00078144 0 0.00078136 0 0.00078146 3.3 0.00078138 3.3 0.00078148 0 0.0007814 0 0.0007815 3.3 0.00078142 3.3 0.00078152 0 0.00078144 0 0.00078154 3.3 0.00078146 3.3 0.0007815599999999999 0 0.0007814800000000001 0 0.00078158 3.3 0.0007815000000000001 3.3 0.0007816 0 0.0007815200000000001 0 0.00078162 3.3 0.0007815400000000001 3.3 0.00078164 0 0.00078156 0 0.00078166 3.3 0.00078158 3.3 0.00078168 0 0.0007816 0 0.0007817 3.3 0.00078162 3.3 0.00078172 0 0.00078164 0 0.00078174 3.3 0.00078166 3.3 0.0007817599999999999 0 0.00078168 0 0.0007817799999999999 3.3 0.0007817000000000001 3.3 0.0007818 0 0.0007817200000000001 0 0.00078182 3.3 0.0007817400000000001 3.3 0.00078184 0 0.00078176 0 0.00078186 3.3 0.00078178 3.3 0.00078188 0 0.0007818 0 0.0007819 3.3 0.00078182 3.3 0.00078192 0 0.00078184 0 0.00078194 3.3 0.00078186 3.3 0.00078196 0 0.00078188 0 0.0007819799999999999 3.3 0.0007819000000000001 3.3 0.000782 0 0.0007819200000000001 0 0.00078202 3.3 0.0007819400000000001 3.3 0.00078204 0 0.0007819600000000001 0 0.00078206 3.3 0.00078198 3.3 0.00078208 0 0.000782 0 0.0007821 3.3 0.00078202 3.3 0.00078212 0 0.00078204 0 0.00078214 3.3 0.00078206 3.3 0.00078216 0 0.00078208 0 0.0007821799999999999 3.3 0.0007821 3.3 0.0007821999999999999 0 0.0007821200000000001 0 0.00078222 3.3 0.0007821400000000001 3.3 0.00078224 0 0.0007821600000000001 0 0.00078226 3.3 0.00078218 3.3 0.00078228 0 0.0007822 0 0.0007823 3.3 0.00078222 3.3 0.00078232 0 0.00078224 0 0.00078234 3.3 0.00078226 3.3 0.00078236 0 0.00078228 0 0.00078238 3.3 0.0007823 3.3 0.0007823999999999999 0 0.0007823200000000001 0 0.00078242 3.3 0.0007823400000000001 3.3 0.00078244 0 0.0007823600000000001 0 0.00078246 3.3 0.0007823800000000001 3.3 0.00078248 0 0.0007824 0 0.0007825 3.3 0.00078242 3.3 0.00078252 0 0.00078244 0 0.00078254 3.3 0.00078246 3.3 0.00078256 0 0.00078248 0 0.00078258 3.3 0.0007825 3.3 0.0007825999999999999 0 0.00078252 0 0.0007826199999999999 3.3 0.0007825400000000001 3.3 0.00078264 0 0.0007825600000000001 0 0.00078266 3.3 0.0007825800000000001 3.3 0.00078268 0 0.0007826 0 0.0007827 3.3 0.00078262 3.3 0.00078272 0 0.00078264 0 0.00078274 3.3 0.00078266 3.3 0.00078276 0 0.00078268 0 0.00078278 3.3 0.0007827 3.3 0.0007827999999999999 0 0.00078272 0 0.0007828199999999999 3.3 0.0007827400000000001 3.3 0.00078284 0 0.0007827600000000001 0 0.00078286 3.3 0.0007827800000000001 3.3 0.00078288 0 0.0007828 0 0.0007829 3.3 0.00078282 3.3 0.00078292 0 0.00078284 0 0.00078294 3.3 0.00078286 3.3 0.00078296 0 0.00078288 0 0.00078298 3.3 0.0007829 3.3 0.000783 0 0.00078292 0 0.0007830199999999999 3.3 0.0007829400000000001 3.3 0.00078304 0 0.0007829600000000001 0 0.00078306 3.3 0.0007829800000000001 3.3 0.00078308 0 0.0007830000000000001 0 0.0007831 3.3 0.00078302 3.3 0.00078312 0 0.00078304 0 0.00078314 3.3 0.00078306 3.3 0.00078316 0 0.00078308 0 0.00078318 3.3 0.0007831 3.3 0.0007832 0 0.00078312 0 0.0007832199999999999 3.3 0.00078314 3.3 0.0007832399999999999 0 0.0007831600000000001 0 0.00078326 3.3 0.0007831800000000001 3.3 0.00078328 0 0.0007832000000000001 0 0.0007833 3.3 0.00078322 3.3 0.00078332 0 0.00078324 0 0.00078334 3.3 0.00078326 3.3 0.00078336 0 0.00078328 0 0.00078338 3.3 0.0007833 3.3 0.0007834 0 0.00078332 0 0.00078342 3.3 0.00078334 3.3 0.0007834399999999999 0 0.0007833600000000001 0 0.00078346 3.3 0.0007833800000000001 3.3 0.00078348 0 0.0007834000000000001 0 0.0007835 3.3 0.0007834200000000001 3.3 0.00078352 0 0.00078344 0 0.00078354 3.3 0.00078346 3.3 0.00078356 0 0.00078348 0 0.00078358 3.3 0.0007835 3.3 0.0007836 0 0.00078352 0 0.00078362 3.3 0.00078354 3.3 0.0007836399999999999 0 0.00078356 0 0.0007836599999999999 3.3 0.0007835800000000001 3.3 0.00078368 0 0.0007836000000000001 0 0.0007837 3.3 0.0007836200000000001 3.3 0.00078372 0 0.00078364 0 0.00078374 3.3 0.00078366 3.3 0.00078376 0 0.00078368 0 0.00078378 3.3 0.0007837 3.3 0.0007838 0 0.00078372 0 0.00078382 3.3 0.00078374 3.3 0.00078384 0 0.00078376 0 0.0007838599999999999 3.3 0.0007837800000000001 3.3 0.00078388 0 0.0007838000000000001 0 0.0007839 3.3 0.0007838200000000001 3.3 0.00078392 0 0.0007838400000000001 0 0.00078394 3.3 0.00078386 3.3 0.00078396 0 0.00078388 0 0.00078398 3.3 0.0007839 3.3 0.000784 0 0.00078392 0 0.00078402 3.3 0.00078394 3.3 0.00078404 0 0.00078396 0 0.0007840599999999999 3.3 0.00078398 3.3 0.0007840799999999999 0 0.0007840000000000001 0 0.0007841 3.3 0.0007840200000000001 3.3 0.00078412 0 0.0007840400000000001 0 0.00078414 3.3 0.00078406 3.3 0.00078416 0 0.00078408 0 0.00078418 3.3 0.0007841 3.3 0.0007842 0 0.00078412 0 0.00078422 3.3 0.00078414 3.3 0.00078424 0 0.00078416 0 0.00078426 3.3 0.00078418 3.3 0.0007842799999999999 0 0.0007842000000000001 0 0.0007843 3.3 0.0007842200000000001 3.3 0.00078432 0 0.0007842400000000001 0 0.00078434 3.3 0.0007842600000000001 3.3 0.00078436 0 0.00078428 0 0.00078438 3.3 0.0007843 3.3 0.0007844 0 0.00078432 0 0.00078442 3.3 0.00078434 3.3 0.00078444 0 0.00078436 0 0.00078446 3.3 0.00078438 3.3 0.0007844799999999999 0 0.0007844 0 0.0007844999999999999 3.3 0.0007844200000000001 3.3 0.00078452 0 0.0007844400000000001 0 0.00078454 3.3 0.0007844600000000001 3.3 0.00078456 0 0.00078448 0 0.00078458 3.3 0.0007845 3.3 0.0007846 0 0.00078452 0 0.00078462 3.3 0.00078454 3.3 0.00078464 0 0.00078456 0 0.00078466 3.3 0.00078458 3.3 0.00078468 0 0.0007846 0 0.0007846999999999999 3.3 0.0007846200000000001 3.3 0.00078472 0 0.0007846400000000001 0 0.00078474 3.3 0.0007846600000000001 3.3 0.00078476 0 0.0007846800000000001 0 0.00078478 3.3 0.0007847 3.3 0.0007848 0 0.00078472 0 0.00078482 3.3 0.00078474 3.3 0.00078484 0 0.00078476 0 0.00078486 3.3 0.00078478 3.3 0.00078488 0 0.0007848 0 0.0007848999999999999 3.3 0.00078482 3.3 0.0007849199999999999 0 0.0007848400000000001 0 0.00078494 3.3 0.0007848600000000001 3.3 0.00078496 0 0.0007848800000000001 0 0.00078498 3.3 0.0007849 3.3 0.000785 0 0.00078492 0 0.00078502 3.3 0.00078494 3.3 0.00078504 0 0.00078496 0 0.00078506 3.3 0.00078498 3.3 0.00078508 0 0.000785 0 0.0007851 3.3 0.00078502 3.3 0.0007851199999999999 0 0.0007850400000000001 0 0.00078514 3.3 0.0007850600000000001 3.3 0.00078516 0 0.0007850800000000001 0 0.00078518 3.3 0.0007851000000000001 3.3 0.0007852 0 0.00078512 0 0.00078522 3.3 0.00078514 3.3 0.00078524 0 0.00078516 0 0.00078526 3.3 0.00078518 3.3 0.00078528 0 0.0007852 0 0.0007853 3.3 0.00078522 3.3 0.0007853199999999999 0 0.00078524 0 0.0007853399999999999 3.3 0.0007852600000000001 3.3 0.00078536 0 0.0007852800000000001 0 0.00078538 3.3 0.0007853000000000001 3.3 0.0007854 0 0.00078532 0 0.00078542 3.3 0.00078534 3.3 0.00078544 0 0.00078536 0 0.00078546 3.3 0.00078538 3.3 0.00078548 0 0.0007854 0 0.0007855 3.3 0.00078542 3.3 0.00078552 0 0.00078544 0 0.0007855399999999999 3.3 0.0007854600000000001 3.3 0.00078556 0 0.0007854800000000001 0 0.00078558 3.3 0.0007855000000000001 3.3 0.0007856 0 0.0007855200000000001 0 0.00078562 3.3 0.00078554 3.3 0.00078564 0 0.00078556 0 0.00078566 3.3 0.00078558 3.3 0.00078568 0 0.0007856 0 0.0007857 3.3 0.00078562 3.3 0.00078572 0 0.00078564 0 0.0007857399999999999 3.3 0.00078566 3.3 0.0007857599999999999 0 0.0007856800000000001 0 0.00078578 3.3 0.0007857000000000001 3.3 0.0007858 0 0.0007857200000000001 0 0.00078582 3.3 0.00078574 3.3 0.00078584 0 0.00078576 0 0.00078586 3.3 0.00078578 3.3 0.00078588 0 0.0007858 0 0.0007859 3.3 0.00078582 3.3 0.00078592 0 0.00078584 0 0.00078594 3.3 0.00078586 3.3 0.0007859599999999999 0 0.0007858800000000001 0 0.00078598 3.3 0.0007859000000000001 3.3 0.000786 0 0.0007859200000000001 0 0.00078602 3.3 0.0007859400000000001 3.3 0.00078604 0 0.00078596 0 0.00078606 3.3 0.00078598 3.3 0.00078608 0 0.000786 0 0.0007861 3.3 0.00078602 3.3 0.00078612 0 0.00078604 0 0.00078614 3.3 0.00078606 3.3 0.0007861599999999999 0 0.00078608 0 0.0007861799999999999 3.3 0.0007861000000000001 3.3 0.0007862 0 0.0007861200000000001 0 0.00078622 3.3 0.0007861400000000001 3.3 0.00078624 0 0.00078616 0 0.00078626 3.3 0.00078618 3.3 0.00078628 0 0.0007862 0 0.0007863 3.3 0.00078622 3.3 0.00078632 0 0.00078624 0 0.00078634 3.3 0.00078626 3.3 0.0007863599999999999 0 0.00078628 0 0.0007863799999999999 3.3 0.0007863000000000001 3.3 0.0007864 0 0.0007863200000000001 0 0.00078642 3.3 0.0007863400000000001 3.3 0.00078644 0 0.00078636 0 0.00078646 3.3 0.00078638 3.3 0.00078648 0 0.0007864 0 0.0007865 3.3 0.00078642 3.3 0.00078652 0 0.00078644 0 0.00078654 3.3 0.00078646 3.3 0.00078656 0 0.00078648 0 0.0007865799999999999 3.3 0.0007865000000000001 3.3 0.0007866 0 0.0007865200000000001 0 0.00078662 3.3 0.0007865400000000001 3.3 0.00078664 0 0.0007865600000000001 0 0.00078666 3.3 0.00078658 3.3 0.00078668 0 0.0007866 0 0.0007867 3.3 0.00078662 3.3 0.00078672 0 0.00078664 0 0.00078674 3.3 0.00078666 3.3 0.00078676 0 0.00078668 0 0.0007867799999999999 3.3 0.0007867 3.3 0.0007867999999999999 0 0.0007867200000000001 0 0.00078682 3.3 0.0007867400000000001 3.3 0.00078684 0 0.0007867600000000001 0 0.00078686 3.3 0.00078678 3.3 0.00078688 0 0.0007868 0 0.0007869 3.3 0.00078682 3.3 0.00078692 0 0.00078684 0 0.00078694 3.3 0.00078686 3.3 0.00078696 0 0.00078688 0 0.00078698 3.3 0.0007869 3.3 0.0007869999999999999 0 0.0007869200000000001 0 0.00078702 3.3 0.0007869400000000001 3.3 0.00078704 0 0.0007869600000000001 0 0.00078706 3.3 0.0007869800000000001 3.3 0.00078708 0 0.000787 0 0.0007871 3.3 0.00078702 3.3 0.00078712 0 0.00078704 0 0.00078714 3.3 0.00078706 3.3 0.00078716 0 0.00078708 0 0.00078718 3.3 0.0007871 3.3 0.0007871999999999999 0 0.00078712 0 0.0007872199999999999 3.3 0.0007871400000000001 3.3 0.00078724 0 0.0007871600000000001 0 0.00078726 3.3 0.0007871800000000001 3.3 0.00078728 0 0.0007872 0 0.0007873 3.3 0.00078722 3.3 0.00078732 0 0.00078724 0 0.00078734 3.3 0.00078726 3.3 0.00078736 0 0.00078728 0 0.00078738 3.3 0.0007873 3.3 0.0007874 0 0.00078732 0 0.0007874199999999999 3.3 0.0007873400000000001 3.3 0.00078744 0 0.0007873600000000001 0 0.00078746 3.3 0.0007873800000000001 3.3 0.00078748 0 0.0007874000000000001 0 0.0007875 3.3 0.00078742 3.3 0.00078752 0 0.00078744 0 0.00078754 3.3 0.00078746 3.3 0.00078756 0 0.00078748 0 0.00078758 3.3 0.0007875 3.3 0.0007876 0 0.00078752 0 0.0007876199999999999 3.3 0.00078754 3.3 0.0007876399999999999 0 0.0007875600000000001 0 0.00078766 3.3 0.0007875800000000001 3.3 0.00078768 0 0.0007876000000000001 0 0.0007877 3.3 0.00078762 3.3 0.00078772 0 0.00078764 0 0.00078774 3.3 0.00078766 3.3 0.00078776 0 0.00078768 0 0.00078778 3.3 0.0007877 3.3 0.0007878 0 0.00078772 0 0.00078782 3.3 0.00078774 3.3 0.0007878399999999999 0 0.0007877600000000001 0 0.00078786 3.3 0.0007877800000000001 3.3 0.00078788 0 0.0007878000000000001 0 0.0007879 3.3 0.0007878200000000001 3.3 0.00078792 0 0.00078784 0 0.00078794 3.3 0.00078786 3.3 0.00078796 0 0.00078788 0 0.00078798 3.3 0.0007879 3.3 0.000788 0 0.00078792 0 0.00078802 3.3 0.00078794 3.3 0.0007880399999999999 0 0.00078796 0 0.0007880599999999999 3.3 0.0007879800000000001 3.3 0.00078808 0 0.0007880000000000001 0 0.0007881 3.3 0.0007880200000000001 3.3 0.00078812 0 0.00078804 0 0.00078814 3.3 0.00078806 3.3 0.00078816 0 0.00078808 0 0.00078818 3.3 0.0007881 3.3 0.0007882 0 0.00078812 0 0.00078822 3.3 0.00078814 3.3 0.00078824 0 0.00078816 0 0.0007882599999999999 3.3 0.0007881800000000001 3.3 0.00078828 0 0.0007882000000000001 0 0.0007883 3.3 0.0007882200000000001 3.3 0.00078832 0 0.0007882400000000001 0 0.00078834 3.3 0.00078826 3.3 0.00078836 0 0.00078828 0 0.00078838 3.3 0.0007883 3.3 0.0007884 0 0.00078832 0 0.00078842 3.3 0.00078834 3.3 0.00078844 0 0.00078836 0 0.0007884599999999999 3.3 0.00078838 3.3 0.0007884799999999999 0 0.0007884000000000001 0 0.0007885 3.3 0.0007884200000000001 3.3 0.00078852 0 0.0007884400000000001 0 0.00078854 3.3 0.00078846 3.3 0.00078856 0 0.00078848 0 0.00078858 3.3 0.0007885 3.3 0.0007886 0 0.00078852 0 0.00078862 3.3 0.00078854 3.3 0.00078864 0 0.00078856 0 0.00078866 3.3 0.00078858 3.3 0.0007886799999999999 0 0.0007886000000000001 0 0.0007887 3.3 0.0007886200000000001 3.3 0.00078872 0 0.0007886400000000001 0 0.00078874 3.3 0.0007886600000000001 3.3 0.00078876 0 0.00078868 0 0.00078878 3.3 0.0007887 3.3 0.0007888 0 0.00078872 0 0.00078882 3.3 0.00078874 3.3 0.00078884 0 0.00078876 0 0.00078886 3.3 0.00078878 3.3 0.0007888799999999999 0 0.0007888 0 0.0007888999999999999 3.3 0.0007888200000000001 3.3 0.00078892 0 0.0007888400000000001 0 0.00078894 3.3 0.0007888600000000001 3.3 0.00078896 0 0.00078888 0 0.00078898 3.3 0.0007889 3.3 0.000789 0 0.00078892 0 0.00078902 3.3 0.00078894 3.3 0.00078904 0 0.00078896 0 0.00078906 3.3 0.00078898 3.3 0.00078908 0 0.000789 0 0.0007890999999999999 3.3 0.0007890200000000001 3.3 0.00078912 0 0.0007890400000000001 0 0.00078914 3.3 0.0007890600000000001 3.3 0.00078916 0 0.0007890800000000001 0 0.00078918 3.3 0.0007891 3.3 0.0007892 0 0.00078912 0 0.00078922 3.3 0.00078914 3.3 0.00078924 0 0.00078916 0 0.00078926 3.3 0.00078918 3.3 0.00078928 0 0.0007892 0 0.0007892999999999999 3.3 0.00078922 3.3 0.0007893199999999999 0 0.0007892400000000001 0 0.00078934 3.3 0.0007892600000000001 3.3 0.00078936 0 0.0007892800000000001 0 0.00078938 3.3 0.0007893 3.3 0.0007894 0 0.00078932 0 0.00078942 3.3 0.00078934 3.3 0.00078944 0 0.00078936 0 0.00078946 3.3 0.00078938 3.3 0.00078948 0 0.0007894 0 0.0007894999999999999 3.3 0.00078942 3.3 0.0007895199999999999 0 0.0007894400000000001 0 0.00078954 3.3 0.0007894600000000001 3.3 0.00078956 0 0.0007894800000000001 0 0.00078958 3.3 0.0007895 3.3 0.0007896 0 0.00078952 0 0.00078962 3.3 0.00078954 3.3 0.00078964 0 0.00078956 0 0.00078966 3.3 0.00078958 3.3 0.00078968 0 0.0007896 0 0.0007897 3.3 0.00078962 3.3 0.0007897199999999999 0 0.0007896400000000001 0 0.00078974 3.3 0.0007896600000000001 3.3 0.00078976 0 0.0007896800000000001 0 0.00078978 3.3 0.0007897000000000001 3.3 0.0007898 0 0.00078972 0 0.00078982 3.3 0.00078974 3.3 0.00078984 0 0.00078976 0 0.00078986 3.3 0.00078978 3.3 0.00078988 0 0.0007898 0 0.0007899 3.3 0.00078982 3.3 0.0007899199999999999 0 0.00078984 0 0.0007899399999999999 3.3 0.0007898600000000001 3.3 0.00078996 0 0.0007898800000000001 0 0.00078998 3.3 0.0007899000000000001 3.3 0.00079 0 0.00078992 0 0.00079002 3.3 0.00078994 3.3 0.00079004 0 0.00078996 0 0.00079006 3.3 0.00078998 3.3 0.00079008 0 0.00079 0 0.0007901 3.3 0.00079002 3.3 0.00079012 0 0.00079004 0 0.0007901399999999999 3.3 0.0007900600000000001 3.3 0.00079016 0 0.0007900800000000001 0 0.00079018 3.3 0.0007901000000000001 3.3 0.0007902 0 0.0007901200000000001 0 0.00079022 3.3 0.00079014 3.3 0.00079024 0 0.00079016 0 0.00079026 3.3 0.00079018 3.3 0.00079028 0 0.0007902 0 0.0007903 3.3 0.00079022 3.3 0.00079032 0 0.00079024 0 0.0007903399999999999 3.3 0.00079026 3.3 0.0007903599999999999 0 0.0007902800000000001 0 0.00079038 3.3 0.0007903000000000001 3.3 0.0007904 0 0.0007903200000000001 0 0.00079042 3.3 0.00079034 3.3 0.00079044 0 0.00079036 0 0.00079046 3.3 0.00079038 3.3 0.00079048 0 0.0007904 0 0.0007905 3.3 0.00079042 3.3 0.00079052 0 0.00079044 0 0.00079054 3.3 0.00079046 3.3 0.0007905599999999999 0 0.0007904800000000001 0 0.00079058 3.3 0.0007905000000000001 3.3 0.0007906 0 0.0007905200000000001 0 0.00079062 3.3 0.0007905400000000001 3.3 0.00079064 0 0.00079056 0 0.00079066 3.3 0.00079058 3.3 0.00079068 0 0.0007906 0 0.0007907 3.3 0.00079062 3.3 0.00079072 0 0.00079064 0 0.00079074 3.3 0.00079066 3.3 0.0007907599999999999 0 0.00079068 0 0.0007907799999999999 3.3 0.0007907000000000001 3.3 0.0007908 0 0.0007907200000000001 0 0.00079082 3.3 0.0007907400000000001 3.3 0.00079084 0 0.00079076 0 0.00079086 3.3 0.00079078 3.3 0.00079088 0 0.0007908 0 0.0007909 3.3 0.00079082 3.3 0.00079092 0 0.00079084 0 0.00079094 3.3 0.00079086 3.3 0.00079096 0 0.00079088 0 0.0007909799999999999 3.3 0.0007909000000000001 3.3 0.000791 0 0.0007909200000000001 0 0.00079102 3.3 0.0007909400000000001 3.3 0.00079104 0 0.0007909600000000001 0 0.00079106 3.3 0.00079098 3.3 0.00079108 0 0.000791 0 0.0007911 3.3 0.00079102 3.3 0.00079112 0 0.00079104 0 0.00079114 3.3 0.00079106 3.3 0.00079116 0 0.00079108 0 0.0007911799999999999 3.3 0.0007911 3.3 0.0007911999999999999 0 0.0007911200000000001 0 0.00079122 3.3 0.0007911400000000001 3.3 0.00079124 0 0.0007911600000000001 0 0.00079126 3.3 0.00079118 3.3 0.00079128 0 0.0007912 0 0.0007913 3.3 0.00079122 3.3 0.00079132 0 0.00079124 0 0.00079134 3.3 0.00079126 3.3 0.00079136 0 0.00079128 0 0.00079138 3.3 0.0007913 3.3 0.0007913999999999999 0 0.0007913200000000001 0 0.00079142 3.3 0.0007913400000000001 3.3 0.00079144 0 0.0007913600000000001 0 0.00079146 3.3 0.0007913800000000001 3.3 0.00079148 0 0.0007914 0 0.0007915 3.3 0.00079142 3.3 0.00079152 0 0.00079144 0 0.00079154 3.3 0.00079146 3.3 0.00079156 0 0.00079148 0 0.00079158 3.3 0.0007915 3.3 0.0007915999999999999 0 0.00079152 0 0.0007916199999999999 3.3 0.0007915400000000001 3.3 0.00079164 0 0.0007915600000000001 0 0.00079166 3.3 0.0007915800000000001 3.3 0.00079168 0 0.0007916 0 0.0007917 3.3 0.00079162 3.3 0.00079172 0 0.00079164 0 0.00079174 3.3 0.00079166 3.3 0.00079176 0 0.00079168 0 0.00079178 3.3 0.0007917 3.3 0.0007918 0 0.00079172 0 0.0007918199999999999 3.3 0.0007917400000000001 3.3 0.00079184 0 0.0007917600000000001 0 0.00079186 3.3 0.0007917800000000001 3.3 0.00079188 0 0.0007918000000000001 0 0.0007919 3.3 0.00079182 3.3 0.00079192 0 0.00079184 0 0.00079194 3.3 0.00079186 3.3 0.00079196 0 0.00079188 0 0.00079198 3.3 0.0007919 3.3 0.000792 0 0.00079192 0 0.0007920199999999999 3.3 0.00079194 3.3 0.0007920399999999999 0 0.0007919600000000001 0 0.00079206 3.3 0.0007919800000000001 3.3 0.00079208 0 0.0007920000000000001 0 0.0007921 3.3 0.00079202 3.3 0.00079212 0 0.00079204 0 0.00079214 3.3 0.00079206 3.3 0.00079216 0 0.00079208 0 0.00079218 3.3 0.0007921 3.3 0.0007922 0 0.00079212 0 0.00079222 3.3 0.00079214 3.3 0.0007922399999999999 0 0.0007921600000000001 0 0.00079226 3.3 0.0007921800000000001 3.3 0.00079228 0 0.0007922000000000001 0 0.0007923 3.3 0.0007922200000000001 3.3 0.00079232 0 0.00079224 0 0.00079234 3.3 0.00079226 3.3 0.00079236 0 0.00079228 0 0.00079238 3.3 0.0007923 3.3 0.0007924 0 0.00079232 0 0.00079242 3.3 0.00079234 3.3 0.0007924399999999999 0 0.00079236 0 0.0007924599999999999 3.3 0.0007923800000000001 3.3 0.00079248 0 0.0007924000000000001 0 0.0007925 3.3 0.0007924200000000001 3.3 0.00079252 0 0.00079244 0 0.00079254 3.3 0.00079246 3.3 0.00079256 0 0.00079248 0 0.00079258 3.3 0.0007925 3.3 0.0007926 0 0.00079252 0 0.00079262 3.3 0.00079254 3.3 0.00079264 0 0.00079256 0 0.0007926599999999999 3.3 0.0007925800000000001 3.3 0.00079268 0 0.0007926000000000001 0 0.0007927 3.3 0.0007926200000000001 3.3 0.00079272 0 0.0007926400000000001 0 0.00079274 3.3 0.00079266 3.3 0.00079276 0 0.00079268 0 0.00079278 3.3 0.0007927 3.3 0.0007928 0 0.00079272 0 0.00079282 3.3 0.00079274 3.3 0.00079284 0 0.00079276 0 0.0007928599999999999 3.3 0.00079278 3.3 0.0007928799999999999 0 0.0007928000000000001 0 0.0007929 3.3 0.0007928200000000001 3.3 0.00079292 0 0.0007928400000000001 0 0.00079294 3.3 0.00079286 3.3 0.00079296 0 0.00079288 0 0.00079298 3.3 0.0007929 3.3 0.000793 0 0.00079292 0 0.00079302 3.3 0.00079294 3.3 0.00079304 0 0.00079296 0 0.0007930599999999999 3.3 0.00079298 3.3 0.0007930799999999999 0 0.0007930000000000001 0 0.0007931 3.3 0.0007930200000000001 3.3 0.00079312 0 0.0007930400000000001 0 0.00079314 3.3 0.00079306 3.3 0.00079316 0 0.00079308 0 0.00079318 3.3 0.0007931 3.3 0.0007932 0 0.00079312 0 0.00079322 3.3 0.00079314 3.3 0.00079324 0 0.00079316 0 0.00079326 3.3 0.00079318 3.3 0.0007932799999999999 0 0.0007932000000000001 0 0.0007933 3.3 0.0007932200000000001 3.3 0.00079332 0 0.0007932400000000001 0 0.00079334 3.3 0.0007932600000000001 3.3 0.00079336 0 0.00079328 0 0.00079338 3.3 0.0007933 3.3 0.0007934 0 0.00079332 0 0.00079342 3.3 0.00079334 3.3 0.00079344 0 0.00079336 0 0.00079346 3.3 0.00079338 3.3 0.0007934799999999999 0 0.0007934 0 0.0007934999999999999 3.3 0.0007934200000000001 3.3 0.00079352 0 0.0007934400000000001 0 0.00079354 3.3 0.0007934600000000001 3.3 0.00079356 0 0.00079348 0 0.00079358 3.3 0.0007935 3.3 0.0007936 0 0.00079352 0 0.00079362 3.3 0.00079354 3.3 0.00079364 0 0.00079356 0 0.00079366 3.3 0.00079358 3.3 0.00079368 0 0.0007936 0 0.0007936999999999999 3.3 0.0007936200000000001 3.3 0.00079372 0 0.0007936400000000001 0 0.00079374 3.3 0.0007936600000000001 3.3 0.00079376 0 0.0007936800000000001 0 0.00079378 3.3 0.0007937 3.3 0.0007938 0 0.00079372 0 0.00079382 3.3 0.00079374 3.3 0.00079384 0 0.00079376 0 0.00079386 3.3 0.00079378 3.3 0.00079388 0 0.0007938 0 0.0007938999999999999 3.3 0.00079382 3.3 0.0007939199999999999 0 0.0007938400000000001 0 0.00079394 3.3 0.0007938600000000001 3.3 0.00079396 0 0.0007938800000000001 0 0.00079398 3.3 0.0007939 3.3 0.000794 0 0.00079392 0 0.00079402 3.3 0.00079394 3.3 0.00079404 0 0.00079396 0 0.00079406 3.3 0.00079398 3.3 0.00079408 0 0.000794 0 0.0007941 3.3 0.00079402 3.3 0.0007941199999999999 0 0.0007940400000000001 0 0.00079414 3.3 0.0007940600000000001 3.3 0.00079416 0 0.0007940800000000001 0 0.00079418 3.3 0.0007941000000000001 3.3 0.0007942 0 0.00079412 0 0.00079422 3.3 0.00079414 3.3 0.00079424 0 0.00079416 0 0.00079426 3.3 0.00079418 3.3 0.00079428 0 0.0007942 0 0.0007943 3.3 0.00079422 3.3 0.0007943199999999999 0 0.00079424 0 0.0007943399999999999 3.3 0.0007942600000000001 3.3 0.00079436 0 0.0007942800000000001 0 0.00079438 3.3 0.0007943000000000001 3.3 0.0007944 0 0.00079432 0 0.00079442 3.3 0.00079434 3.3 0.00079444 0 0.00079436 0 0.00079446 3.3 0.00079438 3.3 0.00079448 0 0.0007944 0 0.0007945 3.3 0.00079442 3.3 0.00079452 0 0.00079444 0 0.0007945399999999999 3.3 0.0007944600000000001 3.3 0.00079456 0 0.0007944800000000001 0 0.00079458 3.3 0.0007945000000000001 3.3 0.0007946 0 0.0007945200000000001 0 0.00079462 3.3 0.00079454 3.3 0.00079464 0 0.00079456 0 0.00079466 3.3 0.00079458 3.3 0.00079468 0 0.0007946 0 0.0007947 3.3 0.00079462 3.3 0.00079472 0 0.00079464 0 0.0007947399999999999 3.3 0.00079466 3.3 0.0007947599999999999 0 0.0007946800000000001 0 0.00079478 3.3 0.0007947000000000001 3.3 0.0007948 0 0.0007947200000000001 0 0.00079482 3.3 0.00079474 3.3 0.00079484 0 0.00079476 0 0.00079486 3.3 0.00079478 3.3 0.00079488 0 0.0007948 0 0.0007949 3.3 0.00079482 3.3 0.00079492 0 0.00079484 0 0.00079494 3.3 0.00079486 3.3 0.0007949599999999999 0 0.0007948800000000001 0 0.00079498 3.3 0.0007949000000000001 3.3 0.000795 0 0.0007949200000000001 0 0.00079502 3.3 0.0007949400000000001 3.3 0.00079504 0 0.00079496 0 0.00079506 3.3 0.00079498 3.3 0.00079508 0 0.000795 0 0.0007951 3.3 0.00079502 3.3 0.00079512 0 0.00079504 0 0.00079514 3.3 0.00079506 3.3 0.0007951599999999999 0 0.00079508 0 0.0007951799999999999 3.3 0.0007951000000000001 3.3 0.0007952 0 0.0007951200000000001 0 0.00079522 3.3 0.0007951400000000001 3.3 0.00079524 0 0.00079516 0 0.00079526 3.3 0.00079518 3.3 0.00079528 0 0.0007952 0 0.0007953 3.3 0.00079522 3.3 0.00079532 0 0.00079524 0 0.00079534 3.3 0.00079526 3.3 0.00079536 0 0.00079528 0 0.0007953799999999999 3.3 0.0007953000000000001 3.3 0.0007954 0 0.0007953200000000001 0 0.00079542 3.3 0.0007953400000000001 3.3 0.00079544 0 0.0007953600000000001 0 0.00079546 3.3 0.00079538 3.3 0.00079548 0 0.0007954 0 0.0007955 3.3 0.00079542 3.3 0.00079552 0 0.00079544 0 0.00079554 3.3 0.00079546 3.3 0.00079556 0 0.00079548 0 0.0007955799999999999 3.3 0.0007955 3.3 0.0007955999999999999 0 0.0007955200000000001 0 0.00079562 3.3 0.0007955400000000001 3.3 0.00079564 0 0.0007955600000000001 0 0.00079566 3.3 0.00079558 3.3 0.00079568 0 0.0007956 0 0.0007957 3.3 0.00079562 3.3 0.00079572 0 0.00079564 0 0.00079574 3.3 0.00079566 3.3 0.00079576 0 0.00079568 0 0.00079578 3.3 0.0007957 3.3 0.0007957999999999999 0 0.0007957200000000001 0 0.00079582 3.3 0.0007957400000000001 3.3 0.00079584 0 0.0007957600000000001 0 0.00079586 3.3 0.0007957800000000001 3.3 0.00079588 0 0.0007958 0 0.0007959 3.3 0.00079582 3.3 0.00079592 0 0.00079584 0 0.00079594 3.3 0.00079586 3.3 0.00079596 0 0.00079588 0 0.00079598 3.3 0.0007959 3.3 0.0007959999999999999 0 0.00079592 0 0.0007960199999999999 3.3 0.0007959400000000001 3.3 0.00079604 0 0.0007959600000000001 0 0.00079606 3.3 0.0007959800000000001 3.3 0.00079608 0 0.000796 0 0.0007961 3.3 0.00079602 3.3 0.00079612 0 0.00079604 0 0.00079614 3.3 0.00079606 3.3 0.00079616 0 0.00079608 0 0.00079618 3.3 0.0007961 3.3 0.0007962 0 0.00079612 0 0.0007962199999999999 3.3 0.0007961400000000001 3.3 0.00079624 0 0.0007961600000000001 0 0.00079626 3.3 0.0007961800000000001 3.3 0.00079628 0 0.0007962000000000001 0 0.0007963 3.3 0.00079622 3.3 0.00079632 0 0.00079624 0 0.00079634 3.3 0.00079626 3.3 0.00079636 0 0.00079628 0 0.00079638 3.3 0.0007963 3.3 0.0007964 0 0.00079632 0 0.0007964199999999999 3.3 0.00079634 3.3 0.0007964399999999999 0 0.0007963600000000001 0 0.00079646 3.3 0.0007963800000000001 3.3 0.00079648 0 0.0007964000000000001 0 0.0007965 3.3 0.00079642 3.3 0.00079652 0 0.00079644 0 0.00079654 3.3 0.00079646 3.3 0.00079656 0 0.00079648 0 0.00079658 3.3 0.0007965 3.3 0.0007966 0 0.00079652 0 0.0007966199999999999 3.3 0.00079654 3.3 0.0007966399999999999 0 0.0007965600000000001 0 0.00079666 3.3 0.0007965800000000001 3.3 0.00079668 0 0.0007966000000000001 0 0.0007967 3.3 0.00079662 3.3 0.00079672 0 0.00079664 0 0.00079674 3.3 0.00079666 3.3 0.00079676 0 0.00079668 0 0.00079678 3.3 0.0007967 3.3 0.0007968 0 0.00079672 0 0.00079682 3.3 0.00079674 3.3 0.0007968399999999999 0 0.0007967600000000001 0 0.00079686 3.3 0.0007967800000000001 3.3 0.00079688 0 0.0007968000000000001 0 0.0007969 3.3 0.0007968200000000001 3.3 0.00079692 0 0.00079684 0 0.00079694 3.3 0.00079686 3.3 0.00079696 0 0.00079688 0 0.00079698 3.3 0.0007969 3.3 0.000797 0 0.00079692 0 0.00079702 3.3 0.00079694 3.3 0.0007970399999999999 0 0.00079696 0 0.0007970599999999999 3.3 0.0007969800000000001 3.3 0.00079708 0 0.0007970000000000001 0 0.0007971 3.3 0.0007970200000000001 3.3 0.00079712 0 0.00079704 0 0.00079714 3.3 0.00079706 3.3 0.00079716 0 0.00079708 0 0.00079718 3.3 0.0007971 3.3 0.0007972 0 0.00079712 0 0.00079722 3.3 0.00079714 3.3 0.00079724 0 0.00079716 0 0.0007972599999999999 3.3 0.0007971800000000001 3.3 0.00079728 0 0.0007972000000000001 0 0.0007973 3.3 0.0007972200000000001 3.3 0.00079732 0 0.0007972400000000001 0 0.00079734 3.3 0.00079726 3.3 0.00079736 0 0.00079728 0 0.00079738 3.3 0.0007973 3.3 0.0007974 0 0.00079732 0 0.00079742 3.3 0.00079734 3.3 0.00079744 0 0.00079736 0 0.0007974599999999999 3.3 0.00079738 3.3 0.0007974799999999999 0 0.0007974000000000001 0 0.0007975 3.3 0.0007974200000000001 3.3 0.00079752 0 0.0007974400000000001 0 0.00079754 3.3 0.00079746 3.3 0.00079756 0 0.00079748 0 0.00079758 3.3 0.0007975 3.3 0.0007976 0 0.00079752 0 0.00079762 3.3 0.00079754 3.3 0.00079764 0 0.00079756 0 0.00079766 3.3 0.00079758 3.3 0.0007976799999999999 0 0.0007976000000000001 0 0.0007977 3.3 0.0007976200000000001 3.3 0.00079772 0 0.0007976400000000001 0 0.00079774 3.3 0.0007976600000000001 3.3 0.00079776 0 0.00079768 0 0.00079778 3.3 0.0007977 3.3 0.0007978 0 0.00079772 0 0.00079782 3.3 0.00079774 3.3 0.00079784 0 0.00079776 0 0.00079786 3.3 0.00079778 3.3 0.0007978799999999999 0 0.0007978 0 0.0007978999999999999 3.3 0.0007978200000000001 3.3 0.00079792 0 0.0007978400000000001 0 0.00079794 3.3 0.0007978600000000001 3.3 0.00079796 0 0.00079788 0 0.00079798 3.3 0.0007979 3.3 0.000798 0 0.00079792 0 0.00079802 3.3 0.00079794 3.3 0.00079804 0 0.00079796 0 0.00079806 3.3 0.00079798 3.3 0.00079808 0 0.000798 0 0.0007980999999999999 3.3 0.0007980200000000001 3.3 0.00079812 0 0.0007980400000000001 0 0.00079814 3.3 0.0007980600000000001 3.3 0.00079816 0 0.0007980800000000001 0 0.00079818 3.3 0.0007981 3.3 0.0007982 0 0.00079812 0 0.00079822 3.3 0.00079814 3.3 0.00079824 0 0.00079816 0 0.00079826 3.3 0.00079818 3.3 0.00079828 0 0.0007982 0 0.0007982999999999999 3.3 0.00079822 3.3 0.0007983199999999999 0 0.0007982400000000001 0 0.00079834 3.3 0.0007982600000000001 3.3 0.00079836 0 0.0007982800000000001 0 0.00079838 3.3 0.0007983 3.3 0.0007984 0 0.00079832 0 0.00079842 3.3 0.00079834 3.3 0.00079844 0 0.00079836 0 0.00079846 3.3 0.00079838 3.3 0.00079848 0 0.0007984 0 0.0007985 3.3 0.00079842 3.3 0.0007985199999999999 0 0.0007984400000000001 0 0.00079854 3.3 0.0007984600000000001 3.3 0.00079856 0 0.0007984800000000001 0 0.00079858 3.3 0.0007985000000000001 3.3 0.0007986 0 0.00079852 0 0.00079862 3.3 0.00079854 3.3 0.00079864 0 0.00079856 0 0.00079866 3.3 0.00079858 3.3 0.00079868 0 0.0007986 0 0.0007987 3.3 0.00079862 3.3 0.0007987199999999999 0 0.00079864 0 0.0007987399999999999 3.3 0.0007986600000000001 3.3 0.00079876 0 0.0007986800000000001 0 0.00079878 3.3 0.0007987000000000001 3.3 0.0007988 0 0.00079872 0 0.00079882 3.3 0.00079874 3.3 0.00079884 0 0.00079876 0 0.00079886 3.3 0.00079878 3.3 0.00079888 0 0.0007988 0 0.0007989 3.3 0.00079882 3.3 0.00079892 0 0.00079884 0 0.0007989399999999999 3.3 0.0007988600000000001 3.3 0.00079896 0 0.0007988800000000001 0 0.00079898 3.3 0.0007989000000000001 3.3 0.000799 0 0.0007989200000000001 0 0.00079902 3.3 0.00079894 3.3 0.00079904 0 0.00079896 0 0.00079906 3.3 0.00079898 3.3 0.00079908 0 0.000799 0 0.0007991 3.3 0.00079902 3.3 0.00079912 0 0.00079904 0 0.0007991399999999999 3.3 0.00079906 3.3 0.0007991599999999999 0 0.0007990800000000001 0 0.00079918 3.3 0.0007991000000000001 3.3 0.0007992 0 0.0007991200000000001 0 0.00079922 3.3 0.00079914 3.3 0.00079924 0 0.00079916 0 0.00079926 3.3 0.00079918 3.3 0.00079928 0 0.0007992 0 0.0007993 3.3 0.00079922 3.3 0.00079932 0 0.00079924 0 0.00079934 3.3 0.00079926 3.3 0.0007993599999999999 0 0.0007992800000000001 0 0.00079938 3.3 0.0007993000000000001 3.3 0.0007994 0 0.0007993200000000001 0 0.00079942 3.3 0.0007993400000000001 3.3 0.00079944 0 0.00079936 0 0.00079946 3.3 0.00079938 3.3 0.00079948 0 0.0007994 0 0.0007995 3.3 0.00079942 3.3 0.00079952 0 0.00079944 0 0.00079954 3.3 0.00079946 3.3 0.0007995599999999999 0 0.00079948 0 0.0007995799999999999 3.3 0.0007995000000000001 3.3 0.0007996 0 0.0007995200000000001 0 0.00079962 3.3 0.0007995400000000001 3.3 0.00079964 0 0.00079956 0 0.00079966 3.3 0.00079958 3.3 0.00079968 0 0.0007996 0 0.0007997 3.3 0.00079962 3.3 0.00079972 0 0.00079964 0 0.00079974 3.3 0.00079966 3.3 0.0007997599999999999 0 0.00079968 0 0.0007997799999999999 3.3 0.0007997000000000001 3.3 0.0007998 0 0.0007997200000000001 0 0.00079982 3.3 0.0007997400000000001 3.3 0.00079984 0 0.00079976 0 0.00079986 3.3 0.00079978 3.3 0.00079988 0 0.0007998 0 0.0007999 3.3 0.00079982 3.3 0.00079992 0 0.00079984 0 0.00079994 3.3 0.00079986 3.3 0.00079996 0 0.00079988 0 0.0007999799999999999 3.3 0.0007999 3.3 0.0007999999999999999 0 0.0007999200000000001 0 0.00080002 3.3 0.0007999400000000001 3.3 0.00080004 0 0.0007999600000000001 0 0.00080006 3.3 0.00079998 3.3 0.00080008 0 0.0008 0 0.0008001 3.3 0.00080002 3.3 0.00080012 0 0.00080004 0 0.00080014 3.3 0.00080006 3.3 0.00080016 0 0.00080008 0 0.0008001799999999999 3.3 0.0008001 3.3 0.0008001999999999999 0 0.0008001200000000001 0 0.00080022 3.3 0.0008001400000000001 3.3 0.00080024 0 0.0008001600000000001 0 0.00080026 3.3 0.00080018 3.3 0.00080028 0 0.0008002 0 0.0008003 3.3 0.00080022 3.3 0.00080032 0 0.00080024 0 0.00080034 3.3 0.00080026 3.3 0.00080036 0 0.00080028 0 0.00080038 3.3 0.0008003 3.3 0.0008003999999999999 0 0.0008003200000000001 0 0.00080042 3.3 0.0008003400000000001 3.3 0.00080044 0 0.0008003600000000001 0 0.00080046 3.3 0.0008003800000000001 3.3 0.00080048 0 0.0008004 0 0.0008005 3.3 0.00080042 3.3 0.00080052 0 0.00080044 0 0.00080054 3.3 0.00080046 3.3 0.00080056 0 0.00080048 0 0.00080058 3.3 0.0008005 3.3 0.0008005999999999999 0 0.00080052 0 0.0008006199999999999 3.3 0.0008005400000000001 3.3 0.00080064 0 0.0008005600000000001 0 0.00080066 3.3 0.0008005800000000001 3.3 0.00080068 0 0.0008006 0 0.0008007 3.3 0.00080062 3.3 0.00080072 0 0.00080064 0 0.00080074 3.3 0.00080066 3.3 0.00080076 0 0.00080068 0 0.00080078 3.3 0.0008007 3.3 0.0008008 0 0.00080072 0 0.0008008199999999999 3.3 0.0008007400000000001 3.3 0.00080084 0 0.0008007600000000001 0 0.00080086 3.3 0.0008007800000000001 3.3 0.00080088 0 0.0008008000000000001 0 0.0008009 3.3 0.00080082 3.3 0.00080092 0 0.00080084 0 0.00080094 3.3 0.00080086 3.3 0.00080096 0 0.00080088 0 0.00080098 3.3 0.0008009 3.3 0.000801 0 0.00080092 0 0.0008010199999999999 3.3 0.00080094 3.3 0.0008010399999999999 0 0.0008009600000000001 0 0.00080106 3.3 0.0008009800000000001 3.3 0.00080108 0 0.0008010000000000001 0 0.0008011 3.3 0.00080102 3.3 0.00080112 0 0.00080104 0 0.00080114 3.3 0.00080106 3.3 0.00080116 0 0.00080108 0 0.00080118 3.3 0.0008011 3.3 0.0008012 0 0.00080112 0 0.00080122 3.3 0.00080114 3.3 0.0008012399999999999 0 0.0008011600000000001 0 0.00080126 3.3 0.0008011800000000001 3.3 0.00080128 0 0.0008012000000000001 0 0.0008013 3.3 0.0008012200000000001 3.3 0.00080132 0 0.00080124 0 0.00080134 3.3 0.00080126 3.3 0.00080136 0 0.00080128 0 0.00080138 3.3 0.0008013 3.3 0.0008014 0 0.00080132 0 0.00080142 3.3 0.00080134 3.3 0.0008014399999999999 0 0.00080136 0 0.0008014599999999999 3.3 0.0008013800000000001 3.3 0.00080148 0 0.0008014000000000001 0 0.0008015 3.3 0.0008014200000000001 3.3 0.00080152 0 0.00080144 0 0.00080154 3.3 0.00080146 3.3 0.00080156 0 0.00080148 0 0.00080158 3.3 0.0008015 3.3 0.0008016 0 0.00080152 0 0.00080162 3.3 0.00080154 3.3 0.00080164 0 0.00080156 0 0.0008016599999999999 3.3 0.0008015800000000001 3.3 0.00080168 0 0.0008016000000000001 0 0.0008017 3.3 0.0008016200000000001 3.3 0.00080172 0 0.0008016400000000001 0 0.00080174 3.3 0.00080166 3.3 0.00080176 0 0.00080168 0 0.00080178 3.3 0.0008017 3.3 0.0008018 0 0.00080172 0 0.00080182 3.3 0.00080174 3.3 0.00080184 0 0.00080176 0 0.0008018599999999999 3.3 0.00080178 3.3 0.0008018799999999999 0 0.0008018000000000001 0 0.0008019 3.3 0.0008018200000000001 3.3 0.00080192 0 0.0008018400000000001 0 0.00080194 3.3 0.00080186 3.3 0.00080196 0 0.00080188 0 0.00080198 3.3 0.0008019 3.3 0.000802 0 0.00080192 0 0.00080202 3.3 0.00080194 3.3 0.00080204 0 0.00080196 0 0.00080206 3.3 0.00080198 3.3 0.0008020799999999999 0 0.0008020000000000001 0 0.0008021 3.3 0.0008020200000000001 3.3 0.00080212 0 0.0008020400000000001 0 0.00080214 3.3 0.0008020600000000001 3.3 0.00080216 0 0.00080208 0 0.00080218 3.3 0.0008021 3.3 0.0008022 0 0.00080212 0 0.00080222 3.3 0.00080214 3.3 0.00080224 0 0.00080216 0 0.00080226 3.3 0.00080218 3.3 0.0008022799999999999 0 0.0008022 0 0.0008022999999999999 3.3 0.0008022200000000001 3.3 0.00080232 0 0.0008022400000000001 0 0.00080234 3.3 0.0008022600000000001 3.3 0.00080236 0 0.00080228 0 0.00080238 3.3 0.0008023 3.3 0.0008024 0 0.00080232 0 0.00080242 3.3 0.00080234 3.3 0.00080244 0 0.00080236 0 0.00080246 3.3 0.00080238 3.3 0.00080248 0 0.0008024 0 0.0008024999999999999 3.3 0.0008024200000000001 3.3 0.00080252 0 0.0008024400000000001 0 0.00080254 3.3 0.0008024600000000001 3.3 0.00080256 0 0.0008024800000000001 0 0.00080258 3.3 0.0008025 3.3 0.0008026 0 0.00080252 0 0.00080262 3.3 0.00080254 3.3 0.00080264 0 0.00080256 0 0.00080266 3.3 0.00080258 3.3 0.00080268 0 0.0008026 0 0.0008026999999999999 3.3 0.00080262 3.3 0.0008027199999999999 0 0.0008026400000000001 0 0.00080274 3.3 0.0008026600000000001 3.3 0.00080276 0 0.0008026800000000001 0 0.00080278 3.3 0.0008027 3.3 0.0008028 0 0.00080272 0 0.00080282 3.3 0.00080274 3.3 0.00080284 0 0.00080276 0 0.00080286 3.3 0.00080278 3.3 0.00080288 0 0.0008028 0 0.0008029 3.3 0.00080282 3.3 0.0008029199999999999 0 0.0008028400000000001 0 0.00080294 3.3 0.0008028600000000001 3.3 0.00080296 0 0.0008028800000000001 0 0.00080298 3.3 0.0008029000000000001 3.3 0.000803 0 0.00080292 0 0.00080302 3.3 0.00080294 3.3 0.00080304 0 0.00080296 0 0.00080306 3.3 0.00080298 3.3 0.00080308 0 0.000803 0 0.0008031 3.3 0.00080302 3.3 0.0008031199999999999 0 0.00080304 0 0.0008031399999999999 3.3 0.0008030600000000001 3.3 0.00080316 0 0.0008030800000000001 0 0.00080318 3.3 0.0008031000000000001 3.3 0.0008032 0 0.00080312 0 0.00080322 3.3 0.00080314 3.3 0.00080324 0 0.00080316 0 0.00080326 3.3 0.00080318 3.3 0.00080328 0 0.0008032 0 0.0008033 3.3 0.00080322 3.3 0.0008033199999999999 0 0.00080324 0 0.0008033399999999999 3.3 0.0008032600000000001 3.3 0.00080336 0 0.0008032800000000001 0 0.00080338 3.3 0.0008033000000000001 3.3 0.0008034 0 0.00080332 0 0.00080342 3.3 0.00080334 3.3 0.00080344 0 0.00080336 0 0.00080346 3.3 0.00080338 3.3 0.00080348 0 0.0008034 0 0.0008035 3.3 0.00080342 3.3 0.00080352 0 0.00080344 0 0.0008035399999999999 3.3 0.00080346 3.3 0.0008035599999999999 0 0.0008034800000000001 0 0.00080358 3.3 0.0008035000000000001 3.3 0.0008036 0 0.0008035200000000001 0 0.00080362 3.3 0.00080354 3.3 0.00080364 0 0.00080356 0 0.00080366 3.3 0.00080358 3.3 0.00080368 0 0.0008036 0 0.0008037 3.3 0.00080362 3.3 0.00080372 0 0.00080364 0 0.0008037399999999999 3.3 0.00080366 3.3 0.0008037599999999999 0 0.0008036800000000001 0 0.00080378 3.3 0.0008037000000000001 3.3 0.0008038 0 0.0008037200000000001 0 0.00080382 3.3 0.00080374 3.3 0.00080384 0 0.00080376 0 0.00080386 3.3 0.00080378 3.3 0.00080388 0 0.0008038 0 0.0008039 3.3 0.00080382 3.3 0.00080392 0 0.00080384 0 0.00080394 3.3 0.00080386 3.3 0.0008039599999999999 0 0.0008038800000000001 0 0.00080398 3.3 0.0008039000000000001 3.3 0.000804 0 0.0008039200000000001 0 0.00080402 3.3 0.0008039400000000001 3.3 0.00080404 0 0.00080396 0 0.00080406 3.3 0.00080398 3.3 0.00080408 0 0.000804 0 0.0008041 3.3 0.00080402 3.3 0.00080412 0 0.00080404 0 0.00080414 3.3 0.00080406 3.3 0.0008041599999999999 0 0.00080408 0 0.0008041799999999999 3.3 0.0008041000000000001 3.3 0.0008042 0 0.0008041200000000001 0 0.00080422 3.3 0.0008041400000000001 3.3 0.00080424 0 0.00080416 0 0.00080426 3.3 0.00080418 3.3 0.00080428 0 0.0008042 0 0.0008043 3.3 0.00080422 3.3 0.00080432 0 0.00080424 0 0.00080434 3.3 0.00080426 3.3 0.00080436 0 0.00080428 0 0.0008043799999999999 3.3 0.0008043000000000001 3.3 0.0008044 0 0.0008043200000000001 0 0.00080442 3.3 0.0008043400000000001 3.3 0.00080444 0 0.0008043600000000001 0 0.00080446 3.3 0.00080438 3.3 0.00080448 0 0.0008044 0 0.0008045 3.3 0.00080442 3.3 0.00080452 0 0.00080444 0 0.00080454 3.3 0.00080446 3.3 0.00080456 0 0.00080448 0 0.0008045799999999999 3.3 0.0008045 3.3 0.0008045999999999999 0 0.0008045200000000001 0 0.00080462 3.3 0.0008045400000000001 3.3 0.00080464 0 0.0008045600000000001 0 0.00080466 3.3 0.00080458 3.3 0.00080468 0 0.0008046 0 0.0008047 3.3 0.00080462 3.3 0.00080472 0 0.00080464 0 0.00080474 3.3 0.00080466 3.3 0.00080476 0 0.00080468 0 0.00080478 3.3 0.0008047 3.3 0.0008047999999999999 0 0.0008047200000000001 0 0.00080482 3.3 0.0008047400000000001 3.3 0.00080484 0 0.0008047600000000001 0 0.00080486 3.3 0.0008047800000000001 3.3 0.00080488 0 0.0008048 0 0.0008049 3.3 0.00080482 3.3 0.00080492 0 0.00080484 0 0.00080494 3.3 0.00080486 3.3 0.00080496 0 0.00080488 0 0.00080498 3.3 0.0008049 3.3 0.0008049999999999999 0 0.00080492 0 0.0008050199999999999 3.3 0.0008049400000000001 3.3 0.00080504 0 0.0008049600000000001 0 0.00080506 3.3 0.0008049800000000001 3.3 0.00080508 0 0.000805 0 0.0008051 3.3 0.00080502 3.3 0.00080512 0 0.00080504 0 0.00080514 3.3 0.00080506 3.3 0.00080516 0 0.00080508 0 0.00080518 3.3 0.0008051 3.3 0.0008052 0 0.00080512 0 0.0008052199999999999 3.3 0.0008051400000000001 3.3 0.00080524 0 0.0008051600000000001 0 0.00080526 3.3 0.0008051800000000001 3.3 0.00080528 0 0.0008052000000000001 0 0.0008053 3.3 0.00080522 3.3 0.00080532 0 0.00080524 0 0.00080534 3.3 0.00080526 3.3 0.00080536 0 0.00080528 0 0.00080538 3.3 0.0008053 3.3 0.0008054 0 0.00080532 0 0.0008054199999999999 3.3 0.00080534 3.3 0.0008054399999999999 0 0.0008053600000000001 0 0.00080546 3.3 0.0008053800000000001 3.3 0.00080548 0 0.0008054000000000001 0 0.0008055 3.3 0.00080542 3.3 0.00080552 0 0.00080544 0 0.00080554 3.3 0.00080546 3.3 0.00080556 0 0.00080548 0 0.00080558 3.3 0.0008055 3.3 0.0008056 0 0.00080552 0 0.00080562 3.3 0.00080554 3.3 0.0008056399999999999 0 0.0008055600000000001 0 0.00080566 3.3 0.0008055800000000001 3.3 0.00080568 0 0.0008056000000000001 0 0.0008057 3.3 0.0008056200000000001 3.3 0.00080572 0 0.00080564 0 0.00080574 3.3 0.00080566 3.3 0.00080576 0 0.00080568 0 0.00080578 3.3 0.0008057 3.3 0.0008058 0 0.00080572 0 0.00080582 3.3 0.00080574 3.3 0.0008058399999999999 0 0.00080576 0 0.0008058599999999999 3.3 0.0008057800000000001 3.3 0.00080588 0 0.0008058000000000001 0 0.0008059 3.3 0.0008058200000000001 3.3 0.00080592 0 0.00080584 0 0.00080594 3.3 0.00080586 3.3 0.00080596 0 0.00080588 0 0.00080598 3.3 0.0008059 3.3 0.000806 0 0.00080592 0 0.00080602 3.3 0.00080594 3.3 0.00080604 0 0.00080596 0 0.0008060599999999999 3.3 0.0008059800000000001 3.3 0.00080608 0 0.0008060000000000001 0 0.0008061 3.3 0.0008060200000000001 3.3 0.00080612 0 0.0008060400000000001 0 0.00080614 3.3 0.00080606 3.3 0.00080616 0 0.00080608 0 0.00080618 3.3 0.0008061 3.3 0.0008062 0 0.00080612 0 0.00080622 3.3 0.00080614 3.3 0.00080624 0 0.00080616 0 0.0008062599999999999 3.3 0.00080618 3.3 0.0008062799999999999 0 0.0008062000000000001 0 0.0008063 3.3 0.0008062200000000001 3.3 0.00080632 0 0.0008062400000000001 0 0.00080634 3.3 0.00080626 3.3 0.00080636 0 0.00080628 0 0.00080638 3.3 0.0008063 3.3 0.0008064 0 0.00080632 0 0.00080642 3.3 0.00080634 3.3 0.00080644 0 0.00080636 0 0.00080646 3.3 0.00080638 3.3 0.0008064799999999999 0 0.0008064000000000001 0 0.0008065 3.3 0.0008064200000000001 3.3 0.00080652 0 0.0008064400000000001 0 0.00080654 3.3 0.0008064600000000001 3.3 0.00080656 0 0.00080648 0 0.00080658 3.3 0.0008065 3.3 0.0008066 0 0.00080652 0 0.00080662 3.3 0.00080654 3.3 0.00080664 0 0.00080656 0 0.00080666 3.3 0.00080658 3.3 0.0008066799999999999 0 0.0008066 0 0.0008066999999999999 3.3 0.0008066200000000001 3.3 0.00080672 0 0.0008066400000000001 0 0.00080674 3.3 0.0008066600000000001 3.3 0.00080676 0 0.00080668 0 0.00080678 3.3 0.0008067 3.3 0.0008068 0 0.00080672 0 0.00080682 3.3 0.00080674 3.3 0.00080684 0 0.00080676 0 0.00080686 3.3 0.00080678 3.3 0.0008068799999999999 0 0.0008068 0 0.0008068999999999999 3.3 0.0008068200000000001 3.3 0.00080692 0 0.0008068400000000001 0 0.00080694 3.3 0.0008068600000000001 3.3 0.00080696 0 0.00080688 0 0.00080698 3.3 0.0008069 3.3 0.000807 0 0.00080692 0 0.00080702 3.3 0.00080694 3.3 0.00080704 0 0.00080696 0 0.00080706 3.3 0.00080698 3.3 0.00080708 0 0.000807 0 0.0008070999999999999 3.3 0.0008070200000000001 3.3 0.00080712 0 0.0008070400000000001 0 0.00080714 3.3 0.0008070600000000001 3.3 0.00080716 0 0.0008070800000000001 0 0.00080718 3.3 0.0008071 3.3 0.0008072 0 0.00080712 0 0.00080722 3.3 0.00080714 3.3 0.00080724 0 0.00080716 0 0.00080726 3.3 0.00080718 3.3 0.00080728 0 0.0008072 0 0.0008072999999999999 3.3 0.00080722 3.3 0.0008073199999999999 0 0.0008072400000000001 0 0.00080734 3.3 0.0008072600000000001 3.3 0.00080736 0 0.0008072800000000001 0 0.00080738 3.3 0.0008073 3.3 0.0008074 0 0.00080732 0 0.00080742 3.3 0.00080734 3.3 0.00080744 0 0.00080736 0 0.00080746 3.3 0.00080738 3.3 0.00080748 0 0.0008074 0 0.0008075 3.3 0.00080742 3.3 0.0008075199999999999 0 0.0008074400000000001 0 0.00080754 3.3 0.0008074600000000001 3.3 0.00080756 0 0.0008074800000000001 0 0.00080758 3.3 0.0008075000000000001 3.3 0.0008076 0 0.00080752 0 0.00080762 3.3 0.00080754 3.3 0.00080764 0 0.00080756 0 0.00080766 3.3 0.00080758 3.3 0.00080768 0 0.0008076 0 0.0008077 3.3 0.00080762 3.3 0.0008077199999999999 0 0.00080764 0 0.0008077399999999999 3.3 0.0008076600000000001 3.3 0.00080776 0 0.0008076800000000001 0 0.00080778 3.3 0.0008077000000000001 3.3 0.0008078 0 0.00080772 0 0.00080782 3.3 0.00080774 3.3 0.00080784 0 0.00080776 0 0.00080786 3.3 0.00080778 3.3 0.00080788 0 0.0008078 0 0.0008079 3.3 0.00080782 3.3 0.00080792 0 0.00080784 0 0.0008079399999999999 3.3 0.0008078600000000001 3.3 0.00080796 0 0.0008078800000000001 0 0.00080798 3.3 0.0008079000000000001 3.3 0.000808 0 0.0008079200000000001 0 0.00080802 3.3 0.00080794 3.3 0.00080804 0 0.00080796 0 0.00080806 3.3 0.00080798 3.3 0.00080808 0 0.000808 0 0.0008081 3.3 0.00080802 3.3 0.00080812 0 0.00080804 0 0.0008081399999999999 3.3 0.00080806 3.3 0.0008081599999999999 0 0.0008080800000000001 0 0.00080818 3.3 0.0008081000000000001 3.3 0.0008082 0 0.0008081200000000001 0 0.00080822 3.3 0.00080814 3.3 0.00080824 0 0.00080816 0 0.00080826 3.3 0.00080818 3.3 0.00080828 0 0.0008082 0 0.0008083 3.3 0.00080822 3.3 0.00080832 0 0.00080824 0 0.00080834 3.3 0.00080826 3.3 0.0008083599999999999 0 0.0008082800000000001 0 0.00080838 3.3 0.0008083000000000001 3.3 0.0008084 0 0.0008083200000000001 0 0.00080842 3.3 0.0008083400000000001 3.3 0.00080844 0 0.00080836 0 0.00080846 3.3 0.00080838 3.3 0.00080848 0 0.0008084 0 0.0008085 3.3 0.00080842 3.3 0.00080852 0 0.00080844 0 0.00080854 3.3 0.00080846 3.3 0.0008085599999999999 0 0.00080848 0 0.0008085799999999999 3.3 0.0008085000000000001 3.3 0.0008086 0 0.0008085200000000001 0 0.00080862 3.3 0.0008085400000000001 3.3 0.00080864 0 0.00080856 0 0.00080866 3.3 0.00080858 3.3 0.00080868 0 0.0008086 0 0.0008087 3.3 0.00080862 3.3 0.00080872 0 0.00080864 0 0.00080874 3.3 0.00080866 3.3 0.00080876 0 0.00080868 0 0.0008087799999999999 3.3 0.0008087000000000001 3.3 0.0008088 0 0.0008087200000000001 0 0.00080882 3.3 0.0008087400000000001 3.3 0.00080884 0 0.0008087600000000001 0 0.00080886 3.3 0.00080878 3.3 0.00080888 0 0.0008088 0 0.0008089 3.3 0.00080882 3.3 0.00080892 0 0.00080884 0 0.00080894 3.3 0.00080886 3.3 0.00080896 0 0.00080888 0 0.0008089799999999999 3.3 0.0008089 3.3 0.0008089999999999999 0 0.0008089200000000001 0 0.00080902 3.3 0.0008089400000000001 3.3 0.00080904 0 0.0008089600000000001 0 0.00080906 3.3 0.00080898 3.3 0.00080908 0 0.000809 0 0.0008091 3.3 0.00080902 3.3 0.00080912 0 0.00080904 0 0.00080914 3.3 0.00080906 3.3 0.00080916 0 0.00080908 0 0.00080918 3.3 0.0008091 3.3 0.0008091999999999999 0 0.0008091200000000001 0 0.00080922 3.3 0.0008091400000000001 3.3 0.00080924 0 0.0008091600000000001 0 0.00080926 3.3 0.0008091800000000001 3.3 0.00080928 0 0.0008092 0 0.0008093 3.3 0.00080922 3.3 0.00080932 0 0.00080924 0 0.00080934 3.3 0.00080926 3.3 0.00080936 0 0.00080928 0 0.00080938 3.3 0.0008093 3.3 0.0008093999999999999 0 0.00080932 0 0.0008094199999999999 3.3 0.0008093400000000001 3.3 0.00080944 0 0.0008093600000000001 0 0.00080946 3.3 0.0008093800000000001 3.3 0.00080948 0 0.0008094 0 0.0008095 3.3 0.00080942 3.3 0.00080952 0 0.00080944 0 0.00080954 3.3 0.00080946 3.3 0.00080956 0 0.00080948 0 0.00080958 3.3 0.0008095 3.3 0.0008096 0 0.00080952 0 0.0008096199999999999 3.3 0.0008095400000000001 3.3 0.00080964 0 0.0008095600000000001 0 0.00080966 3.3 0.0008095800000000001 3.3 0.00080968 0 0.0008096000000000001 0 0.0008097 3.3 0.00080962 3.3 0.00080972 0 0.00080964 0 0.00080974 3.3 0.00080966 3.3 0.00080976 0 0.00080968 0 0.00080978 3.3 0.0008097 3.3 0.0008098 0 0.00080972 0 0.0008098199999999999 3.3 0.00080974 3.3 0.0008098399999999999 0 0.0008097600000000001 0 0.00080986 3.3 0.0008097800000000001 3.3 0.00080988 0 0.0008098000000000001 0 0.0008099 3.3 0.00080982 3.3 0.00080992 0 0.00080984 0 0.00080994 3.3 0.00080986 3.3 0.00080996 0 0.00080988 0 0.00080998 3.3 0.0008099 3.3 0.00081 0 0.00080992 0 0.00081002 3.3 0.00080994 3.3 0.0008100399999999999 0 0.0008099600000000001 0 0.00081006 3.3 0.0008099800000000001 3.3 0.00081008 0 0.0008100000000000001 0 0.0008101 3.3 0.0008100200000000001 3.3 0.00081012 0 0.00081004 0 0.00081014 3.3 0.00081006 3.3 0.00081016 0 0.00081008 0 0.00081018 3.3 0.0008101 3.3 0.0008102 0 0.00081012 0 0.00081022 3.3 0.00081014 3.3 0.0008102399999999999 0 0.00081016 0 0.0008102599999999999 3.3 0.0008101800000000001 3.3 0.00081028 0 0.0008102000000000001 0 0.0008103 3.3 0.0008102200000000001 3.3 0.00081032 0 0.00081024 0 0.00081034 3.3 0.00081026 3.3 0.00081036 0 0.00081028 0 0.00081038 3.3 0.0008103 3.3 0.0008104 0 0.00081032 0 0.00081042 3.3 0.00081034 3.3 0.0008104399999999999 0 0.00081036 0 0.0008104599999999999 3.3 0.0008103800000000001 3.3 0.00081048 0 0.0008104000000000001 0 0.0008105 3.3 0.0008104200000000001 3.3 0.00081052 0 0.00081044 0 0.00081054 3.3 0.00081046 3.3 0.00081056 0 0.00081048 0 0.00081058 3.3 0.0008105 3.3 0.0008106 0 0.00081052 0 0.00081062 3.3 0.00081054 3.3 0.00081064 0 0.00081056 0 0.0008106599999999999 3.3 0.0008105800000000001 3.3 0.00081068 0 0.0008106000000000001 0 0.0008107 3.3 0.0008106200000000001 3.3 0.00081072 0 0.0008106400000000001 0 0.00081074 3.3 0.00081066 3.3 0.00081076 0 0.00081068 0 0.00081078 3.3 0.0008107 3.3 0.0008108 0 0.00081072 0 0.00081082 3.3 0.00081074 3.3 0.00081084 0 0.00081076 0 0.0008108599999999999 3.3 0.00081078 3.3 0.0008108799999999999 0 0.0008108000000000001 0 0.0008109 3.3 0.0008108200000000001 3.3 0.00081092 0 0.0008108400000000001 0 0.00081094 3.3 0.00081086 3.3 0.00081096 0 0.00081088 0 0.00081098 3.3 0.0008109 3.3 0.000811 0 0.00081092 0 0.00081102 3.3 0.00081094 3.3 0.00081104 0 0.00081096 0 0.00081106 3.3 0.00081098 3.3 0.0008110799999999999 0 0.0008110000000000001 0 0.0008111 3.3 0.0008110200000000001 3.3 0.00081112 0 0.0008110400000000001 0 0.00081114 3.3 0.0008110600000000001 3.3 0.00081116 0 0.00081108 0 0.00081118 3.3 0.0008111 3.3 0.0008112 0 0.00081112 0 0.00081122 3.3 0.00081114 3.3 0.00081124 0 0.00081116 0 0.00081126 3.3 0.00081118 3.3 0.0008112799999999999 0 0.0008112 0 0.0008112999999999999 3.3 0.0008112200000000001 3.3 0.00081132 0 0.0008112400000000001 0 0.00081134 3.3 0.0008112600000000001 3.3 0.00081136 0 0.00081128 0 0.00081138 3.3 0.0008113 3.3 0.0008114 0 0.00081132 0 0.00081142 3.3 0.00081134 3.3 0.00081144 0 0.00081136 0 0.00081146 3.3 0.00081138 3.3 0.00081148 0 0.0008114 0 0.0008114999999999999 3.3 0.0008114200000000001 3.3 0.00081152 0 0.0008114400000000001 0 0.00081154 3.3 0.0008114600000000001 3.3 0.00081156 0 0.0008114800000000001 0 0.00081158 3.3 0.0008115 3.3 0.0008116 0 0.00081152 0 0.00081162 3.3 0.00081154 3.3 0.00081164 0 0.00081156 0 0.00081166 3.3 0.00081158 3.3 0.00081168 0 0.0008116 0 0.0008116999999999999 3.3 0.00081162 3.3 0.0008117199999999999 0 0.0008116400000000001 0 0.00081174 3.3 0.0008116600000000001 3.3 0.00081176 0 0.0008116800000000001 0 0.00081178 3.3 0.0008117 3.3 0.0008118 0 0.00081172 0 0.00081182 3.3 0.00081174 3.3 0.00081184 0 0.00081176 0 0.00081186 3.3 0.00081178 3.3 0.00081188 0 0.0008118 0 0.0008119 3.3 0.00081182 3.3 0.0008119199999999999 0 0.0008118400000000001 0 0.00081194 3.3 0.0008118600000000001 3.3 0.00081196 0 0.0008118800000000001 0 0.00081198 3.3 0.0008119000000000001 3.3 0.000812 0 0.00081192 0 0.00081202 3.3 0.00081194 3.3 0.00081204 0 0.00081196 0 0.00081206 3.3 0.00081198 3.3 0.00081208 0 0.000812 0 0.0008121 3.3 0.00081202 3.3 0.0008121199999999999 0 0.00081204 0 0.0008121399999999999 3.3 0.0008120600000000001 3.3 0.00081216 0 0.0008120800000000001 0 0.00081218 3.3 0.0008121000000000001 3.3 0.0008122 0 0.00081212 0 0.00081222 3.3 0.00081214 3.3 0.00081224 0 0.00081216 0 0.00081226 3.3 0.00081218 3.3 0.00081228 0 0.0008122 0 0.0008123 3.3 0.00081222 3.3 0.00081232 0 0.00081224 0 0.0008123399999999999 3.3 0.0008122600000000001 3.3 0.00081236 0 0.0008122800000000001 0 0.00081238 3.3 0.0008123000000000001 3.3 0.0008124 0 0.0008123200000000001 0 0.00081242 3.3 0.00081234 3.3 0.00081244 0 0.00081236 0 0.00081246 3.3 0.00081238 3.3 0.00081248 0 0.0008124 0 0.0008125 3.3 0.00081242 3.3 0.00081252 0 0.00081244 0 0.0008125399999999999 3.3 0.00081246 3.3 0.0008125599999999999 0 0.0008124800000000001 0 0.00081258 3.3 0.0008125000000000001 3.3 0.0008126 0 0.0008125200000000001 0 0.00081262 3.3 0.00081254 3.3 0.00081264 0 0.00081256 0 0.00081266 3.3 0.00081258 3.3 0.00081268 0 0.0008126 0 0.0008127 3.3 0.00081262 3.3 0.00081272 0 0.00081264 0 0.00081274 3.3 0.00081266 3.3 0.0008127599999999999 0 0.0008126800000000001 0 0.00081278 3.3 0.0008127000000000001 3.3 0.0008128 0 0.0008127200000000001 0 0.00081282 3.3 0.0008127400000000001 3.3 0.00081284 0 0.00081276 0 0.00081286 3.3 0.00081278 3.3 0.00081288 0 0.0008128 0 0.0008129 3.3 0.00081282 3.3 0.00081292 0 0.00081284 0 0.00081294 3.3 0.00081286 3.3 0.0008129599999999999 0 0.00081288 0 0.0008129799999999999 3.3 0.0008129000000000001 3.3 0.000813 0 0.0008129200000000001 0 0.00081302 3.3 0.0008129400000000001 3.3 0.00081304 0 0.00081296 0 0.00081306 3.3 0.00081298 3.3 0.00081308 0 0.000813 0 0.0008131 3.3 0.00081302 3.3 0.00081312 0 0.00081304 0 0.00081314 3.3 0.00081306 3.3 0.00081316 0 0.00081308 0 0.0008131799999999999 3.3 0.0008131000000000001 3.3 0.0008132 0 0.0008131200000000001 0 0.00081322 3.3 0.0008131400000000001 3.3 0.00081324 0 0.0008131600000000001 0 0.00081326 3.3 0.00081318 3.3 0.00081328 0 0.0008132 0 0.0008133 3.3 0.00081322 3.3 0.00081332 0 0.00081324 0 0.00081334 3.3 0.00081326 3.3 0.00081336 0 0.00081328 0 0.0008133799999999999 3.3 0.0008133 3.3 0.0008133999999999999 0 0.0008133200000000001 0 0.00081342 3.3 0.0008133400000000001 3.3 0.00081344 0 0.0008133600000000001 0 0.00081346 3.3 0.00081338 3.3 0.00081348 0 0.0008134 0 0.0008135 3.3 0.00081342 3.3 0.00081352 0 0.00081344 0 0.00081354 3.3 0.00081346 3.3 0.00081356 0 0.00081348 0 0.0008135799999999999 3.3 0.0008135 3.3 0.0008135999999999999 0 0.0008135200000000001 0 0.00081362 3.3 0.0008135400000000001 3.3 0.00081364 0 0.0008135600000000001 0 0.00081366 3.3 0.00081358 3.3 0.00081368 0 0.0008136 0 0.0008137 3.3 0.00081362 3.3 0.00081372 0 0.00081364 0 0.00081374 3.3 0.00081366 3.3 0.00081376 0 0.00081368 0 0.00081378 3.3 0.0008137 3.3 0.0008137999999999999 0 0.00081372 0 0.0008138199999999999 3.3 0.0008137400000000001 3.3 0.00081384 0 0.0008137600000000001 0 0.00081386 3.3 0.0008137800000000001 3.3 0.00081388 0 0.0008138 0 0.0008139 3.3 0.00081382 3.3 0.00081392 0 0.00081384 0 0.00081394 3.3 0.00081386 3.3 0.00081396 0 0.00081388 0 0.00081398 3.3 0.0008139 3.3 0.0008139999999999999 0 0.00081392 0 0.0008140199999999999 3.3 0.0008139400000000001 3.3 0.00081404 0 0.0008139600000000001 0 0.00081406 3.3 0.0008139800000000001 3.3 0.00081408 0 0.000814 0 0.0008141 3.3 0.00081402 3.3 0.00081412 0 0.00081404 0 0.00081414 3.3 0.00081406 3.3 0.00081416 0 0.00081408 0 0.00081418 3.3 0.0008141 3.3 0.0008142 0 0.00081412 0 0.0008142199999999999 3.3 0.0008141400000000001 3.3 0.00081424 0 0.0008141600000000001 0 0.00081426 3.3 0.0008141800000000001 3.3 0.00081428 0 0.0008142000000000001 0 0.0008143 3.3 0.00081422 3.3 0.00081432 0 0.00081424 0 0.00081434 3.3 0.00081426 3.3 0.00081436 0 0.00081428 0 0.00081438 3.3 0.0008143 3.3 0.0008144 0 0.00081432 0 0.0008144199999999999 3.3 0.00081434 3.3 0.0008144399999999999 0 0.0008143600000000001 0 0.00081446 3.3 0.0008143800000000001 3.3 0.00081448 0 0.0008144000000000001 0 0.0008145 3.3 0.00081442 3.3 0.00081452 0 0.00081444 0 0.00081454 3.3 0.00081446 3.3 0.00081456 0 0.00081448 0 0.00081458 3.3 0.0008145 3.3 0.0008146 0 0.00081452 0 0.00081462 3.3 0.00081454 3.3 0.0008146399999999999 0 0.0008145600000000001 0 0.00081466 3.3 0.0008145800000000001 3.3 0.00081468 0 0.0008146000000000001 0 0.0008147 3.3 0.0008146200000000001 3.3 0.00081472 0 0.00081464 0 0.00081474 3.3 0.00081466 3.3 0.00081476 0 0.00081468 0 0.00081478 3.3 0.0008147 3.3 0.0008148 0 0.00081472 0 0.00081482 3.3 0.00081474 3.3 0.0008148399999999999 0 0.00081476 0 0.0008148599999999999 3.3 0.0008147800000000001 3.3 0.00081488 0 0.0008148000000000001 0 0.0008149 3.3 0.0008148200000000001 3.3 0.00081492 0 0.00081484 0 0.00081494 3.3 0.00081486 3.3 0.00081496 0 0.00081488 0 0.00081498 3.3 0.0008149 3.3 0.000815 0 0.00081492 0 0.00081502 3.3 0.00081494 3.3 0.00081504 0 0.00081496 0 0.0008150599999999999 3.3 0.0008149800000000001 3.3 0.00081508 0 0.0008150000000000001 0 0.0008151 3.3 0.0008150200000000001 3.3 0.00081512 0 0.0008150400000000001 0 0.00081514 3.3 0.00081506 3.3 0.00081516 0 0.00081508 0 0.00081518 3.3 0.0008151 3.3 0.0008152 0 0.00081512 0 0.00081522 3.3 0.00081514 3.3 0.00081524 0 0.00081516 0 0.0008152599999999999 3.3 0.00081518 3.3 0.0008152799999999999 0 0.0008152000000000001 0 0.0008153 3.3 0.0008152200000000001 3.3 0.00081532 0 0.0008152400000000001 0 0.00081534 3.3 0.00081526 3.3 0.00081536 0 0.00081528 0 0.00081538 3.3 0.0008153 3.3 0.0008154 0 0.00081532 0 0.00081542 3.3 0.00081534 3.3 0.00081544 0 0.00081536 0 0.00081546 3.3 0.00081538 3.3 0.0008154799999999999 0 0.0008154000000000001 0 0.0008155 3.3 0.0008154200000000001 3.3 0.00081552 0 0.0008154400000000001 0 0.00081554 3.3 0.0008154600000000001 3.3 0.00081556 0 0.00081548 0 0.00081558 3.3 0.0008155 3.3 0.0008156 0 0.00081552 0 0.00081562 3.3 0.00081554 3.3 0.00081564 0 0.00081556 0 0.00081566 3.3 0.00081558 3.3 0.0008156799999999999 0 0.0008156 0 0.0008156999999999999 3.3 0.0008156200000000001 3.3 0.00081572 0 0.0008156400000000001 0 0.00081574 3.3 0.0008156600000000001 3.3 0.00081576 0 0.00081568 0 0.00081578 3.3 0.0008157 3.3 0.0008158 0 0.00081572 0 0.00081582 3.3 0.00081574 3.3 0.00081584 0 0.00081576 0 0.00081586 3.3 0.00081578 3.3 0.00081588 0 0.0008158 0 0.0008158999999999999 3.3 0.0008158200000000001 3.3 0.00081592 0 0.0008158400000000001 0 0.00081594 3.3 0.0008158600000000001 3.3 0.00081596 0 0.0008158800000000001 0 0.00081598 3.3 0.0008159 3.3 0.000816 0 0.00081592 0 0.00081602 3.3 0.00081594 3.3 0.00081604 0 0.00081596 0 0.00081606 3.3 0.00081598 3.3 0.00081608 0 0.000816 0 0.0008160999999999999 3.3 0.00081602 3.3 0.0008161199999999999 0 0.0008160400000000001 0 0.00081614 3.3 0.0008160600000000001 3.3 0.00081616 0 0.0008160800000000001 0 0.00081618 3.3 0.0008161 3.3 0.0008162 0 0.00081612 0 0.00081622 3.3 0.00081614 3.3 0.00081624 0 0.00081616 0 0.00081626 3.3 0.00081618 3.3 0.00081628 0 0.0008162 0 0.0008163 3.3 0.00081622 3.3 0.0008163199999999999 0 0.0008162400000000001 0 0.00081634 3.3 0.0008162600000000001 3.3 0.00081636 0 0.0008162800000000001 0 0.00081638 3.3 0.0008163000000000001 3.3 0.0008164 0 0.00081632 0 0.00081642 3.3 0.00081634 3.3 0.00081644 0 0.00081636 0 0.00081646 3.3 0.00081638 3.3 0.00081648 0 0.0008164 0 0.0008165 3.3 0.00081642 3.3 0.0008165199999999999 0 0.00081644 0 0.0008165399999999999 3.3 0.0008164600000000001 3.3 0.00081656 0 0.0008164800000000001 0 0.00081658 3.3 0.0008165000000000001 3.3 0.0008166 0 0.00081652 0 0.00081662 3.3 0.00081654 3.3 0.00081664 0 0.00081656 0 0.00081666 3.3 0.00081658 3.3 0.00081668 0 0.0008166 0 0.0008167 3.3 0.00081662 3.3 0.00081672 0 0.00081664 0 0.0008167399999999999 3.3 0.0008166600000000001 3.3 0.00081676 0 0.0008166800000000001 0 0.00081678 3.3 0.0008167000000000001 3.3 0.0008168 0 0.0008167200000000001 0 0.00081682 3.3 0.00081674 3.3 0.00081684 0 0.00081676 0 0.00081686 3.3 0.00081678 3.3 0.00081688 0 0.0008168 0 0.0008169 3.3 0.00081682 3.3 0.00081692 0 0.00081684 0 0.0008169399999999999 3.3 0.00081686 3.3 0.0008169599999999999 0 0.0008168800000000001 0 0.00081698 3.3 0.0008169000000000001 3.3 0.000817 0 0.0008169200000000001 0 0.00081702 3.3 0.00081694 3.3 0.00081704 0 0.00081696 0 0.00081706 3.3 0.00081698 3.3 0.00081708 0 0.000817 0 0.0008171 3.3 0.00081702 3.3 0.00081712 0 0.00081704 0 0.0008171399999999999 3.3 0.00081706 3.3 0.0008171599999999999 0 0.0008170800000000001 0 0.00081718 3.3 0.0008171000000000001 3.3 0.0008172 0 0.0008171200000000001 0 0.00081722 3.3 0.00081714 3.3 0.00081724 0 0.00081716 0 0.00081726 3.3 0.00081718 3.3 0.00081728 0 0.0008172 0 0.0008173 3.3 0.00081722 3.3 0.00081732 0 0.00081724 0 0.00081734 3.3 0.00081726 3.3 0.0008173599999999999 0 0.00081728 0 0.0008173799999999999 3.3 0.0008173000000000001 3.3 0.0008174 0 0.0008173200000000001 0 0.00081742 3.3 0.0008173400000000001 3.3 0.00081744 0 0.00081736 0 0.00081746 3.3 0.00081738 3.3 0.00081748 0 0.0008174 0 0.0008175 3.3 0.00081742 3.3 0.00081752 0 0.00081744 0 0.00081754 3.3 0.00081746 3.3 0.0008175599999999999 0 0.00081748 0 0.0008175799999999999 3.3 0.0008175000000000001 3.3 0.0008176 0 0.0008175200000000001 0 0.00081762 3.3 0.0008175400000000001 3.3 0.00081764 0 0.00081756 0 0.00081766 3.3 0.00081758 3.3 0.00081768 0 0.0008176 0 0.0008177 3.3 0.00081762 3.3 0.00081772 0 0.00081764 0 0.00081774 3.3 0.00081766 3.3 0.00081776 0 0.00081768 0 0.0008177799999999999 3.3 0.0008177000000000001 3.3 0.0008178 0 0.0008177200000000001 0 0.00081782 3.3 0.0008177400000000001 3.3 0.00081784 0 0.0008177600000000001 0 0.00081786 3.3 0.00081778 3.3 0.00081788 0 0.0008178 0 0.0008179 3.3 0.00081782 3.3 0.00081792 0 0.00081784 0 0.00081794 3.3 0.00081786 3.3 0.00081796 0 0.00081788 0 0.0008179799999999999 3.3 0.0008179 3.3 0.0008179999999999999 0 0.0008179200000000001 0 0.00081802 3.3 0.0008179400000000001 3.3 0.00081804 0 0.0008179600000000001 0 0.00081806 3.3 0.00081798 3.3 0.00081808 0 0.000818 0 0.0008181 3.3 0.00081802 3.3 0.00081812 0 0.00081804 0 0.00081814 3.3 0.00081806 3.3 0.00081816 0 0.00081808 0 0.00081818 3.3 0.0008181 3.3 0.0008181999999999999 0 0.0008181200000000001 0 0.00081822 3.3 0.0008181400000000001 3.3 0.00081824 0 0.0008181600000000001 0 0.00081826 3.3 0.0008181800000000001 3.3 0.00081828 0 0.0008182 0 0.0008183 3.3 0.00081822 3.3 0.00081832 0 0.00081824 0 0.00081834 3.3 0.00081826 3.3 0.00081836 0 0.00081828 0 0.00081838 3.3 0.0008183 3.3 0.0008183999999999999 0 0.00081832 0 0.0008184199999999999 3.3 0.0008183400000000001 3.3 0.00081844 0 0.0008183600000000001 0 0.00081846 3.3 0.0008183800000000001 3.3 0.00081848 0 0.0008184 0 0.0008185 3.3 0.00081842 3.3 0.00081852 0 0.00081844 0 0.00081854 3.3 0.00081846 3.3 0.00081856 0 0.00081848 0 0.00081858 3.3 0.0008185 3.3 0.0008186 0 0.00081852 0 0.0008186199999999999 3.3 0.0008185400000000001 3.3 0.00081864 0 0.0008185600000000001 0 0.00081866 3.3 0.0008185800000000001 3.3 0.00081868 0 0.0008186000000000001 0 0.0008187 3.3 0.00081862 3.3 0.00081872 0 0.00081864 0 0.00081874 3.3 0.00081866 3.3 0.00081876 0 0.00081868 0 0.00081878 3.3 0.0008187 3.3 0.0008188 0 0.00081872 0 0.0008188199999999999 3.3 0.00081874 3.3 0.0008188399999999999 0 0.0008187600000000001 0 0.00081886 3.3 0.0008187800000000001 3.3 0.00081888 0 0.0008188000000000001 0 0.0008189 3.3 0.00081882 3.3 0.00081892 0 0.00081884 0 0.00081894 3.3 0.00081886 3.3 0.00081896 0 0.00081888 0 0.00081898 3.3 0.0008189 3.3 0.000819 0 0.00081892 0 0.00081902 3.3 0.00081894 3.3 0.0008190399999999999 0 0.0008189600000000001 0 0.00081906 3.3 0.0008189800000000001 3.3 0.00081908 0 0.0008190000000000001 0 0.0008191 3.3 0.0008190200000000001 3.3 0.00081912 0 0.00081904 0 0.00081914 3.3 0.00081906 3.3 0.00081916 0 0.00081908 0 0.00081918 3.3 0.0008191 3.3 0.0008192 0 0.00081912 0 0.00081922 3.3 0.00081914 3.3 0.0008192399999999999 0 0.00081916 0 0.0008192599999999999 3.3 0.0008191800000000001 3.3 0.00081928 0 0.0008192000000000001 0 0.0008193 3.3 0.0008192200000000001 3.3 0.00081932 0 0.00081924 0 0.00081934 3.3 0.00081926 3.3 0.00081936 0 0.00081928 0 0.00081938 3.3 0.0008193 3.3 0.0008194 0 0.00081932 0 0.00081942 3.3 0.00081934 3.3 0.00081944 0 0.00081936 0 0.0008194599999999999 3.3 0.0008193800000000001 3.3 0.00081948 0 0.0008194000000000001 0 0.0008195 3.3 0.0008194200000000001 3.3 0.00081952 0 0.0008194400000000001 0 0.00081954 3.3 0.00081946 3.3 0.00081956 0 0.00081948 0 0.00081958 3.3 0.0008195 3.3 0.0008196 0 0.00081952 0 0.00081962 3.3 0.00081954 3.3 0.00081964 0 0.00081956 0 0.0008196599999999999 3.3 0.00081958 3.3 0.0008196799999999999 0 0.0008196000000000001 0 0.0008197 3.3 0.0008196200000000001 3.3 0.00081972 0 0.0008196400000000001 0 0.00081974 3.3 0.00081966 3.3 0.00081976 0 0.00081968 0 0.00081978 3.3 0.0008197 3.3 0.0008198 0 0.00081972 0 0.00081982 3.3 0.00081974 3.3 0.00081984 0 0.00081976 0 0.00081986 3.3 0.00081978 3.3 0.0008198799999999999 0 0.0008198000000000001 0 0.0008199 3.3 0.0008198200000000001 3.3 0.00081992 0 0.0008198400000000001 0 0.00081994 3.3 0.0008198600000000001 3.3 0.00081996 0 0.00081988 0 0.00081998 3.3 0.0008199 3.3 0.00082 0 0.00081992 0 0.00082002 3.3 0.00081994 3.3 0.00082004 0 0.00081996 0 0.00082006 3.3 0.00081998 3.3 0.0008200799999999999 0 0.00082 0 0.0008200999999999999 3.3 0.0008200200000000001 3.3 0.00082012 0 0.0008200400000000001 0 0.00082014 3.3 0.0008200600000000001 3.3 0.00082016 0 0.00082008 0 0.00082018 3.3 0.0008201 3.3 0.0008202 0 0.00082012 0 0.00082022 3.3 0.00082014 3.3 0.00082024 0 0.00082016 0 0.00082026 3.3 0.00082018 3.3 0.00082028 0 0.0008202 0 0.0008202999999999999 3.3 0.0008202200000000001 3.3 0.00082032 0 0.0008202400000000001 0 0.00082034 3.3 0.0008202600000000001 3.3 0.00082036 0 0.0008202800000000001 0 0.00082038 3.3 0.0008203 3.3 0.0008204 0 0.00082032 0 0.00082042 3.3 0.00082034 3.3 0.00082044 0 0.00082036 0 0.00082046 3.3 0.00082038 3.3 0.00082048 0 0.0008204 0 0.0008204999999999999 3.3 0.00082042 3.3 0.0008205199999999999 0 0.0008204400000000001 0 0.00082054 3.3 0.0008204600000000001 3.3 0.00082056 0 0.0008204800000000001 0 0.00082058 3.3 0.0008205 3.3 0.0008206 0 0.00082052 0 0.00082062 3.3 0.00082054 3.3 0.00082064 0 0.00082056 0 0.00082066 3.3 0.00082058 3.3 0.00082068 0 0.0008206 0 0.0008206999999999999 3.3 0.00082062 3.3 0.0008207199999999999 0 0.0008206400000000001 0 0.00082074 3.3 0.0008206600000000001 3.3 0.00082076 0 0.0008206800000000001 0 0.00082078 3.3 0.0008207 3.3 0.0008208 0 0.00082072 0 0.00082082 3.3 0.00082074 3.3 0.00082084 0 0.00082076 0 0.00082086 3.3 0.00082078 3.3 0.00082088 0 0.0008208 0 0.0008209 3.3 0.00082082 3.3 0.0008209199999999999 0 0.00082084 0 0.0008209399999999999 3.3 0.0008208600000000001 3.3 0.00082096 0 0.0008208800000000001 0 0.00082098 3.3 0.0008209000000000001 3.3 0.000821 0 0.00082092 0 0.00082102 3.3 0.00082094 3.3 0.00082104 0 0.00082096 0 0.00082106 3.3 0.00082098 3.3 0.00082108 0 0.000821 0 0.0008211 3.3 0.00082102 3.3 0.0008211199999999999 0 0.00082104 0 0.0008211399999999999 3.3 0.0008210600000000001 3.3 0.00082116 0 0.0008210800000000001 0 0.00082118 3.3 0.0008211000000000001 3.3 0.0008212 0 0.00082112 0 0.00082122 3.3 0.00082114 3.3 0.00082124 0 0.00082116 0 0.00082126 3.3 0.00082118 3.3 0.00082128 0 0.0008212 0 0.0008213 3.3 0.00082122 3.3 0.00082132 0 0.00082124 0 0.0008213399999999999 3.3 0.0008212600000000001 3.3 0.00082136 0 0.0008212800000000001 0 0.00082138 3.3 0.0008213000000000001 3.3 0.0008214 0 0.0008213200000000001 0 0.00082142 3.3 0.00082134 3.3 0.00082144 0 0.00082136 0 0.00082146 3.3 0.00082138 3.3 0.00082148 0 0.0008214 0 0.0008215 3.3 0.00082142 3.3 0.00082152 0 0.00082144 0 0.0008215399999999999 3.3 0.00082146 3.3 0.0008215599999999999 0 0.0008214800000000001 0 0.00082158 3.3 0.0008215000000000001 3.3 0.0008216 0 0.0008215200000000001 0 0.00082162 3.3 0.00082154 3.3 0.00082164 0 0.00082156 0 0.00082166 3.3 0.00082158 3.3 0.00082168 0 0.0008216 0 0.0008217 3.3 0.00082162 3.3 0.00082172 0 0.00082164 0 0.00082174 3.3 0.00082166 3.3 0.0008217599999999999 0 0.0008216800000000001 0 0.00082178 3.3 0.0008217000000000001 3.3 0.0008218 0 0.0008217200000000001 0 0.00082182 3.3 0.0008217400000000001 3.3 0.00082184 0 0.00082176 0 0.00082186 3.3 0.00082178 3.3 0.00082188 0 0.0008218 0 0.0008219 3.3 0.00082182 3.3 0.00082192 0 0.00082184 0 0.00082194 3.3 0.00082186 3.3 0.0008219599999999999 0 0.00082188 0 0.0008219799999999999 3.3 0.0008219000000000001 3.3 0.000822 0 0.0008219200000000001 0 0.00082202 3.3 0.0008219400000000001 3.3 0.00082204 0 0.00082196 0 0.00082206 3.3 0.00082198 3.3 0.00082208 0 0.000822 0 0.0008221 3.3 0.00082202 3.3 0.00082212 0 0.00082204 0 0.00082214 3.3 0.00082206 3.3 0.00082216 0 0.00082208 0 0.0008221799999999999 3.3 0.0008221000000000001 3.3 0.0008222 0 0.0008221200000000001 0 0.00082222 3.3 0.0008221400000000001 3.3 0.00082224 0 0.0008221600000000001 0 0.00082226 3.3 0.00082218 3.3 0.00082228 0 0.0008222 0 0.0008223 3.3 0.00082222 3.3 0.00082232 0 0.00082224 0 0.00082234 3.3 0.00082226 3.3 0.00082236 0 0.00082228 0 0.0008223799999999999 3.3 0.0008223 3.3 0.0008223999999999999 0 0.0008223200000000001 0 0.00082242 3.3 0.0008223400000000001 3.3 0.00082244 0 0.0008223600000000001 0 0.00082246 3.3 0.00082238 3.3 0.00082248 0 0.0008224 0 0.0008225 3.3 0.00082242 3.3 0.00082252 0 0.00082244 0 0.00082254 3.3 0.00082246 3.3 0.00082256 0 0.00082248 0 0.00082258 3.3 0.0008225 3.3 0.0008225999999999999 0 0.0008225200000000001 0 0.00082262 3.3 0.0008225400000000001 3.3 0.00082264 0 0.0008225600000000001 0 0.00082266 3.3 0.0008225800000000001 3.3 0.00082268 0 0.0008226 0 0.0008227 3.3 0.00082262 3.3 0.00082272 0 0.00082264 0 0.00082274 3.3 0.00082266 3.3 0.00082276 0 0.00082268 0 0.00082278 3.3 0.0008227 3.3 0.0008227999999999999 0 0.00082272 0 0.0008228199999999999 3.3 0.0008227400000000001 3.3 0.00082284 0 0.0008227600000000001 0 0.00082286 3.3 0.0008227800000000001 3.3 0.00082288 0 0.0008228 0 0.0008229 3.3 0.00082282 3.3 0.00082292 0 0.00082284 0 0.00082294 3.3 0.00082286 3.3 0.00082296 0 0.00082288 0 0.00082298 3.3 0.0008229 3.3 0.000823 0 0.00082292 0 0.0008230199999999999 3.3 0.0008229400000000001 3.3 0.00082304 0 0.0008229600000000001 0 0.00082306 3.3 0.0008229800000000001 3.3 0.00082308 0 0.0008230000000000001 0 0.0008231 3.3 0.00082302 3.3 0.00082312 0 0.00082304 0 0.00082314 3.3 0.00082306 3.3 0.00082316 0 0.00082308 0 0.00082318 3.3 0.0008231 3.3 0.0008232 0 0.00082312 0 0.0008232199999999999 3.3 0.00082314 3.3 0.0008232399999999999 0 0.0008231600000000001 0 0.00082326 3.3 0.0008231800000000001 3.3 0.00082328 0 0.0008232000000000001 0 0.0008233 3.3 0.00082322 3.3 0.00082332 0 0.00082324 0 0.00082334 3.3 0.00082326 3.3 0.00082336 0 0.00082328 0 0.00082338 3.3 0.0008233 3.3 0.0008234 0 0.00082332 0 0.00082342 3.3 0.00082334 3.3 0.0008234399999999999 0 0.0008233600000000001 0 0.00082346 3.3 0.0008233800000000001 3.3 0.00082348 0 0.0008234000000000001 0 0.0008235 3.3 0.0008234200000000001 3.3 0.00082352 0 0.00082344 0 0.00082354 3.3 0.00082346 3.3 0.00082356 0 0.00082348 0 0.00082358 3.3 0.0008235 3.3 0.0008236 0 0.00082352 0 0.00082362 3.3 0.00082354 3.3 0.0008236399999999999 0 0.00082356 0 0.0008236599999999999 3.3 0.0008235800000000001 3.3 0.00082368 0 0.0008236000000000001 0 0.0008237 3.3 0.0008236200000000001 3.3 0.00082372 0 0.00082364 0 0.00082374 3.3 0.00082366 3.3 0.00082376 0 0.00082368 0 0.00082378 3.3 0.0008237 3.3 0.0008238 0 0.00082372 0 0.00082382 3.3 0.00082374 3.3 0.0008238399999999999 0 0.00082376 0 0.0008238599999999999 3.3 0.0008237800000000001 3.3 0.00082388 0 0.0008238000000000001 0 0.0008239 3.3 0.0008238200000000001 3.3 0.00082392 0 0.00082384 0 0.00082394 3.3 0.00082386 3.3 0.00082396 0 0.00082388 0 0.00082398 3.3 0.0008239 3.3 0.000824 0 0.00082392 0 0.00082402 3.3 0.00082394 3.3 0.00082404 0 0.00082396 0 0.0008240599999999999 3.3 0.00082398 3.3 0.0008240799999999999 0 0.0008240000000000001 0 0.0008241 3.3 0.0008240200000000001 3.3 0.00082412 0 0.0008240400000000001 0 0.00082414 3.3 0.00082406 3.3 0.00082416 0 0.00082408 0 0.00082418 3.3 0.0008241 3.3 0.0008242 0 0.00082412 0 0.00082422 3.3 0.00082414 3.3 0.00082424 0 0.00082416 0 0.0008242599999999999 3.3 0.00082418 3.3 0.0008242799999999999 0 0.0008242000000000001 0 0.0008243 3.3 0.0008242200000000001 3.3 0.00082432 0 0.0008242400000000001 0 0.00082434 3.3 0.00082426 3.3 0.00082436 0 0.00082428 0 0.00082438 3.3 0.0008243 3.3 0.0008244 0 0.00082432 0 0.00082442 3.3 0.00082434 3.3 0.00082444 0 0.00082436 0 0.00082446 3.3 0.00082438 3.3 0.0008244799999999999 0 0.0008244000000000001 0 0.0008245 3.3 0.0008244200000000001 3.3 0.00082452 0 0.0008244400000000001 0 0.00082454 3.3 0.0008244600000000001 3.3 0.00082456 0 0.00082448 0 0.00082458 3.3 0.0008245 3.3 0.0008246 0 0.00082452 0 0.00082462 3.3 0.00082454 3.3 0.00082464 0 0.00082456 0 0.00082466 3.3 0.00082458 3.3 0.0008246799999999999 0 0.0008246 0 0.0008246999999999999 3.3 0.0008246200000000001 3.3 0.00082472 0 0.0008246400000000001 0 0.00082474 3.3 0.0008246600000000001 3.3 0.00082476 0 0.00082468 0 0.00082478 3.3 0.0008247 3.3 0.0008248 0 0.00082472 0 0.00082482 3.3 0.00082474 3.3 0.00082484 0 0.00082476 0 0.00082486 3.3 0.00082478 3.3 0.00082488 0 0.0008248 0 0.0008248999999999999 3.3 0.0008248200000000001 3.3 0.00082492 0 0.0008248400000000001 0 0.00082494 3.3 0.0008248600000000001 3.3 0.00082496 0 0.0008248800000000001 0 0.00082498 3.3 0.0008249 3.3 0.000825 0 0.00082492 0 0.00082502 3.3 0.00082494 3.3 0.00082504 0 0.00082496 0 0.00082506 3.3 0.00082498 3.3 0.00082508 0 0.000825 0 0.0008250999999999999 3.3 0.00082502 3.3 0.0008251199999999999 0 0.0008250400000000001 0 0.00082514 3.3 0.0008250600000000001 3.3 0.00082516 0 0.0008250800000000001 0 0.00082518 3.3 0.0008251 3.3 0.0008252 0 0.00082512 0 0.00082522 3.3 0.00082514 3.3 0.00082524 0 0.00082516 0 0.00082526 3.3 0.00082518 3.3 0.00082528 0 0.0008252 0 0.0008253 3.3 0.00082522 3.3 0.0008253199999999999 0 0.0008252400000000001 0 0.00082534 3.3 0.0008252600000000001 3.3 0.00082536 0 0.0008252800000000001 0 0.00082538 3.3 0.0008253000000000001 3.3 0.0008254 0 0.00082532 0 0.00082542 3.3 0.00082534 3.3 0.00082544 0 0.00082536 0 0.00082546 3.3 0.00082538 3.3 0.00082548 0 0.0008254 0 0.0008255 3.3 0.00082542 3.3 0.0008255199999999999 0 0.00082544 0 0.0008255399999999999 3.3 0.0008254600000000001 3.3 0.00082556 0 0.0008254800000000001 0 0.00082558 3.3 0.0008255000000000001 3.3 0.0008256 0 0.00082552 0 0.00082562 3.3 0.00082554 3.3 0.00082564 0 0.00082556 0 0.00082566 3.3 0.00082558 3.3 0.00082568 0 0.0008256 0 0.0008257 3.3 0.00082562 3.3 0.00082572 0 0.00082564 0 0.0008257399999999999 3.3 0.0008256600000000001 3.3 0.00082576 0 0.0008256800000000001 0 0.00082578 3.3 0.0008257000000000001 3.3 0.0008258 0 0.0008257200000000001 0 0.00082582 3.3 0.00082574 3.3 0.00082584 0 0.00082576 0 0.00082586 3.3 0.00082578 3.3 0.00082588 0 0.0008258 0 0.0008259 3.3 0.00082582 3.3 0.00082592 0 0.00082584 0 0.0008259399999999999 3.3 0.00082586 3.3 0.0008259599999999999 0 0.0008258800000000001 0 0.00082598 3.3 0.0008259000000000001 3.3 0.000826 0 0.0008259200000000001 0 0.00082602 3.3 0.00082594 3.3 0.00082604 0 0.00082596 0 0.00082606 3.3 0.00082598 3.3 0.00082608 0 0.000826 0 0.0008261 3.3 0.00082602 3.3 0.00082612 0 0.00082604 0 0.00082614 3.3 0.00082606 3.3 0.0008261599999999999 0 0.0008260800000000001 0 0.00082618 3.3 0.0008261000000000001 3.3 0.0008262 0 0.0008261200000000001 0 0.00082622 3.3 0.0008261400000000001 3.3 0.00082624 0 0.00082616 0 0.00082626 3.3 0.00082618 3.3 0.00082628 0 0.0008262 0 0.0008263 3.3 0.00082622 3.3 0.00082632 0 0.00082624 0 0.00082634 3.3 0.00082626 3.3 0.0008263599999999999 0 0.00082628 0 0.0008263799999999999 3.3 0.0008263000000000001 3.3 0.0008264 0 0.0008263200000000001 0 0.00082642 3.3 0.0008263400000000001 3.3 0.00082644 0 0.00082636 0 0.00082646 3.3 0.00082638 3.3 0.00082648 0 0.0008264 0 0.0008265 3.3 0.00082642 3.3 0.00082652 0 0.00082644 0 0.00082654 3.3 0.00082646 3.3 0.00082656 0 0.00082648 0 0.0008265799999999999 3.3 0.0008265000000000001 3.3 0.0008266 0 0.0008265200000000001 0 0.00082662 3.3 0.0008265400000000001 3.3 0.00082664 0 0.0008265600000000001 0 0.00082666 3.3 0.00082658 3.3 0.00082668 0 0.0008266 0 0.0008267 3.3 0.00082662 3.3 0.00082672 0 0.00082664 0 0.00082674 3.3 0.00082666 3.3 0.00082676 0 0.00082668 0 0.0008267799999999999 3.3 0.0008267 3.3 0.0008267999999999999 0 0.0008267200000000001 0 0.00082682 3.3 0.0008267400000000001 3.3 0.00082684 0 0.0008267600000000001 0 0.00082686 3.3 0.00082678 3.3 0.00082688 0 0.0008268 0 0.0008269 3.3 0.00082682 3.3 0.00082692 0 0.00082684 0 0.00082694 3.3 0.00082686 3.3 0.00082696 0 0.00082688 0 0.00082698 3.3 0.0008269 3.3 0.0008269999999999999 0 0.0008269200000000001 0 0.00082702 3.3 0.0008269400000000001 3.3 0.00082704 0 0.0008269600000000001 0 0.00082706 3.3 0.0008269800000000001 3.3 0.00082708 0 0.000827 0 0.0008271 3.3 0.00082702 3.3 0.00082712 0 0.00082704 0 0.00082714 3.3 0.00082706 3.3 0.00082716 0 0.00082708 0 0.00082718 3.3 0.0008271 3.3 0.0008271999999999999 0 0.00082712 0 0.0008272199999999999 3.3 0.0008271400000000001 3.3 0.00082724 0 0.0008271600000000001 0 0.00082726 3.3 0.0008271800000000001 3.3 0.00082728 0 0.0008272 0 0.0008273 3.3 0.00082722 3.3 0.00082732 0 0.00082724 0 0.00082734 3.3 0.00082726 3.3 0.00082736 0 0.00082728 0 0.00082738 3.3 0.0008273 3.3 0.0008273999999999999 0 0.00082732 0 0.0008274199999999999 3.3 0.0008273400000000001 3.3 0.00082744 0 0.0008273600000000001 0 0.00082746 3.3 0.0008273800000000001 3.3 0.00082748 0 0.0008274 0 0.0008275 3.3 0.00082742 3.3 0.00082752 0 0.00082744 0 0.00082754 3.3 0.00082746 3.3 0.00082756 0 0.00082748 0 0.00082758 3.3 0.0008275 3.3 0.0008276 0 0.00082752 0 0.0008276199999999999 3.3 0.00082754 3.3 0.0008276399999999999 0 0.0008275600000000001 0 0.00082766 3.3 0.0008275800000000001 3.3 0.00082768 0 0.0008276000000000001 0 0.0008277 3.3 0.00082762 3.3 0.00082772 0 0.00082764 0 0.00082774 3.3 0.00082766 3.3 0.00082776 0 0.00082768 0 0.00082778 3.3 0.0008277 3.3 0.0008278 0 0.00082772 0 0.0008278199999999999 3.3 0.00082774 3.3 0.0008278399999999999 0 0.0008277600000000001 0 0.00082786 3.3 0.0008277800000000001 3.3 0.00082788 0 0.0008278000000000001 0 0.0008279 3.3 0.00082782 3.3 0.00082792 0 0.00082784 0 0.00082794 3.3 0.00082786 3.3 0.00082796 0 0.00082788 0 0.00082798 3.3 0.0008279 3.3 0.000828 0 0.00082792 0 0.00082802 3.3 0.00082794 3.3 0.0008280399999999999 0 0.0008279600000000001 0 0.00082806 3.3 0.0008279800000000001 3.3 0.00082808 0 0.0008280000000000001 0 0.0008281 3.3 0.0008280200000000001 3.3 0.00082812 0 0.00082804 0 0.00082814 3.3 0.00082806 3.3 0.00082816 0 0.00082808 0 0.00082818 3.3 0.0008281 3.3 0.0008282 0 0.00082812 0 0.00082822 3.3 0.00082814 3.3 0.0008282399999999999 0 0.00082816 0 0.0008282599999999999 3.3 0.0008281800000000001 3.3 0.00082828 0 0.0008282000000000001 0 0.0008283 3.3 0.0008282200000000001 3.3 0.00082832 0 0.00082824 0 0.00082834 3.3 0.00082826 3.3 0.00082836 0 0.00082828 0 0.00082838 3.3 0.0008283 3.3 0.0008284 0 0.00082832 0 0.00082842 3.3 0.00082834 3.3 0.00082844 0 0.00082836 0 0.0008284599999999999 3.3 0.0008283800000000001 3.3 0.00082848 0 0.0008284000000000001 0 0.0008285 3.3 0.0008284200000000001 3.3 0.00082852 0 0.0008284400000000001 0 0.00082854 3.3 0.00082846 3.3 0.00082856 0 0.00082848 0 0.00082858 3.3 0.0008285 3.3 0.0008286 0 0.00082852 0 0.00082862 3.3 0.00082854 3.3 0.00082864 0 0.00082856 0 0.0008286599999999999 3.3 0.00082858 3.3 0.0008286799999999999 0 0.0008286000000000001 0 0.0008287 3.3 0.0008286200000000001 3.3 0.00082872 0 0.0008286400000000001 0 0.00082874 3.3 0.00082866 3.3 0.00082876 0 0.00082868 0 0.00082878 3.3 0.0008287 3.3 0.0008288 0 0.00082872 0 0.00082882 3.3 0.00082874 3.3 0.00082884 0 0.00082876 0 0.00082886 3.3 0.00082878 3.3 0.0008288799999999999 0 0.0008288000000000001 0 0.0008289 3.3 0.0008288200000000001 3.3 0.00082892 0 0.0008288400000000001 0 0.00082894 3.3 0.0008288600000000001 3.3 0.00082896 0 0.00082888 0 0.00082898 3.3 0.0008289 3.3 0.000829 0 0.00082892 0 0.00082902 3.3 0.00082894 3.3 0.00082904 0 0.00082896 0 0.00082906 3.3 0.00082898 3.3 0.0008290799999999999 0 0.000829 0 0.0008290999999999999 3.3 0.0008290200000000001 3.3 0.00082912 0 0.0008290400000000001 0 0.00082914 3.3 0.0008290600000000001 3.3 0.00082916 0 0.00082908 0 0.00082918 3.3 0.0008291 3.3 0.0008292 0 0.00082912 0 0.00082922 3.3 0.00082914 3.3 0.00082924 0 0.00082916 0 0.00082926 3.3 0.00082918 3.3 0.00082928 0 0.0008292 0 0.0008292999999999999 3.3 0.0008292200000000001 3.3 0.00082932 0 0.0008292400000000001 0 0.00082934 3.3 0.0008292600000000001 3.3 0.00082936 0 0.0008292800000000001 0 0.00082938 3.3 0.0008293 3.3 0.0008294 0 0.00082932 0 0.00082942 3.3 0.00082934 3.3 0.00082944 0 0.00082936 0 0.00082946 3.3 0.00082938 3.3 0.00082948 0 0.0008294 0 0.0008294999999999999 3.3 0.00082942 3.3 0.0008295199999999999 0 0.0008294400000000001 0 0.00082954 3.3 0.0008294600000000001 3.3 0.00082956 0 0.0008294800000000001 0 0.00082958 3.3 0.0008295 3.3 0.0008296 0 0.00082952 0 0.00082962 3.3 0.00082954 3.3 0.00082964 0 0.00082956 0 0.00082966 3.3 0.00082958 3.3 0.00082968 0 0.0008296 0 0.0008297 3.3 0.00082962 3.3 0.0008297199999999999 0 0.0008296400000000001 0 0.00082974 3.3 0.0008296600000000001 3.3 0.00082976 0 0.0008296800000000001 0 0.00082978 3.3 0.0008297000000000001 3.3 0.0008298 0 0.00082972 0 0.00082982 3.3 0.00082974 3.3 0.00082984 0 0.00082976 0 0.00082986 3.3 0.00082978 3.3 0.00082988 0 0.0008298 0 0.0008299 3.3 0.00082982 3.3 0.0008299199999999999 0 0.00082984 0 0.0008299399999999999 3.3 0.0008298600000000001 3.3 0.00082996 0 0.0008298800000000001 0 0.00082998 3.3 0.0008299000000000001 3.3 0.00083 0 0.00082992 0 0.00083002 3.3 0.00082994 3.3 0.00083004 0 0.00082996 0 0.00083006 3.3 0.00082998 3.3 0.00083008 0 0.00083 0 0.0008301 3.3 0.00083002 3.3 0.00083012 0 0.00083004 0 0.0008301399999999999 3.3 0.0008300600000000001 3.3 0.00083016 0 0.0008300800000000001 0 0.00083018 3.3 0.0008301000000000001 3.3 0.0008302 0 0.0008301200000000001 0 0.00083022 3.3 0.00083014 3.3 0.00083024 0 0.00083016 0 0.00083026 3.3 0.00083018 3.3 0.00083028 0 0.0008302 0 0.0008303 3.3 0.00083022 3.3 0.00083032 0 0.00083024 0 0.0008303399999999999 3.3 0.00083026 3.3 0.0008303599999999999 0 0.0008302800000000001 0 0.00083038 3.3 0.0008303000000000001 3.3 0.0008304 0 0.0008303200000000001 0 0.00083042 3.3 0.00083034 3.3 0.00083044 0 0.00083036 0 0.00083046 3.3 0.00083038 3.3 0.00083048 0 0.0008304 0 0.0008305 3.3 0.00083042 3.3 0.00083052 0 0.00083044 0 0.00083054 3.3 0.00083046 3.3 0.0008305599999999999 0 0.0008304800000000001 0 0.00083058 3.3 0.0008305000000000001 3.3 0.0008306 0 0.0008305200000000001 0 0.00083062 3.3 0.0008305400000000001 3.3 0.00083064 0 0.00083056 0 0.00083066 3.3 0.00083058 3.3 0.00083068 0 0.0008306 0 0.0008307 3.3 0.00083062 3.3 0.00083072 0 0.00083064 0 0.00083074 3.3 0.00083066 3.3 0.0008307599999999999 0 0.00083068 0 0.0008307799999999999 3.3 0.0008307000000000001 3.3 0.0008308 0 0.0008307200000000001 0 0.00083082 3.3 0.0008307400000000001 3.3 0.00083084 0 0.00083076 0 0.00083086 3.3 0.00083078 3.3 0.00083088 0 0.0008308 0 0.0008309 3.3 0.00083082 3.3 0.00083092 0 0.00083084 0 0.00083094 3.3 0.00083086 3.3 0.0008309599999999999 0 0.00083088 0 0.0008309799999999999 3.3 0.0008309000000000001 3.3 0.000831 0 0.0008309200000000001 0 0.00083102 3.3 0.0008309400000000001 3.3 0.00083104 0 0.00083096 0 0.00083106 3.3 0.00083098 3.3 0.00083108 0 0.000831 0 0.0008311 3.3 0.00083102 3.3 0.00083112 0 0.00083104 0 0.00083114 3.3 0.00083106 3.3 0.00083116 0 0.00083108 0 0.0008311799999999999 3.3 0.0008311 3.3 0.0008311999999999999 0 0.0008311200000000001 0 0.00083122 3.3 0.0008311400000000001 3.3 0.00083124 0 0.0008311600000000001 0 0.00083126 3.3 0.00083118 3.3 0.00083128 0 0.0008312 0 0.0008313 3.3 0.00083122 3.3 0.00083132 0 0.00083124 0 0.00083134 3.3 0.00083126 3.3 0.00083136 0 0.00083128 0 0.0008313799999999999 3.3 0.0008313 3.3 0.0008313999999999999 0 0.0008313200000000001 0 0.00083142 3.3 0.0008313400000000001 3.3 0.00083144 0 0.0008313600000000001 0 0.00083146 3.3 0.00083138 3.3 0.00083148 0 0.0008314 0 0.0008315 3.3 0.00083142 3.3 0.00083152 0 0.00083144 0 0.00083154 3.3 0.00083146 3.3 0.00083156 0 0.00083148 0 0.00083158 3.3 0.0008315 3.3 0.0008315999999999999 0 0.0008315200000000001 0 0.00083162 3.3 0.0008315400000000001 3.3 0.00083164 0 0.0008315600000000001 0 0.00083166 3.3 0.0008315800000000001 3.3 0.00083168 0 0.0008316 0 0.0008317 3.3 0.00083162 3.3 0.00083172 0 0.00083164 0 0.00083174 3.3 0.00083166 3.3 0.00083176 0 0.00083168 0 0.00083178 3.3 0.0008317 3.3 0.0008317999999999999 0 0.00083172 0 0.0008318199999999999 3.3 0.0008317400000000001 3.3 0.00083184 0 0.0008317600000000001 0 0.00083186 3.3 0.0008317800000000001 3.3 0.00083188 0 0.0008318 0 0.0008319 3.3 0.00083182 3.3 0.00083192 0 0.00083184 0 0.00083194 3.3 0.00083186 3.3 0.00083196 0 0.00083188 0 0.00083198 3.3 0.0008319 3.3 0.000832 0 0.00083192 0 0.0008320199999999999 3.3 0.0008319400000000001 3.3 0.00083204 0 0.0008319600000000001 0 0.00083206 3.3 0.0008319800000000001 3.3 0.00083208 0 0.0008320000000000001 0 0.0008321 3.3 0.00083202 3.3 0.00083212 0 0.00083204 0 0.00083214 3.3 0.00083206 3.3 0.00083216 0 0.00083208 0 0.00083218 3.3 0.0008321 3.3 0.0008322 0 0.00083212 0 0.0008322199999999999 3.3 0.00083214 3.3 0.0008322399999999999 0 0.0008321600000000001 0 0.00083226 3.3 0.0008321800000000001 3.3 0.00083228 0 0.0008322000000000001 0 0.0008323 3.3 0.00083222 3.3 0.00083232 0 0.00083224 0 0.00083234 3.3 0.00083226 3.3 0.00083236 0 0.00083228 0 0.00083238 3.3 0.0008323 3.3 0.0008324 0 0.00083232 0 0.00083242 3.3 0.00083234 3.3 0.0008324399999999999 0 0.0008323600000000001 0 0.00083246 3.3 0.0008323800000000001 3.3 0.00083248 0 0.0008324000000000001 0 0.0008325 3.3 0.0008324200000000001 3.3 0.00083252 0 0.00083244 0 0.00083254 3.3 0.00083246 3.3 0.00083256 0 0.00083248 0 0.00083258 3.3 0.0008325 3.3 0.0008326 0 0.00083252 0 0.00083262 3.3 0.00083254 3.3 0.0008326399999999999 0 0.00083256 0 0.0008326599999999999 3.3 0.0008325800000000001 3.3 0.00083268 0 0.0008326000000000001 0 0.0008327 3.3 0.0008326200000000001 3.3 0.00083272 0 0.00083264 0 0.00083274 3.3 0.00083266 3.3 0.00083276 0 0.00083268 0 0.00083278 3.3 0.0008327 3.3 0.0008328 0 0.00083272 0 0.00083282 3.3 0.00083274 3.3 0.00083284 0 0.00083276 0 0.0008328599999999999 3.3 0.0008327800000000001 3.3 0.00083288 0 0.0008328000000000001 0 0.0008329 3.3 0.0008328200000000001 3.3 0.00083292 0 0.0008328400000000001 0 0.00083294 3.3 0.00083286 3.3 0.00083296 0 0.00083288 0 0.00083298 3.3 0.0008329 3.3 0.000833 0 0.00083292 0 0.00083302 3.3 0.00083294 3.3 0.00083304 0 0.00083296 0 0.0008330599999999999 3.3 0.00083298 3.3 0.0008330799999999999 0 0.0008330000000000001 0 0.0008331 3.3 0.0008330200000000001 3.3 0.00083312 0 0.0008330400000000001 0 0.00083314 3.3 0.00083306 3.3 0.00083316 0 0.00083308 0 0.00083318 3.3 0.0008331 3.3 0.0008332 0 0.00083312 0 0.00083322 3.3 0.00083314 3.3 0.00083324 0 0.00083316 0 0.00083326 3.3 0.00083318 3.3 0.0008332799999999999 0 0.0008332000000000001 0 0.0008333 3.3 0.0008332200000000001 3.3 0.00083332 0 0.0008332400000000001 0 0.00083334 3.3 0.0008332600000000001 3.3 0.00083336 0 0.00083328 0 0.00083338 3.3 0.0008333 3.3 0.0008334 0 0.00083332 0 0.00083342 3.3 0.00083334 3.3 0.00083344 0 0.00083336 0 0.00083346 3.3 0.00083338 3.3 0.0008334799999999999 0 0.0008334 0 0.0008334999999999999 3.3 0.0008334200000000001 3.3 0.00083352 0 0.0008334400000000001 0 0.00083354 3.3 0.0008334600000000001 3.3 0.00083356 0 0.00083348 0 0.00083358 3.3 0.0008335 3.3 0.0008336 0 0.00083352 0 0.00083362 3.3 0.00083354 3.3 0.00083364 0 0.00083356 0 0.00083366 3.3 0.00083358 3.3 0.00083368 0 0.0008336 0 0.0008336999999999999 3.3 0.0008336200000000001 3.3 0.00083372 0 0.0008336400000000001 0 0.00083374 3.3 0.0008336600000000001 3.3 0.00083376 0 0.0008336800000000001 0 0.00083378 3.3 0.0008337 3.3 0.0008338 0 0.00083372 0 0.00083382 3.3 0.00083374 3.3 0.00083384 0 0.00083376 0 0.00083386 3.3 0.00083378 3.3 0.00083388 0 0.0008338 0 0.0008338999999999999 3.3 0.00083382 3.3 0.0008339199999999999 0 0.0008338400000000001 0 0.00083394 3.3 0.0008338600000000001 3.3 0.00083396 0 0.0008338800000000001 0 0.00083398 3.3 0.0008339 3.3 0.000834 0 0.00083392 0 0.00083402 3.3 0.00083394 3.3 0.00083404 0 0.00083396 0 0.00083406 3.3 0.00083398 3.3 0.00083408 0 0.000834 0 0.0008340999999999999 3.3 0.00083402 3.3 0.0008341199999999999 0 0.0008340400000000001 0 0.00083414 3.3 0.0008340600000000001 3.3 0.00083416 0 0.0008340800000000001 0 0.00083418 3.3 0.0008341 3.3 0.0008342 0 0.00083412 0 0.00083422 3.3 0.00083414 3.3 0.00083424 0 0.00083416 0 0.00083426 3.3 0.00083418 3.3 0.00083428 0 0.0008342 0 0.0008343 3.3 0.00083422 3.3 0.0008343199999999999 0 0.00083424 0 0.0008343399999999999 3.3 0.0008342600000000001 3.3 0.00083436 0 0.0008342800000000001 0 0.00083438 3.3 0.0008343000000000001 3.3 0.0008344 0 0.00083432 0 0.00083442 3.3 0.00083434 3.3 0.00083444 0 0.00083436 0 0.00083446 3.3 0.00083438 3.3 0.00083448 0 0.0008344 0 0.0008345 3.3 0.00083442 3.3 0.0008345199999999999 0 0.00083444 0 0.0008345399999999999 3.3 0.0008344600000000001 3.3 0.00083456 0 0.0008344800000000001 0 0.00083458 3.3 0.0008345000000000001 3.3 0.0008346 0 0.00083452 0 0.00083462 3.3 0.00083454 3.3 0.00083464 0 0.00083456 0 0.00083466 3.3 0.00083458 3.3 0.00083468 0 0.0008346 0 0.0008347 3.3 0.00083462 3.3 0.00083472 0 0.00083464 0 0.0008347399999999999 3.3 0.00083466 3.3 0.0008347599999999999 0 0.0008346800000000001 0 0.00083478 3.3 0.0008347000000000001 3.3 0.0008348 0 0.0008347200000000001 0 0.00083482 3.3 0.00083474 3.3 0.00083484 0 0.00083476 0 0.00083486 3.3 0.00083478 3.3 0.00083488 0 0.0008348 0 0.0008349 3.3 0.00083482 3.3 0.00083492 0 0.00083484 0 0.0008349399999999999 3.3 0.00083486 3.3 0.0008349599999999999 0 0.0008348800000000001 0 0.00083498 3.3 0.0008349000000000001 3.3 0.000835 0 0.0008349200000000001 0 0.00083502 3.3 0.00083494 3.3 0.00083504 0 0.00083496 0 0.00083506 3.3 0.00083498 3.3 0.00083508 0 0.000835 0 0.0008351 3.3 0.00083502 3.3 0.00083512 0 0.00083504 0 0.00083514 3.3 0.00083506 3.3 0.0008351599999999999 0 0.0008350800000000001 0 0.00083518 3.3 0.0008351000000000001 3.3 0.0008352 0 0.0008351200000000001 0 0.00083522 3.3 0.0008351400000000001 3.3 0.00083524 0 0.00083516 0 0.00083526 3.3 0.00083518 3.3 0.00083528 0 0.0008352 0 0.0008353 3.3 0.00083522 3.3 0.00083532 0 0.00083524 0 0.00083534 3.3 0.00083526 3.3 0.0008353599999999999 0 0.00083528 0 0.0008353799999999999 3.3 0.0008353000000000001 3.3 0.0008354 0 0.0008353200000000001 0 0.00083542 3.3 0.0008353400000000001 3.3 0.00083544 0 0.00083536 0 0.00083546 3.3 0.00083538 3.3 0.00083548 0 0.0008354 0 0.0008355 3.3 0.00083542 3.3 0.00083552 0 0.00083544 0 0.00083554 3.3 0.00083546 3.3 0.00083556 0 0.00083548 0 0.0008355799999999999 3.3 0.0008355000000000001 3.3 0.0008356 0 0.0008355200000000001 0 0.00083562 3.3 0.0008355400000000001 3.3 0.00083564 0 0.0008355600000000001 0 0.00083566 3.3 0.00083558 3.3 0.00083568 0 0.0008356 0 0.0008357 3.3 0.00083562 3.3 0.00083572 0 0.00083564 0 0.00083574 3.3 0.00083566 3.3 0.00083576 0 0.00083568 0 0.0008357799999999999 3.3 0.0008357 3.3 0.0008357999999999999 0 0.0008357200000000001 0 0.00083582 3.3 0.0008357400000000001 3.3 0.00083584 0 0.0008357600000000001 0 0.00083586 3.3 0.00083578 3.3 0.00083588 0 0.0008358 0 0.0008359 3.3 0.00083582 3.3 0.00083592 0 0.00083584 0 0.00083594 3.3 0.00083586 3.3 0.00083596 0 0.00083588 0 0.00083598 3.3 0.0008359 3.3 0.0008359999999999999 0 0.0008359200000000001 0 0.00083602 3.3 0.0008359400000000001 3.3 0.00083604 0 0.0008359600000000001 0 0.00083606 3.3 0.0008359800000000001 3.3 0.00083608 0 0.000836 0 0.0008361 3.3 0.00083602 3.3 0.00083612 0 0.00083604 0 0.00083614 3.3 0.00083606 3.3 0.00083616 0 0.00083608 0 0.00083618 3.3 0.0008361 3.3 0.0008361999999999999 0 0.00083612 0 0.0008362199999999999 3.3 0.0008361400000000001 3.3 0.00083624 0 0.0008361600000000001 0 0.00083626 3.3 0.0008361800000000001 3.3 0.00083628 0 0.0008362 0 0.0008363 3.3 0.00083622 3.3 0.00083632 0 0.00083624 0 0.00083634 3.3 0.00083626 3.3 0.00083636 0 0.00083628 0 0.00083638 3.3 0.0008363 3.3 0.0008364 0 0.00083632 0 0.0008364199999999999 3.3 0.0008363400000000001 3.3 0.00083644 0 0.0008363600000000001 0 0.00083646 3.3 0.0008363800000000001 3.3 0.00083648 0 0.0008364000000000001 0 0.0008365 3.3 0.00083642 3.3 0.00083652 0 0.00083644 0 0.00083654 3.3 0.00083646 3.3 0.00083656 0 0.00083648 0 0.00083658 3.3 0.0008365 3.3 0.0008366 0 0.00083652 0 0.0008366199999999999 3.3 0.00083654 3.3 0.0008366399999999999 0 0.0008365600000000001 0 0.00083666 3.3 0.0008365800000000001 3.3 0.00083668 0 0.0008366000000000001 0 0.0008367 3.3 0.00083662 3.3 0.00083672 0 0.00083664 0 0.00083674 3.3 0.00083666 3.3 0.00083676 0 0.00083668 0 0.00083678 3.3 0.0008367 3.3 0.0008368 0 0.00083672 0 0.00083682 3.3 0.00083674 3.3 0.0008368399999999999 0 0.0008367600000000001 0 0.00083686 3.3 0.0008367800000000001 3.3 0.00083688 0 0.0008368000000000001 0 0.0008369 3.3 0.0008368200000000001 3.3 0.00083692 0 0.00083684 0 0.00083694 3.3 0.00083686 3.3 0.00083696 0 0.00083688 0 0.00083698 3.3 0.0008369 3.3 0.000837 0 0.00083692 0 0.00083702 3.3 0.00083694 3.3 0.0008370399999999999 0 0.00083696 0 0.0008370599999999999 3.3 0.0008369800000000001 3.3 0.00083708 0 0.0008370000000000001 0 0.0008371 3.3 0.0008370200000000001 3.3 0.00083712 0 0.00083704 0 0.00083714 3.3 0.00083706 3.3 0.00083716 0 0.00083708 0 0.00083718 3.3 0.0008371 3.3 0.0008372 0 0.00083712 0 0.00083722 3.3 0.00083714 3.3 0.00083724 0 0.00083716 0 0.0008372599999999999 3.3 0.0008371800000000001 3.3 0.00083728 0 0.0008372000000000001 0 0.0008373 3.3 0.0008372200000000001 3.3 0.00083732 0 0.0008372400000000001 0 0.00083734 3.3 0.00083726 3.3 0.00083736 0 0.00083728 0 0.00083738 3.3 0.0008373 3.3 0.0008374 0 0.00083732 0 0.00083742 3.3 0.00083734 3.3 0.00083744 0 0.00083736 0 0.0008374599999999999 3.3 0.00083738 3.3 0.0008374799999999999 0 0.0008374000000000001 0 0.0008375 3.3 0.0008374200000000001 3.3 0.00083752 0 0.0008374400000000001 0 0.00083754 3.3 0.00083746 3.3 0.00083756 0 0.00083748 0 0.00083758 3.3 0.0008375 3.3 0.0008376 0 0.00083752 0 0.00083762 3.3 0.00083754 3.3 0.00083764 0 0.00083756 0 0.0008376599999999999 3.3 0.00083758 3.3 0.0008376799999999999 0 0.0008376000000000001 0 0.0008377 3.3 0.0008376200000000001 3.3 0.00083772 0 0.0008376400000000001 0 0.00083774 3.3 0.00083766 3.3 0.00083776 0 0.00083768 0 0.00083778 3.3 0.0008377 3.3 0.0008378 0 0.00083772 0 0.00083782 3.3 0.00083774 3.3 0.00083784 0 0.00083776 0 0.00083786 3.3 0.00083778 3.3 0.0008378799999999999 0 0.0008378 0 0.0008378999999999999 3.3 0.0008378200000000001 3.3 0.00083792 0 0.0008378400000000001 0 0.00083794 3.3 0.0008378600000000001 3.3 0.00083796 0 0.00083788 0 0.00083798 3.3 0.0008379 3.3 0.000838 0 0.00083792 0 0.00083802 3.3 0.00083794 3.3 0.00083804 0 0.00083796 0 0.00083806 3.3 0.00083798 3.3 0.0008380799999999999 0 0.000838 0 0.0008380999999999999 3.3 0.0008380200000000001 3.3 0.00083812 0 0.0008380400000000001 0 0.00083814 3.3 0.0008380600000000001 3.3 0.00083816 0 0.00083808 0 0.00083818 3.3 0.0008381 3.3 0.0008382 0 0.00083812 0 0.00083822 3.3 0.00083814 3.3 0.00083824 0 0.00083816 0 0.00083826 3.3 0.00083818 3.3 0.00083828 0 0.0008382 0 0.0008382999999999999 3.3 0.00083822 3.3 0.0008383199999999999 0 0.0008382400000000001 0 0.00083834 3.3 0.0008382600000000001 3.3 0.00083836 0 0.0008382800000000001 0 0.00083838 3.3 0.0008383 3.3 0.0008384 0 0.00083832 0 0.00083842 3.3 0.00083834 3.3 0.00083844 0 0.00083836 0 0.00083846 3.3 0.00083838 3.3 0.00083848 0 0.0008384 0 0.0008384999999999999 3.3 0.00083842 3.3 0.0008385199999999999 0 0.0008384400000000001 0 0.00083854 3.3 0.0008384600000000001 3.3 0.00083856 0 0.0008384800000000001 0 0.00083858 3.3 0.0008385 3.3 0.0008386 0 0.00083852 0 0.00083862 3.3 0.00083854 3.3 0.00083864 0 0.00083856 0 0.00083866 3.3 0.00083858 3.3 0.00083868 0 0.0008386 0 0.0008387 3.3 0.00083862 3.3 0.0008387199999999999 0 0.0008386400000000001 0 0.00083874 3.3 0.0008386600000000001 3.3 0.00083876 0 0.0008386800000000001 0 0.00083878 3.3 0.0008387000000000001 3.3 0.0008388 0 0.00083872 0 0.00083882 3.3 0.00083874 3.3 0.00083884 0 0.00083876 0 0.00083886 3.3 0.00083878 3.3 0.00083888 0 0.0008388 0 0.0008389 3.3 0.00083882 3.3 0.0008389199999999999 0 0.00083884 0 0.0008389399999999999 3.3 0.0008388600000000001 3.3 0.00083896 0 0.0008388800000000001 0 0.00083898 3.3 0.0008389000000000001 3.3 0.000839 0 0.00083892 0 0.00083902 3.3 0.00083894 3.3 0.00083904 0 0.00083896 0 0.00083906 3.3 0.00083898 3.3 0.00083908 0 0.000839 0 0.0008391 3.3 0.00083902 3.3 0.00083912 0 0.00083904 0 0.0008391399999999999 3.3 0.0008390600000000001 3.3 0.00083916 0 0.0008390800000000001 0 0.00083918 3.3 0.0008391000000000001 3.3 0.0008392 0 0.0008391200000000001 0 0.00083922 3.3 0.00083914 3.3 0.00083924 0 0.00083916 0 0.00083926 3.3 0.00083918 3.3 0.00083928 0 0.0008392 0 0.0008393 3.3 0.00083922 3.3 0.00083932 0 0.00083924 0 0.0008393399999999999 3.3 0.00083926 3.3 0.0008393599999999999 0 0.0008392800000000001 0 0.00083938 3.3 0.0008393000000000001 3.3 0.0008394 0 0.0008393200000000001 0 0.00083942 3.3 0.00083934 3.3 0.00083944 0 0.00083936 0 0.00083946 3.3 0.00083938 3.3 0.00083948 0 0.0008394 0 0.0008395 3.3 0.00083942 3.3 0.00083952 0 0.00083944 0 0.00083954 3.3 0.00083946 3.3 0.0008395599999999999 0 0.0008394800000000001 0 0.00083958 3.3 0.0008395000000000001 3.3 0.0008396 0 0.0008395200000000001 0 0.00083962 3.3 0.0008395400000000001 3.3 0.00083964 0 0.00083956 0 0.00083966 3.3 0.00083958 3.3 0.00083968 0 0.0008396 0 0.0008397 3.3 0.00083962 3.3 0.00083972 0 0.00083964 0 0.00083974 3.3 0.00083966 3.3 0.0008397599999999999 0 0.00083968 0 0.0008397799999999999 3.3 0.0008397000000000001 3.3 0.0008398 0 0.0008397200000000001 0 0.00083982 3.3 0.0008397400000000001 3.3 0.00083984 0 0.00083976 0 0.00083986 3.3 0.00083978 3.3 0.00083988 0 0.0008398 0 0.0008399 3.3 0.00083982 3.3 0.00083992 0 0.00083984 0 0.00083994 3.3 0.00083986 3.3 0.00083996 0 0.00083988 0 0.0008399799999999999 3.3 0.0008399000000000001 3.3 0.00084 0 0.0008399200000000001 0 0.00084002 3.3 0.0008399400000000001 3.3 0.00084004 0 0.0008399600000000001 0 0.00084006 3.3 0.00083998 3.3 0.00084008 0 0.00084 0 0.0008401 3.3 0.00084002 3.3 0.00084012 0 0.00084004 0 0.00084014 3.3 0.00084006 3.3 0.00084016 0 0.00084008 0 0.0008401799999999999 3.3 0.0008401 3.3 0.0008401999999999999 0 0.0008401200000000001 0 0.00084022 3.3 0.0008401400000000001 3.3 0.00084024 0 0.0008401600000000001 0 0.00084026 3.3 0.00084018 3.3 0.00084028 0 0.0008402 0 0.0008403 3.3 0.00084022 3.3 0.00084032 0 0.00084024 0 0.00084034 3.3 0.00084026 3.3 0.00084036 0 0.00084028 0 0.00084038 3.3 0.0008403 3.3 0.0008403999999999999 0 0.0008403200000000001 0 0.00084042 3.3 0.0008403400000000001 3.3 0.00084044 0 0.0008403600000000001 0 0.00084046 3.3 0.0008403800000000001 3.3 0.00084048 0 0.0008404 0 0.0008405 3.3 0.00084042 3.3 0.00084052 0 0.00084044 0 0.00084054 3.3 0.00084046 3.3 0.00084056 0 0.00084048 0 0.00084058 3.3 0.0008405 3.3 0.0008405999999999999 0 0.00084052 0 0.0008406199999999999 3.3 0.0008405400000000001 3.3 0.00084064 0 0.0008405600000000001 0 0.00084066 3.3 0.0008405800000000001 3.3 0.00084068 0 0.0008406 0 0.0008407 3.3 0.00084062 3.3 0.00084072 0 0.00084064 0 0.00084074 3.3 0.00084066 3.3 0.00084076 0 0.00084068 0 0.00084078 3.3 0.0008407 3.3 0.0008408 0 0.00084072 0 0.0008408199999999999 3.3 0.0008407400000000001 3.3 0.00084084 0 0.0008407600000000001 0 0.00084086 3.3 0.0008407800000000001 3.3 0.00084088 0 0.0008408000000000001 0 0.0008409 3.3 0.00084082 3.3 0.00084092 0 0.00084084 0 0.00084094 3.3 0.00084086 3.3 0.00084096 0 0.00084088 0 0.00084098 3.3 0.0008409 3.3 0.000841 0 0.00084092 0 0.0008410199999999999 3.3 0.00084094 3.3 0.0008410399999999999 0 0.0008409600000000001 0 0.00084106 3.3 0.0008409800000000001 3.3 0.00084108 0 0.0008410000000000001 0 0.0008411 3.3 0.00084102 3.3 0.00084112 0 0.00084104 0 0.00084114 3.3 0.00084106 3.3 0.00084116 0 0.00084108 0 0.00084118 3.3 0.0008411 3.3 0.0008412 0 0.00084112 0 0.0008412199999999999 3.3 0.00084114 3.3 0.0008412399999999999 0 0.0008411600000000001 0 0.00084126 3.3 0.0008411800000000001 3.3 0.00084128 0 0.0008412000000000001 0 0.0008413 3.3 0.00084122 3.3 0.00084132 0 0.00084124 0 0.00084134 3.3 0.00084126 3.3 0.00084136 0 0.00084128 0 0.00084138 3.3 0.0008413 3.3 0.0008414 0 0.00084132 0 0.00084142 3.3 0.00084134 3.3 0.0008414399999999999 0 0.00084136 0 0.0008414599999999999 3.3 0.0008413800000000001 3.3 0.00084148 0 0.0008414000000000001 0 0.0008415 3.3 0.0008414200000000001 3.3 0.00084152 0 0.00084144 0 0.00084154 3.3 0.00084146 3.3 0.00084156 0 0.00084148 0 0.00084158 3.3 0.0008415 3.3 0.0008416 0 0.00084152 0 0.00084162 3.3 0.00084154 3.3 0.0008416399999999999 0 0.00084156 0 0.0008416599999999999 3.3 0.0008415800000000001 3.3 0.00084168 0 0.0008416000000000001 0 0.0008417 3.3 0.0008416200000000001 3.3 0.00084172 0 0.00084164 0 0.00084174 3.3 0.00084166 3.3 0.00084176 0 0.00084168 0 0.00084178 3.3 0.0008417 3.3 0.0008418 0 0.00084172 0 0.00084182 3.3 0.00084174 3.3 0.00084184 0 0.00084176 0 0.0008418599999999999 3.3 0.0008417800000000001 3.3 0.00084188 0 0.0008418000000000001 0 0.0008419 3.3 0.0008418200000000001 3.3 0.00084192 0 0.0008418400000000001 0 0.00084194 3.3 0.00084186 3.3 0.00084196 0 0.00084188 0 0.00084198 3.3 0.0008419 3.3 0.000842 0 0.00084192 0 0.00084202 3.3 0.00084194 3.3 0.00084204 0 0.00084196 0 0.0008420599999999999 3.3 0.00084198 3.3 0.0008420799999999999 0 0.0008420000000000001 0 0.0008421 3.3 0.0008420200000000001 3.3 0.00084212 0 0.0008420400000000001 0 0.00084214 3.3 0.00084206 3.3 0.00084216 0 0.00084208 0 0.00084218 3.3 0.0008421 3.3 0.0008422 0 0.00084212 0 0.00084222 3.3 0.00084214 3.3 0.00084224 0 0.00084216 0 0.00084226 3.3 0.00084218 3.3 0.0008422799999999999 0 0.0008422000000000001 0 0.0008423 3.3 0.0008422200000000001 3.3 0.00084232 0 0.0008422400000000001 0 0.00084234 3.3 0.0008422600000000001 3.3 0.00084236 0 0.00084228 0 0.00084238 3.3 0.0008423 3.3 0.0008424 0 0.00084232 0 0.00084242 3.3 0.00084234 3.3 0.00084244 0 0.00084236 0 0.00084246 3.3 0.00084238 3.3 0.0008424799999999999 0 0.0008424 0 0.0008424999999999999 3.3 0.0008424200000000001 3.3 0.00084252 0 0.0008424400000000001 0 0.00084254 3.3 0.0008424600000000001 3.3 0.00084256 0 0.00084248 0 0.00084258 3.3 0.0008425 3.3 0.0008426 0 0.00084252 0 0.00084262 3.3 0.00084254 3.3 0.00084264 0 0.00084256 0 0.00084266 3.3 0.00084258 3.3 0.00084268 0 0.0008426 0 0.0008426999999999999 3.3 0.0008426200000000001 3.3 0.00084272 0 0.0008426400000000001 0 0.00084274 3.3 0.0008426600000000001 3.3 0.00084276 0 0.0008426800000000001 0 0.00084278 3.3 0.0008427 3.3 0.0008428 0 0.00084272 0 0.00084282 3.3 0.00084274 3.3 0.00084284 0 0.00084276 0 0.00084286 3.3 0.00084278 3.3 0.00084288 0 0.0008428 0 0.0008428999999999999 3.3 0.00084282 3.3 0.0008429199999999999 0 0.0008428400000000001 0 0.00084294 3.3 0.0008428600000000001 3.3 0.00084296 0 0.0008428800000000001 0 0.00084298 3.3 0.0008429 3.3 0.000843 0 0.00084292 0 0.00084302 3.3 0.00084294 3.3 0.00084304 0 0.00084296 0 0.00084306 3.3 0.00084298 3.3 0.00084308 0 0.000843 0 0.0008431 3.3 0.00084302 3.3 0.0008431199999999999 0 0.0008430400000000001 0 0.00084314 3.3 0.0008430600000000001 3.3 0.00084316 0 0.0008430800000000001 0 0.00084318 3.3 0.0008431000000000001 3.3 0.0008432 0 0.00084312 0 0.00084322 3.3 0.00084314 3.3 0.00084324 0 0.00084316 0 0.00084326 3.3 0.00084318 3.3 0.00084328 0 0.0008432 0 0.0008433 3.3 0.00084322 3.3 0.0008433199999999999 0 0.00084324 0 0.0008433399999999999 3.3 0.0008432600000000001 3.3 0.00084336 0 0.0008432800000000001 0 0.00084338 3.3 0.0008433000000000001 3.3 0.0008434 0 0.00084332 0 0.00084342 3.3 0.00084334 3.3 0.00084344 0 0.00084336 0 0.00084346 3.3 0.00084338 3.3 0.00084348 0 0.0008434 0 0.0008435 3.3 0.00084342 3.3 0.00084352 0 0.00084344 0 0.0008435399999999999 3.3 0.0008434600000000001 3.3 0.00084356 0 0.0008434800000000001 0 0.00084358 3.3 0.0008435000000000001 3.3 0.0008436 0 0.0008435200000000001 0 0.00084362 3.3 0.00084354 3.3 0.00084364 0 0.00084356 0 0.00084366 3.3 0.00084358 3.3 0.00084368 0 0.0008436 0 0.0008437 3.3 0.00084362 3.3 0.00084372 0 0.00084364 0 0.0008437399999999999 3.3 0.00084366 3.3 0.0008437599999999999 0 0.0008436800000000001 0 0.00084378 3.3 0.0008437000000000001 3.3 0.0008438 0 0.0008437200000000001 0 0.00084382 3.3 0.00084374 3.3 0.00084384 0 0.00084376 0 0.00084386 3.3 0.00084378 3.3 0.00084388 0 0.0008438 0 0.0008439 3.3 0.00084382 3.3 0.00084392 0 0.00084384 0 0.00084394 3.3 0.00084386 3.3 0.0008439599999999999 0 0.0008438800000000001 0 0.00084398 3.3 0.0008439000000000001 3.3 0.000844 0 0.0008439200000000001 0 0.00084402 3.3 0.0008439400000000001 3.3 0.00084404 0 0.00084396 0 0.00084406 3.3 0.00084398 3.3 0.00084408 0 0.000844 0 0.0008441 3.3 0.00084402 3.3 0.00084412 0 0.00084404 0 0.00084414 3.3 0.00084406 3.3 0.0008441599999999999 0 0.00084408 0 0.0008441799999999999 3.3 0.0008441000000000001 3.3 0.0008442 0 0.0008441200000000001 0 0.00084422 3.3 0.0008441400000000001 3.3 0.00084424 0 0.00084416 0 0.00084426 3.3 0.00084418 3.3 0.00084428 0 0.0008442 0 0.0008443 3.3 0.00084422 3.3 0.00084432 0 0.00084424 0 0.00084434 3.3 0.00084426 3.3 0.0008443599999999999 0 0.00084428 0 0.0008443799999999999 3.3 0.0008443000000000001 3.3 0.0008444 0 0.0008443200000000001 0 0.00084442 3.3 0.0008443400000000001 3.3 0.00084444 0 0.00084436 0 0.00084446 3.3 0.00084438 3.3 0.00084448 0 0.0008444 0 0.0008445 3.3 0.00084442 3.3 0.00084452 0 0.00084444 0 0.00084454 3.3 0.00084446 3.3 0.00084456 0 0.00084448 0 0.0008445799999999999 3.3 0.0008445 3.3 0.0008445999999999999 0 0.0008445200000000001 0 0.00084462 3.3 0.0008445400000000001 3.3 0.00084464 0 0.0008445600000000001 0 0.00084466 3.3 0.00084458 3.3 0.00084468 0 0.0008446 0 0.0008447 3.3 0.00084462 3.3 0.00084472 0 0.00084464 0 0.00084474 3.3 0.00084466 3.3 0.00084476 0 0.00084468 0 0.0008447799999999999 3.3 0.0008447 3.3 0.0008447999999999999 0 0.0008447200000000001 0 0.00084482 3.3 0.0008447400000000001 3.3 0.00084484 0 0.0008447600000000001 0 0.00084486 3.3 0.00084478 3.3 0.00084488 0 0.0008448 0 0.0008449 3.3 0.00084482 3.3 0.00084492 0 0.00084484 0 0.00084494 3.3 0.00084486 3.3 0.00084496 0 0.00084488 0 0.00084498 3.3 0.0008449 3.3 0.0008449999999999999 0 0.00084492 0 0.0008450199999999999 3.3 0.0008449400000000001 3.3 0.00084504 0 0.0008449600000000001 0 0.00084506 3.3 0.0008449800000000001 3.3 0.00084508 0 0.000845 0 0.0008451 3.3 0.00084502 3.3 0.00084512 0 0.00084504 0 0.00084514 3.3 0.00084506 3.3 0.00084516 0 0.00084508 0 0.00084518 3.3 0.0008451 3.3 0.0008451999999999999 0 0.00084512 0 0.0008452199999999999 3.3 0.0008451400000000001 3.3 0.00084524 0 0.0008451600000000001 0 0.00084526 3.3 0.0008451800000000001 3.3 0.00084528 0 0.0008452 0 0.0008453 3.3 0.00084522 3.3 0.00084532 0 0.00084524 0 0.00084534 3.3 0.00084526 3.3 0.00084536 0 0.00084528 0 0.00084538 3.3 0.0008453 3.3 0.0008454 0 0.00084532 0 0.0008454199999999999 3.3 0.0008453400000000001 3.3 0.00084544 0 0.0008453600000000001 0 0.00084546 3.3 0.0008453800000000001 3.3 0.00084548 0 0.0008454000000000001 0 0.0008455 3.3 0.00084542 3.3 0.00084552 0 0.00084544 0 0.00084554 3.3 0.00084546 3.3 0.00084556 0 0.00084548 0 0.00084558 3.3 0.0008455 3.3 0.0008456 0 0.00084552 0 0.0008456199999999999 3.3 0.00084554 3.3 0.0008456399999999999 0 0.0008455600000000001 0 0.00084566 3.3 0.0008455800000000001 3.3 0.00084568 0 0.0008456000000000001 0 0.0008457 3.3 0.00084562 3.3 0.00084572 0 0.00084564 0 0.00084574 3.3 0.00084566 3.3 0.00084576 0 0.00084568 0 0.00084578 3.3 0.0008457 3.3 0.0008458 0 0.00084572 0 0.00084582 3.3 0.00084574 3.3 0.0008458399999999999 0 0.0008457600000000001 0 0.00084586 3.3 0.0008457800000000001 3.3 0.00084588 0 0.0008458000000000001 0 0.0008459 3.3 0.0008458200000000001 3.3 0.00084592 0 0.00084584 0 0.00084594 3.3 0.00084586 3.3 0.00084596 0 0.00084588 0 0.00084598 3.3 0.0008459 3.3 0.000846 0 0.00084592 0 0.00084602 3.3 0.00084594 3.3 0.0008460399999999999 0 0.00084596 0 0.0008460599999999999 3.3 0.0008459800000000001 3.3 0.00084608 0 0.0008460000000000001 0 0.0008461 3.3 0.0008460200000000001 3.3 0.00084612 0 0.00084604 0 0.00084614 3.3 0.00084606 3.3 0.00084616 0 0.00084608 0 0.00084618 3.3 0.0008461 3.3 0.0008462 0 0.00084612 0 0.00084622 3.3 0.00084614 3.3 0.00084624 0 0.00084616 0 0.0008462599999999999 3.3 0.0008461800000000001 3.3 0.00084628 0 0.0008462000000000001 0 0.0008463 3.3 0.0008462200000000001 3.3 0.00084632 0 0.0008462400000000001 0 0.00084634 3.3 0.00084626 3.3 0.00084636 0 0.00084628 0 0.00084638 3.3 0.0008463 3.3 0.0008464 0 0.00084632 0 0.00084642 3.3 0.00084634 3.3 0.00084644 0 0.00084636 0 0.0008464599999999999 3.3 0.00084638 3.3 0.0008464799999999999 0 0.0008464000000000001 0 0.0008465 3.3 0.0008464200000000001 3.3 0.00084652 0 0.0008464400000000001 0 0.00084654 3.3 0.00084646 3.3 0.00084656 0 0.00084648 0 0.00084658 3.3 0.0008465 3.3 0.0008466 0 0.00084652 0 0.00084662 3.3 0.00084654 3.3 0.00084664 0 0.00084656 0 0.00084666 3.3 0.00084658 3.3 0.0008466799999999999 0 0.0008466000000000001 0 0.0008467 3.3 0.0008466200000000001 3.3 0.00084672 0 0.0008466400000000001 0 0.00084674 3.3 0.0008466600000000001 3.3 0.00084676 0 0.00084668 0 0.00084678 3.3 0.0008467 3.3 0.0008468 0 0.00084672 0 0.00084682 3.3 0.00084674 3.3 0.00084684 0 0.00084676 0 0.00084686 3.3 0.00084678 3.3 0.0008468799999999999 0 0.0008468 0 0.0008468999999999999 3.3 0.0008468200000000001 3.3 0.00084692 0 0.0008468400000000001 0 0.00084694 3.3 0.0008468600000000001 3.3 0.00084696 0 0.00084688 0 0.00084698 3.3 0.0008469 3.3 0.000847 0 0.00084692 0 0.00084702 3.3 0.00084694 3.3 0.00084704 0 0.00084696 0 0.00084706 3.3 0.00084698 3.3 0.00084708 0 0.000847 0 0.0008470999999999999 3.3 0.0008470200000000001 3.3 0.00084712 0 0.0008470400000000001 0 0.00084714 3.3 0.0008470600000000001 3.3 0.00084716 0 0.0008470800000000001 0 0.00084718 3.3 0.0008471 3.3 0.0008472 0 0.00084712 0 0.00084722 3.3 0.00084714 3.3 0.00084724 0 0.00084716 0 0.00084726 3.3 0.00084718 3.3 0.00084728 0 0.0008472 0 0.0008472999999999999 3.3 0.00084722 3.3 0.0008473199999999999 0 0.0008472400000000001 0 0.00084734 3.3 0.0008472600000000001 3.3 0.00084736 0 0.0008472800000000001 0 0.00084738 3.3 0.0008473 3.3 0.0008474 0 0.00084732 0 0.00084742 3.3 0.00084734 3.3 0.00084744 0 0.00084736 0 0.00084746 3.3 0.00084738 3.3 0.00084748 0 0.0008474 0 0.0008475 3.3 0.00084742 3.3 0.0008475199999999999 0 0.0008474400000000001 0 0.00084754 3.3 0.0008474600000000001 3.3 0.00084756 0 0.0008474800000000001 0 0.00084758 3.3 0.0008475000000000001 3.3 0.0008476 0 0.00084752 0 0.00084762 3.3 0.00084754 3.3 0.00084764 0 0.00084756 0 0.00084766 3.3 0.00084758 3.3 0.00084768 0 0.0008476 0 0.0008477 3.3 0.00084762 3.3 0.0008477199999999999 0 0.00084764 0 0.0008477399999999999 3.3 0.0008476600000000001 3.3 0.00084776 0 0.0008476800000000001 0 0.00084778 3.3 0.0008477000000000001 3.3 0.0008478 0 0.00084772 0 0.00084782 3.3 0.00084774 3.3 0.00084784 0 0.00084776 0 0.00084786 3.3 0.00084778 3.3 0.00084788 0 0.0008478 0 0.0008479 3.3 0.00084782 3.3 0.0008479199999999999 0 0.00084784 0 0.0008479399999999999 3.3 0.0008478600000000001 3.3 0.00084796 0 0.0008478800000000001 0 0.00084798 3.3 0.0008479000000000001 3.3 0.000848 0 0.00084792 0 0.00084802 3.3 0.00084794 3.3 0.00084804 0 0.00084796 0 0.00084806 3.3 0.00084798 3.3 0.00084808 0 0.000848 0 0.0008481 3.3 0.00084802 3.3 0.00084812 0 0.00084804 0 0.0008481399999999999 3.3 0.00084806 3.3 0.0008481599999999999 0 0.0008480800000000001 0 0.00084818 3.3 0.0008481000000000001 3.3 0.0008482 0 0.0008481200000000001 0 0.00084822 3.3 0.00084814 3.3 0.00084824 0 0.00084816 0 0.00084826 3.3 0.00084818 3.3 0.00084828 0 0.0008482 0 0.0008483 3.3 0.00084822 3.3 0.00084832 0 0.00084824 0 0.0008483399999999999 3.3 0.00084826 3.3 0.0008483599999999999 0 0.0008482800000000001 0 0.00084838 3.3 0.0008483000000000001 3.3 0.0008484 0 0.0008483200000000001 0 0.00084842 3.3 0.00084834 3.3 0.00084844 0 0.00084836 0 0.00084846 3.3 0.00084838 3.3 0.00084848 0 0.0008484 0 0.0008485 3.3 0.00084842 3.3 0.00084852 0 0.00084844 0 0.00084854 3.3 0.00084846 3.3 0.0008485599999999999 0 0.00084848 0 0.0008485799999999999 3.3 0.0008485000000000001 3.3 0.0008486 0 0.0008485200000000001 0 0.00084862 3.3 0.0008485400000000001 3.3 0.00084864 0 0.00084856 0 0.00084866 3.3 0.00084858 3.3 0.00084868 0 0.0008486 0 0.0008487 3.3 0.00084862 3.3 0.00084872 0 0.00084864 0 0.00084874 3.3 0.00084866 3.3 0.0008487599999999999 0 0.00084868 0 0.0008487799999999999 3.3 0.0008487000000000001 3.3 0.0008488 0 0.0008487200000000001 0 0.00084882 3.3 0.0008487400000000001 3.3 0.00084884 0 0.00084876 0 0.00084886 3.3 0.00084878 3.3 0.00084888 0 0.0008488 0 0.0008489 3.3 0.00084882 3.3 0.00084892 0 0.00084884 0 0.00084894 3.3 0.00084886 3.3 0.00084896 0 0.00084888 0 0.0008489799999999999 3.3 0.0008489000000000001 3.3 0.000849 0 0.0008489200000000001 0 0.00084902 3.3 0.0008489400000000001 3.3 0.00084904 0 0.0008489600000000001 0 0.00084906 3.3 0.00084898 3.3 0.00084908 0 0.000849 0 0.0008491 3.3 0.00084902 3.3 0.00084912 0 0.00084904 0 0.00084914 3.3 0.00084906 3.3 0.00084916 0 0.00084908 0 0.0008491799999999999 3.3 0.0008491 3.3 0.0008491999999999999 0 0.0008491200000000001 0 0.00084922 3.3 0.0008491400000000001 3.3 0.00084924 0 0.0008491600000000001 0 0.00084926 3.3 0.00084918 3.3 0.00084928 0 0.0008492 0 0.0008493 3.3 0.00084922 3.3 0.00084932 0 0.00084924 0 0.00084934 3.3 0.00084926 3.3 0.00084936 0 0.00084928 0 0.00084938 3.3 0.0008493 3.3 0.0008493999999999999 0 0.0008493200000000001 0 0.00084942 3.3 0.0008493400000000001 3.3 0.00084944 0 0.0008493600000000001 0 0.00084946 3.3 0.0008493800000000001 3.3 0.00084948 0 0.0008494 0 0.0008495 3.3 0.00084942 3.3 0.00084952 0 0.00084944 0 0.00084954 3.3 0.00084946 3.3 0.00084956 0 0.00084948 0 0.00084958 3.3 0.0008495 3.3 0.0008495999999999999 0 0.00084952 0 0.0008496199999999999 3.3 0.0008495400000000001 3.3 0.00084964 0 0.0008495600000000001 0 0.00084966 3.3 0.0008495800000000001 3.3 0.00084968 0 0.0008496 0 0.0008497 3.3 0.00084962 3.3 0.00084972 0 0.00084964 0 0.00084974 3.3 0.00084966 3.3 0.00084976 0 0.00084968 0 0.00084978 3.3 0.0008497 3.3 0.0008498 0 0.00084972 0 0.0008498199999999999 3.3 0.0008497400000000001 3.3 0.00084984 0 0.0008497600000000001 0 0.00084986 3.3 0.0008497800000000001 3.3 0.00084988 0 0.0008498000000000001 0 0.0008499 3.3 0.00084982 3.3 0.00084992 0 0.00084984 0 0.00084994 3.3 0.00084986 3.3 0.00084996 0 0.00084988 0 0.00084998 3.3 0.0008499 3.3 0.00085 0 0.00084992 0 0.0008500199999999999 3.3 0.00084994 3.3 0.0008500399999999999 0 0.0008499600000000001 0 0.00085006 3.3 0.0008499800000000001 3.3 0.00085008 0 0.0008500000000000001 0 0.0008501 3.3 0.00085002 3.3 0.00085012 0 0.00085004 0 0.00085014 3.3 0.00085006 3.3 0.00085016 0 0.00085008 0 0.00085018 3.3 0.0008501 3.3 0.0008502 0 0.00085012 0 0.00085022 3.3 0.00085014 3.3 0.0008502399999999999 0 0.0008501600000000001 0 0.00085026 3.3 0.0008501800000000001 3.3 0.00085028 0 0.0008502000000000001 0 0.0008503 3.3 0.0008502200000000001 3.3 0.00085032 0 0.00085024 0 0.00085034 3.3 0.00085026 3.3 0.00085036 0 0.00085028 0 0.00085038 3.3 0.0008503 3.3 0.0008504 0 0.00085032 0 0.00085042 3.3 0.00085034 3.3 0.0008504399999999999 0 0.00085036 0 0.0008504599999999999 3.3 0.0008503800000000001 3.3 0.00085048 0 0.0008504000000000001 0 0.0008505 3.3 0.0008504200000000001 3.3 0.00085052 0 0.00085044 0 0.00085054 3.3 0.00085046 3.3 0.00085056 0 0.00085048 0 0.00085058 3.3 0.0008505 3.3 0.0008506 0 0.00085052 0 0.00085062 3.3 0.00085054 3.3 0.00085064 0 0.00085056 0 0.0008506599999999999 3.3 0.0008505800000000001 3.3 0.00085068 0 0.0008506000000000001 0 0.0008507 3.3 0.0008506200000000001 3.3 0.00085072 0 0.0008506400000000001 0 0.00085074 3.3 0.00085066 3.3 0.00085076 0 0.00085068 0 0.00085078 3.3 0.0008507 3.3 0.0008508 0 0.00085072 0 0.00085082 3.3 0.00085074 3.3 0.00085084 0 0.00085076 0 0.0008508599999999999 3.3 0.00085078 3.3 0.0008508799999999999 0 0.0008508000000000001 0 0.0008509 3.3 0.0008508200000000001 3.3 0.00085092 0 0.0008508400000000001 0 0.00085094 3.3 0.00085086 3.3 0.00085096 0 0.00085088 0 0.00085098 3.3 0.0008509 3.3 0.000851 0 0.00085092 0 0.00085102 3.3 0.00085094 3.3 0.00085104 0 0.00085096 0 0.00085106 3.3 0.00085098 3.3 0.0008510799999999999 0 0.0008510000000000001 0 0.0008511 3.3 0.0008510200000000001 3.3 0.00085112 0 0.0008510400000000001 0 0.00085114 3.3 0.0008510600000000001 3.3 0.00085116 0 0.00085108 0 0.00085118 3.3 0.0008511 3.3 0.0008512 0 0.00085112 0 0.00085122 3.3 0.00085114 3.3 0.00085124 0 0.00085116 0 0.00085126 3.3 0.00085118 3.3 0.0008512799999999999 0 0.0008512 0 0.0008512999999999999 3.3 0.0008512200000000001 3.3 0.00085132 0 0.0008512400000000001 0 0.00085134 3.3 0.0008512600000000001 3.3 0.00085136 0 0.00085128 0 0.00085138 3.3 0.0008513 3.3 0.0008514 0 0.00085132 0 0.00085142 3.3 0.00085134 3.3 0.00085144 0 0.00085136 0 0.00085146 3.3 0.00085138 3.3 0.0008514799999999999 0 0.0008514 0 0.0008514999999999999 3.3 0.0008514200000000001 3.3 0.00085152 0 0.0008514400000000001 0 0.00085154 3.3 0.0008514600000000001 3.3 0.00085156 0 0.00085148 0 0.00085158 3.3 0.0008515 3.3 0.0008516 0 0.00085152 0 0.00085162 3.3 0.00085154 3.3 0.00085164 0 0.00085156 0 0.00085166 3.3 0.00085158 3.3 0.00085168 0 0.0008516 0 0.0008516999999999999 3.3 0.00085162 3.3 0.0008517199999999999 0 0.0008516400000000001 0 0.00085174 3.3 0.0008516600000000001 3.3 0.00085176 0 0.0008516800000000001 0 0.00085178 3.3 0.0008517 3.3 0.0008518 0 0.00085172 0 0.00085182 3.3 0.00085174 3.3 0.00085184 0 0.00085176 0 0.00085186 3.3 0.00085178 3.3 0.00085188 0 0.0008518 0 0.0008518999999999999 3.3 0.00085182 3.3 0.0008519199999999999 0 0.0008518400000000001 0 0.00085194 3.3 0.0008518600000000001 3.3 0.00085196 0 0.0008518800000000001 0 0.00085198 3.3 0.0008519 3.3 0.000852 0 0.00085192 0 0.00085202 3.3 0.00085194 3.3 0.00085204 0 0.00085196 0 0.00085206 3.3 0.00085198 3.3 0.00085208 0 0.000852 0 0.0008521 3.3 0.00085202 3.3 0.0008521199999999999 0 0.00085204 0 0.0008521399999999999 3.3 0.0008520600000000001 3.3 0.00085216 0 0.0008520800000000001 0 0.00085218 3.3 0.0008521000000000001 3.3 0.0008522 0 0.00085212 0 0.00085222 3.3 0.00085214 3.3 0.00085224 0 0.00085216 0 0.00085226 3.3 0.00085218 3.3 0.00085228 0 0.0008522 0 0.0008523 3.3 0.00085222 3.3 0.0008523199999999999 0 0.00085224 0 0.0008523399999999999 3.3 0.0008522600000000001 3.3 0.00085236 0 0.0008522800000000001 0 0.00085238 3.3 0.0008523000000000001 3.3 0.0008524 0 0.00085232 0 0.00085242 3.3 0.00085234 3.3 0.00085244 0 0.00085236 0 0.00085246 3.3 0.00085238 3.3 0.00085248 0 0.0008524 0 0.0008525 3.3 0.00085242 3.3 0.00085252 0 0.00085244 0 0.0008525399999999999 3.3 0.0008524600000000001 3.3 0.00085256 0 0.0008524800000000001 0 0.00085258 3.3 0.0008525000000000001 3.3 0.0008526 0 0.0008525200000000001 0 0.00085262 3.3 0.00085254 3.3 0.00085264 0 0.00085256 0 0.00085266 3.3 0.00085258 3.3 0.00085268 0 0.0008526 0 0.0008527 3.3 0.00085262 3.3 0.00085272 0 0.00085264 0 0.0008527399999999999 3.3 0.00085266 3.3 0.0008527599999999999 0 0.0008526800000000001 0 0.00085278 3.3 0.0008527000000000001 3.3 0.0008528 0 0.0008527200000000001 0 0.00085282 3.3 0.00085274 3.3 0.00085284 0 0.00085276 0 0.00085286 3.3 0.00085278 3.3 0.00085288 0 0.0008528 0 0.0008529 3.3 0.00085282 3.3 0.00085292 0 0.00085284 0 0.00085294 3.3 0.00085286 3.3 0.0008529599999999999 0 0.0008528800000000001 0 0.00085298 3.3 0.0008529000000000001 3.3 0.000853 0 0.0008529200000000001 0 0.00085302 3.3 0.0008529400000000001 3.3 0.00085304 0 0.00085296 0 0.00085306 3.3 0.00085298 3.3 0.00085308 0 0.000853 0 0.0008531 3.3 0.00085302 3.3 0.00085312 0 0.00085304 0 0.00085314 3.3 0.00085306 3.3 0.0008531599999999999 0 0.00085308 0 0.0008531799999999999 3.3 0.0008531000000000001 3.3 0.0008532 0 0.0008531200000000001 0 0.00085322 3.3 0.0008531400000000001 3.3 0.00085324 0 0.00085316 0 0.00085326 3.3 0.00085318 3.3 0.00085328 0 0.0008532 0 0.0008533 3.3 0.00085322 3.3 0.00085332 0 0.00085324 0 0.00085334 3.3 0.00085326 3.3 0.00085336 0 0.00085328 0 0.0008533799999999999 3.3 0.0008533000000000001 3.3 0.0008534 0 0.0008533200000000001 0 0.00085342 3.3 0.0008533400000000001 3.3 0.00085344 0 0.0008533600000000001 0 0.00085346 3.3 0.00085338 3.3 0.00085348 0 0.0008534 0 0.0008535 3.3 0.00085342 3.3 0.00085352 0 0.00085344 0 0.00085354 3.3 0.00085346 3.3 0.00085356 0 0.00085348 0 0.0008535799999999999 3.3 0.0008535 3.3 0.0008535999999999999 0 0.0008535200000000001 0 0.00085362 3.3 0.0008535400000000001 3.3 0.00085364 0 0.0008535600000000001 0 0.00085366 3.3 0.00085358 3.3 0.00085368 0 0.0008536 0 0.0008537 3.3 0.00085362 3.3 0.00085372 0 0.00085364 0 0.00085374 3.3 0.00085366 3.3 0.00085376 0 0.00085368 0 0.00085378 3.3 0.0008537 3.3 0.0008537999999999999 0 0.0008537200000000001 0 0.00085382 3.3 0.0008537400000000001 3.3 0.00085384 0 0.0008537600000000001 0 0.00085386 3.3 0.0008537800000000001 3.3 0.00085388 0 0.0008538 0 0.0008539 3.3 0.00085382 3.3 0.00085392 0 0.00085384 0 0.00085394 3.3 0.00085386 3.3 0.00085396 0 0.00085388 0 0.00085398 3.3 0.0008539 3.3 0.0008539999999999999 0 0.00085392 0 0.0008540199999999999 3.3 0.0008539400000000001 3.3 0.00085404 0 0.0008539600000000001 0 0.00085406 3.3 0.0008539800000000001 3.3 0.00085408 0 0.000854 0 0.0008541 3.3 0.00085402 3.3 0.00085412 0 0.00085404 0 0.00085414 3.3 0.00085406 3.3 0.00085416 0 0.00085408 0 0.00085418 3.3 0.0008541 3.3 0.0008542 0 0.00085412 0 0.0008542199999999999 3.3 0.0008541400000000001 3.3 0.00085424 0 0.0008541600000000001 0 0.00085426 3.3 0.0008541800000000001 3.3 0.00085428 0 0.0008542000000000001 0 0.0008543 3.3 0.00085422 3.3 0.00085432 0 0.00085424 0 0.00085434 3.3 0.00085426 3.3 0.00085436 0 0.00085428 0 0.00085438 3.3 0.0008543 3.3 0.0008544 0 0.00085432 0 0.0008544199999999999 3.3 0.00085434 3.3 0.0008544399999999999 0 0.0008543600000000001 0 0.00085446 3.3 0.0008543800000000001 3.3 0.00085448 0 0.0008544000000000001 0 0.0008545 3.3 0.00085442 3.3 0.00085452 0 0.00085444 0 0.00085454 3.3 0.00085446 3.3 0.00085456 0 0.00085448 0 0.00085458 3.3 0.0008545 3.3 0.0008546 0 0.00085452 0 0.0008546199999999999 3.3 0.00085454 3.3 0.0008546399999999999 0 0.0008545600000000001 0 0.00085466 3.3 0.0008545800000000001 3.3 0.00085468 0 0.0008546000000000001 0 0.0008547 3.3 0.00085462 3.3 0.00085472 0 0.00085464 0 0.00085474 3.3 0.00085466 3.3 0.00085476 0 0.00085468 0 0.00085478 3.3 0.0008547 3.3 0.0008548 0 0.00085472 0 0.00085482 3.3 0.00085474 3.3 0.0008548399999999999 0 0.00085476 0 0.0008548599999999999 3.3 0.0008547800000000001 3.3 0.00085488 0 0.0008548000000000001 0 0.0008549 3.3 0.0008548200000000001 3.3 0.00085492 0 0.00085484 0 0.00085494 3.3 0.00085486 3.3 0.00085496 0 0.00085488 0 0.00085498 3.3 0.0008549 3.3 0.000855 0 0.00085492 0 0.00085502 3.3 0.00085494 3.3 0.0008550399999999999 0 0.00085496 0 0.0008550599999999999 3.3 0.0008549800000000001 3.3 0.00085508 0 0.0008550000000000001 0 0.0008551 3.3 0.0008550200000000001 3.3 0.00085512 0 0.00085504 0 0.00085514 3.3 0.00085506 3.3 0.00085516 0 0.00085508 0 0.00085518 3.3 0.0008551 3.3 0.0008552 0 0.00085512 0 0.00085522 3.3 0.00085514 3.3 0.00085524 0 0.00085516 0 0.0008552599999999999 3.3 0.00085518 3.3 0.0008552799999999999 0 0.0008552000000000001 0 0.0008553 3.3 0.0008552200000000001 3.3 0.00085532 0 0.0008552400000000001 0 0.00085534 3.3 0.00085526 3.3 0.00085536 0 0.00085528 0 0.00085538 3.3 0.0008553 3.3 0.0008554 0 0.00085532 0 0.00085542 3.3 0.00085534 3.3 0.00085544 0 0.00085536 0 0.0008554599999999999 3.3 0.00085538 3.3 0.0008554799999999999 0 0.0008554000000000001 0 0.0008555 3.3 0.0008554200000000001 3.3 0.00085552 0 0.0008554400000000001 0 0.00085554 3.3 0.00085546 3.3 0.00085556 0 0.00085548 0 0.00085558 3.3 0.0008555 3.3 0.0008556 0 0.00085552 0 0.00085562 3.3 0.00085554 3.3 0.00085564 0 0.00085556 0 0.00085566 3.3 0.00085558 3.3 0.0008556799999999999 0 0.0008556000000000001 0 0.0008557 3.3 0.0008556200000000001 3.3 0.00085572 0 0.0008556400000000001 0 0.00085574 3.3 0.0008556600000000001 3.3 0.00085576 0 0.00085568 0 0.00085578 3.3 0.0008557 3.3 0.0008558 0 0.00085572 0 0.00085582 3.3 0.00085574 3.3 0.00085584 0 0.00085576 0 0.00085586 3.3 0.00085578 3.3 0.0008558799999999999 0 0.0008558 0 0.0008558999999999999 3.3 0.0008558200000000001 3.3 0.00085592 0 0.0008558400000000001 0 0.00085594 3.3 0.0008558600000000001 3.3 0.00085596 0 0.00085588 0 0.00085598 3.3 0.0008559 3.3 0.000856 0 0.00085592 0 0.00085602 3.3 0.00085594 3.3 0.00085604 0 0.00085596 0 0.00085606 3.3 0.00085598 3.3 0.00085608 0 0.000856 0 0.0008560999999999999 3.3 0.0008560200000000001 3.3 0.00085612 0 0.0008560400000000001 0 0.00085614 3.3 0.0008560600000000001 3.3 0.00085616 0 0.0008560800000000001 0 0.00085618 3.3 0.0008561 3.3 0.0008562 0 0.00085612 0 0.00085622 3.3 0.00085614 3.3 0.00085624 0 0.00085616 0 0.00085626 3.3 0.00085618 3.3 0.00085628 0 0.0008562 0 0.0008562999999999999 3.3 0.00085622 3.3 0.0008563199999999999 0 0.0008562400000000001 0 0.00085634 3.3 0.0008562600000000001 3.3 0.00085636 0 0.0008562800000000001 0 0.00085638 3.3 0.0008563 3.3 0.0008564 0 0.00085632 0 0.00085642 3.3 0.00085634 3.3 0.00085644 0 0.00085636 0 0.00085646 3.3 0.00085638 3.3 0.00085648 0 0.0008564 0 0.0008565 3.3 0.00085642 3.3 0.0008565199999999999 0 0.0008564400000000001 0 0.00085654 3.3 0.0008564600000000001 3.3 0.00085656 0 0.0008564800000000001 0 0.00085658 3.3 0.0008565000000000001 3.3 0.0008566 0 0.00085652 0 0.00085662 3.3 0.00085654 3.3 0.00085664 0 0.00085656 0 0.00085666 3.3 0.00085658 3.3 0.00085668 0 0.0008566 0 0.0008567 3.3 0.00085662 3.3 0.0008567199999999999 0 0.00085664 0 0.0008567399999999999 3.3 0.0008566600000000001 3.3 0.00085676 0 0.0008566800000000001 0 0.00085678 3.3 0.0008567000000000001 3.3 0.0008568 0 0.00085672 0 0.00085682 3.3 0.00085674 3.3 0.00085684 0 0.00085676 0 0.00085686 3.3 0.00085678 3.3 0.00085688 0 0.0008568 0 0.0008569 3.3 0.00085682 3.3 0.00085692 0 0.00085684 0 0.0008569399999999999 3.3 0.0008568600000000001 3.3 0.00085696 0 0.0008568800000000001 0 0.00085698 3.3 0.0008569000000000001 3.3 0.000857 0 0.0008569200000000001 0 0.00085702 3.3 0.00085694 3.3 0.00085704 0 0.00085696 0 0.00085706 3.3 0.00085698 3.3 0.00085708 0 0.000857 0 0.0008571 3.3 0.00085702 3.3 0.00085712 0 0.00085704 0 0.0008571399999999999 3.3 0.00085706 3.3 0.0008571599999999999 0 0.0008570800000000001 0 0.00085718 3.3 0.0008571000000000001 3.3 0.0008572 0 0.0008571200000000001 0 0.00085722 3.3 0.00085714 3.3 0.00085724 0 0.00085716 0 0.00085726 3.3 0.00085718 3.3 0.00085728 0 0.0008572 0 0.0008573 3.3 0.00085722 3.3 0.00085732 0 0.00085724 0 0.00085734 3.3 0.00085726 3.3 0.0008573599999999999 0 0.0008572800000000001 0 0.00085738 3.3 0.0008573000000000001 3.3 0.0008574 0 0.0008573200000000001 0 0.00085742 3.3 0.0008573400000000001 3.3 0.00085744 0 0.00085736 0 0.00085746 3.3 0.00085738 3.3 0.00085748 0 0.0008574 0 0.0008575 3.3 0.00085742 3.3 0.00085752 0 0.00085744 0 0.00085754 3.3 0.00085746 3.3 0.0008575599999999999 0 0.00085748 0 0.0008575799999999999 3.3 0.0008575000000000001 3.3 0.0008576 0 0.0008575200000000001 0 0.00085762 3.3 0.0008575400000000001 3.3 0.00085764 0 0.00085756 0 0.00085766 3.3 0.00085758 3.3 0.00085768 0 0.0008576 0 0.0008577 3.3 0.00085762 3.3 0.00085772 0 0.00085764 0 0.00085774 3.3 0.00085766 3.3 0.00085776 0 0.00085768 0 0.0008577799999999999 3.3 0.0008577000000000001 3.3 0.0008578 0 0.0008577200000000001 0 0.00085782 3.3 0.0008577400000000001 3.3 0.00085784 0 0.0008577600000000001 0 0.00085786 3.3 0.00085778 3.3 0.00085788 0 0.0008578 0 0.0008579 3.3 0.00085782 3.3 0.00085792 0 0.00085784 0 0.00085794 3.3 0.00085786 3.3 0.00085796 0 0.00085788 0 0.0008579799999999999 3.3 0.0008579 3.3 0.0008579999999999999 0 0.0008579200000000001 0 0.00085802 3.3 0.0008579400000000001 3.3 0.00085804 0 0.0008579600000000001 0 0.00085806 3.3 0.00085798 3.3 0.00085808 0 0.000858 0 0.0008581 3.3 0.00085802 3.3 0.00085812 0 0.00085804 0 0.00085814 3.3 0.00085806 3.3 0.00085816 0 0.00085808 0 0.0008581799999999999 3.3 0.0008581 3.3 0.0008581999999999999 0 0.0008581200000000001 0 0.00085822 3.3 0.0008581400000000001 3.3 0.00085824 0 0.0008581600000000001 0 0.00085826 3.3 0.00085818 3.3 0.00085828 0 0.0008582 0 0.0008583 3.3 0.00085822 3.3 0.00085832 0 0.00085824 0 0.00085834 3.3 0.00085826 3.3 0.00085836 0 0.00085828 0 0.00085838 3.3 0.0008583 3.3 0.0008583999999999999 0 0.00085832 0 0.0008584199999999999 3.3 0.0008583400000000001 3.3 0.00085844 0 0.0008583600000000001 0 0.00085846 3.3 0.0008583800000000001 3.3 0.00085848 0 0.0008584 0 0.0008585 3.3 0.00085842 3.3 0.00085852 0 0.00085844 0 0.00085854 3.3 0.00085846 3.3 0.00085856 0 0.00085848 0 0.00085858 3.3 0.0008585 3.3 0.0008585999999999999 0 0.00085852 0 0.0008586199999999999 3.3 0.0008585400000000001 3.3 0.00085864 0 0.0008585600000000001 0 0.00085866 3.3 0.0008585800000000001 3.3 0.00085868 0 0.0008586 0 0.0008587 3.3 0.00085862 3.3 0.00085872 0 0.00085864 0 0.00085874 3.3 0.00085866 3.3 0.00085876 0 0.00085868 0 0.00085878 3.3 0.0008587 3.3 0.0008588 0 0.00085872 0 0.0008588199999999999 3.3 0.00085874 3.3 0.0008588399999999999 0 0.0008587600000000001 0 0.00085886 3.3 0.0008587800000000001 3.3 0.00085888 0 0.0008588000000000001 0 0.0008589 3.3 0.00085882 3.3 0.00085892 0 0.00085884 0 0.00085894 3.3 0.00085886 3.3 0.00085896 0 0.00085888 0 0.00085898 3.3 0.0008589 3.3 0.000859 0 0.00085892 0 0.0008590199999999999 3.3 0.00085894 3.3 0.0008590399999999999 0 0.0008589600000000001 0 0.00085906 3.3 0.0008589800000000001 3.3 0.00085908 0 0.0008590000000000001 0 0.0008591 3.3 0.00085902 3.3 0.00085912 0 0.00085904 0 0.00085914 3.3 0.00085906 3.3 0.00085916 0 0.00085908 0 0.00085918 3.3 0.0008591 3.3 0.0008592 0 0.00085912 0 0.00085922 3.3 0.00085914 3.3 0.0008592399999999999 0 0.0008591600000000001 0 0.00085926 3.3 0.0008591800000000001 3.3 0.00085928 0 0.0008592000000000001 0 0.0008593 3.3 0.0008592200000000001 3.3 0.00085932 0 0.00085924 0 0.00085934 3.3 0.00085926 3.3 0.00085936 0 0.00085928 0 0.00085938 3.3 0.0008593 3.3 0.0008594 0 0.00085932 0 0.00085942 3.3 0.00085934 3.3 0.0008594399999999999 0 0.00085936 0 0.0008594599999999999 3.3 0.0008593800000000001 3.3 0.00085948 0 0.0008594000000000001 0 0.0008595 3.3 0.0008594200000000001 3.3 0.00085952 0 0.00085944 0 0.00085954 3.3 0.00085946 3.3 0.00085956 0 0.00085948 0 0.00085958 3.3 0.0008595 3.3 0.0008596 0 0.00085952 0 0.00085962 3.3 0.00085954 3.3 0.00085964 0 0.00085956 0 0.0008596599999999999 3.3 0.0008595800000000001 3.3 0.00085968 0 0.0008596000000000001 0 0.0008597 3.3 0.0008596200000000001 3.3 0.00085972 0 0.0008596400000000001 0 0.00085974 3.3 0.00085966 3.3 0.00085976 0 0.00085968 0 0.00085978 3.3 0.0008597 3.3 0.0008598 0 0.00085972 0 0.00085982 3.3 0.00085974 3.3 0.00085984 0 0.00085976 0 0.0008598599999999999 3.3 0.00085978 3.3 0.0008598799999999999 0 0.0008598000000000001 0 0.0008599 3.3 0.0008598200000000001 3.3 0.00085992 0 0.0008598400000000001 0 0.00085994 3.3 0.00085986 3.3 0.00085996 0 0.00085988 0 0.00085998 3.3 0.0008599 3.3 0.00086 0 0.00085992 0 0.00086002 3.3 0.00085994 3.3 0.00086004 0 0.00085996 0 0.00086006 3.3 0.00085998 3.3 0.0008600799999999999 0 0.0008600000000000001 0 0.0008601 3.3 0.0008600200000000001 3.3 0.00086012 0 0.0008600400000000001 0 0.00086014 3.3 0.0008600600000000001 3.3 0.00086016 0 0.00086008 0 0.00086018 3.3 0.0008601 3.3 0.0008602 0 0.00086012 0 0.00086022 3.3 0.00086014 3.3 0.00086024 0 0.00086016 0 0.00086026 3.3 0.00086018 3.3 0.0008602799999999999 0 0.0008602 0 0.0008602999999999999 3.3 0.0008602200000000001 3.3 0.00086032 0 0.0008602400000000001 0 0.00086034 3.3 0.0008602600000000001 3.3 0.00086036 0 0.00086028 0 0.00086038 3.3 0.0008603 3.3 0.0008604 0 0.00086032 0 0.00086042 3.3 0.00086034 3.3 0.00086044 0 0.00086036 0 0.00086046 3.3 0.00086038 3.3 0.00086048 0 0.0008604 0 0.0008604999999999999 3.3 0.0008604200000000001 3.3 0.00086052 0 0.0008604400000000001 0 0.00086054 3.3 0.0008604600000000001 3.3 0.00086056 0 0.0008604800000000001 0 0.00086058 3.3 0.0008605 3.3 0.0008606 0 0.00086052 0 0.00086062 3.3 0.00086054 3.3 0.00086064 0 0.00086056 0 0.00086066 3.3 0.00086058 3.3 0.00086068 0 0.0008606 0 0.0008606999999999999 3.3 0.00086062 3.3 0.0008607199999999999 0 0.0008606400000000001 0 0.00086074 3.3 0.0008606600000000001 3.3 0.00086076 0 0.0008606800000000001 0 0.00086078 3.3 0.0008607 3.3 0.0008608 0 0.00086072 0 0.00086082 3.3 0.00086074 3.3 0.00086084 0 0.00086076 0 0.00086086 3.3 0.00086078 3.3 0.00086088 0 0.0008608 0 0.0008609 3.3 0.00086082 3.3 0.0008609199999999999 0 0.0008608400000000001 0 0.00086094 3.3 0.0008608600000000001 3.3 0.00086096 0 0.0008608800000000001 0 0.00086098 3.3 0.0008609000000000001 3.3 0.000861 0 0.00086092 0 0.00086102 3.3 0.00086094 3.3 0.00086104 0 0.00086096 0 0.00086106 3.3 0.00086098 3.3 0.00086108 0 0.000861 0 0.0008611 3.3 0.00086102 3.3 0.0008611199999999999 0 0.00086104 0 0.0008611399999999999 3.3 0.0008610600000000001 3.3 0.00086116 0 0.0008610800000000001 0 0.00086118 3.3 0.0008611000000000001 3.3 0.0008612 0 0.00086112 0 0.00086122 3.3 0.00086114 3.3 0.00086124 0 0.00086116 0 0.00086126 3.3 0.00086118 3.3 0.00086128 0 0.0008612 0 0.0008613 3.3 0.00086122 3.3 0.00086132 0 0.00086124 0 0.0008613399999999999 3.3 0.0008612600000000001 3.3 0.00086136 0 0.0008612800000000001 0 0.00086138 3.3 0.0008613000000000001 3.3 0.0008614 0 0.0008613200000000001 0 0.00086142 3.3 0.00086134 3.3 0.00086144 0 0.00086136 0 0.00086146 3.3 0.00086138 3.3 0.00086148 0 0.0008614 0 0.0008615 3.3 0.00086142 3.3 0.00086152 0 0.00086144 0 0.0008615399999999999 3.3 0.00086146 3.3 0.0008615599999999999 0 0.0008614800000000001 0 0.00086158 3.3 0.0008615000000000001 3.3 0.0008616 0 0.0008615200000000001 0 0.00086162 3.3 0.00086154 3.3 0.00086164 0 0.00086156 0 0.00086166 3.3 0.00086158 3.3 0.00086168 0 0.0008616 0 0.0008617 3.3 0.00086162 3.3 0.00086172 0 0.00086164 0 0.0008617399999999999 3.3 0.00086166 3.3 0.0008617599999999999 0 0.0008616800000000001 0 0.00086178 3.3 0.0008617000000000001 3.3 0.0008618 0 0.0008617200000000001 0 0.00086182 3.3 0.00086174 3.3 0.00086184 0 0.00086176 0 0.00086186 3.3 0.00086178 3.3 0.00086188 0 0.0008618 0 0.0008619 3.3 0.00086182 3.3 0.00086192 0 0.00086184 0 0.00086194 3.3 0.00086186 3.3 0.0008619599999999999 0 0.00086188 0 0.0008619799999999999 3.3 0.0008619000000000001 3.3 0.000862 0 0.0008619200000000001 0 0.00086202 3.3 0.0008619400000000001 3.3 0.00086204 0 0.00086196 0 0.00086206 3.3 0.00086198 3.3 0.00086208 0 0.000862 0 0.0008621 3.3 0.00086202 3.3 0.00086212 0 0.00086204 0 0.00086214 3.3 0.00086206 3.3 0.0008621599999999999 0 0.00086208 0 0.0008621799999999999 3.3 0.0008621000000000001 3.3 0.0008622 0 0.0008621200000000001 0 0.00086222 3.3 0.0008621400000000001 3.3 0.00086224 0 0.00086216 0 0.00086226 3.3 0.00086218 3.3 0.00086228 0 0.0008622 0 0.0008623 3.3 0.00086222 3.3 0.00086232 0 0.00086224 0 0.00086234 3.3 0.00086226 3.3 0.00086236 0 0.00086228 0 0.0008623799999999999 3.3 0.0008623 3.3 0.0008623999999999999 0 0.0008623200000000001 0 0.00086242 3.3 0.0008623400000000001 3.3 0.00086244 0 0.0008623600000000001 0 0.00086246 3.3 0.00086238 3.3 0.00086248 0 0.0008624 0 0.0008625 3.3 0.00086242 3.3 0.00086252 0 0.00086244 0 0.00086254 3.3 0.00086246 3.3 0.00086256 0 0.00086248 0 0.0008625799999999999 3.3 0.0008625 3.3 0.0008625999999999999 0 0.0008625200000000001 0 0.00086262 3.3 0.0008625400000000001 3.3 0.00086264 0 0.0008625600000000001 0 0.00086266 3.3 0.00086258 3.3 0.00086268 0 0.0008626 0 0.0008627 3.3 0.00086262 3.3 0.00086272 0 0.00086264 0 0.00086274 3.3 0.00086266 3.3 0.00086276 0 0.00086268 0 0.00086278 3.3 0.0008627 3.3 0.0008627999999999999 0 0.0008627200000000001 0 0.00086282 3.3 0.0008627400000000001 3.3 0.00086284 0 0.0008627600000000001 0 0.00086286 3.3 0.0008627800000000001 3.3 0.00086288 0 0.0008628 0 0.0008629 3.3 0.00086282 3.3 0.00086292 0 0.00086284 0 0.00086294 3.3 0.00086286 3.3 0.00086296 0 0.00086288 0 0.00086298 3.3 0.0008629 3.3 0.0008629999999999999 0 0.00086292 0 0.0008630199999999999 3.3 0.0008629400000000001 3.3 0.00086304 0 0.0008629600000000001 0 0.00086306 3.3 0.0008629800000000001 3.3 0.00086308 0 0.000863 0 0.0008631 3.3 0.00086302 3.3 0.00086312 0 0.00086304 0 0.00086314 3.3 0.00086306 3.3 0.00086316 0 0.00086308 0 0.00086318 3.3 0.0008631 3.3 0.0008632 0 0.00086312 0 0.0008632199999999999 3.3 0.0008631400000000001 3.3 0.00086324 0 0.0008631600000000001 0 0.00086326 3.3 0.0008631800000000001 3.3 0.00086328 0 0.0008632000000000001 0 0.0008633 3.3 0.00086322 3.3 0.00086332 0 0.00086324 0 0.00086334 3.3 0.00086326 3.3 0.00086336 0 0.00086328 0 0.00086338 3.3 0.0008633 3.3 0.0008634 0 0.00086332 0 0.0008634199999999999 3.3 0.00086334 3.3 0.0008634399999999999 0 0.0008633600000000001 0 0.00086346 3.3 0.0008633800000000001 3.3 0.00086348 0 0.0008634000000000001 0 0.0008635 3.3 0.00086342 3.3 0.00086352 0 0.00086344 0 0.00086354 3.3 0.00086346 3.3 0.00086356 0 0.00086348 0 0.00086358 3.3 0.0008635 3.3 0.0008636 0 0.00086352 0 0.00086362 3.3 0.00086354 3.3 0.0008636399999999999 0 0.0008635600000000001 0 0.00086366 3.3 0.0008635800000000001 3.3 0.00086368 0 0.0008636000000000001 0 0.0008637 3.3 0.0008636200000000001 3.3 0.00086372 0 0.00086364 0 0.00086374 3.3 0.00086366 3.3 0.00086376 0 0.00086368 0 0.00086378 3.3 0.0008637 3.3 0.0008638 0 0.00086372 0 0.00086382 3.3 0.00086374 3.3 0.0008638399999999999 0 0.00086376 0 0.0008638599999999999 3.3 0.0008637800000000001 3.3 0.00086388 0 0.0008638000000000001 0 0.0008639 3.3 0.0008638200000000001 3.3 0.00086392 0 0.00086384 0 0.00086394 3.3 0.00086386 3.3 0.00086396 0 0.00086388 0 0.00086398 3.3 0.0008639 3.3 0.000864 0 0.00086392 0 0.00086402 3.3 0.00086394 3.3 0.00086404 0 0.00086396 0 0.0008640599999999999 3.3 0.0008639800000000001 3.3 0.00086408 0 0.0008640000000000001 0 0.0008641 3.3 0.0008640200000000001 3.3 0.00086412 0 0.0008640400000000001 0 0.00086414 3.3 0.00086406 3.3 0.00086416 0 0.00086408 0 0.00086418 3.3 0.0008641 3.3 0.0008642 0 0.00086412 0 0.00086422 3.3 0.00086414 3.3 0.00086424 0 0.00086416 0 0.0008642599999999999 3.3 0.00086418 3.3 0.0008642799999999999 0 0.0008642000000000001 0 0.0008643 3.3 0.0008642200000000001 3.3 0.00086432 0 0.0008642400000000001 0 0.00086434 3.3 0.00086426 3.3 0.00086436 0 0.00086428 0 0.00086438 3.3 0.0008643 3.3 0.0008644 0 0.00086432 0 0.00086442 3.3 0.00086434 3.3 0.00086444 0 0.00086436 0 0.00086446 3.3 0.00086438 3.3 0.0008644799999999999 0 0.0008644000000000001 0 0.0008645 3.3 0.0008644200000000001 3.3 0.00086452 0 0.0008644400000000001 0 0.00086454 3.3 0.0008644600000000001 3.3 0.00086456 0 0.00086448 0 0.00086458 3.3 0.0008645 3.3 0.0008646 0 0.00086452 0 0.00086462 3.3 0.00086454 3.3 0.00086464 0 0.00086456 0 0.00086466 3.3 0.00086458 3.3 0.0008646799999999999 0 0.0008646 0 0.0008646999999999999 3.3 0.0008646200000000001 3.3 0.00086472 0 0.0008646400000000001 0 0.00086474 3.3 0.0008646600000000001 3.3 0.00086476 0 0.00086468 0 0.00086478 3.3 0.0008647 3.3 0.0008648 0 0.00086472 0 0.00086482 3.3 0.00086474 3.3 0.00086484 0 0.00086476 0 0.00086486 3.3 0.00086478 3.3 0.0008648799999999999 0 0.0008648 0 0.0008648999999999999 3.3 0.0008648200000000001 3.3 0.00086492 0 0.0008648400000000001 0 0.00086494 3.3 0.0008648600000000001 3.3 0.00086496 0 0.00086488 0 0.00086498 3.3 0.0008649 3.3 0.000865 0 0.00086492 0 0.00086502 3.3 0.00086494 3.3 0.00086504 0 0.00086496 0 0.00086506 3.3 0.00086498 3.3 0.00086508 0 0.000865 0 0.0008650999999999999 3.3 0.00086502 3.3 0.0008651199999999999 0 0.0008650400000000001 0 0.00086514 3.3 0.0008650600000000001 3.3 0.00086516 0 0.0008650800000000001 0 0.00086518 3.3 0.0008651 3.3 0.0008652 0 0.00086512 0 0.00086522 3.3 0.00086514 3.3 0.00086524 0 0.00086516 0 0.00086526 3.3 0.00086518 3.3 0.00086528 0 0.0008652 0 0.0008652999999999999 3.3 0.00086522 3.3 0.0008653199999999999 0 0.0008652400000000001 0 0.00086534 3.3 0.0008652600000000001 3.3 0.00086536 0 0.0008652800000000001 0 0.00086538 3.3 0.0008653 3.3 0.0008654 0 0.00086532 0 0.00086542 3.3 0.00086534 3.3 0.00086544 0 0.00086536 0 0.00086546 3.3 0.00086538 3.3 0.00086548 0 0.0008654 0 0.0008655 3.3 0.00086542 3.3 0.0008655199999999999 0 0.00086544 0 0.0008655399999999999 3.3 0.0008654600000000001 3.3 0.00086556 0 0.0008654800000000001 0 0.00086558 3.3 0.0008655000000000001 3.3 0.0008656 0 0.00086552 0 0.00086562 3.3 0.00086554 3.3 0.00086564 0 0.00086556 0 0.00086566 3.3 0.00086558 3.3 0.00086568 0 0.0008656 0 0.0008657 3.3 0.00086562 3.3 0.0008657199999999999 0 0.00086564 0 0.0008657399999999999 3.3 0.0008656600000000001 3.3 0.00086576 0 0.0008656800000000001 0 0.00086578 3.3 0.0008657000000000001 3.3 0.0008658 0 0.00086572 0 0.00086582 3.3 0.00086574 3.3 0.00086584 0 0.00086576 0 0.00086586 3.3 0.00086578 3.3 0.00086588 0 0.0008658 0 0.0008659 3.3 0.00086582 3.3 0.00086592 0 0.00086584 0 0.0008659399999999999 3.3 0.00086586 3.3 0.0008659599999999999 0 0.0008658800000000001 0 0.00086598 3.3 0.0008659000000000001 3.3 0.000866 0 0.0008659200000000001 0 0.00086602 3.3 0.00086594 3.3 0.00086604 0 0.00086596 0 0.00086606 3.3 0.00086598 3.3 0.00086608 0 0.000866 0 0.0008661 3.3 0.00086602 3.3 0.00086612 0 0.00086604 0 0.0008661399999999999 3.3 0.00086606 3.3 0.0008661599999999999 0 0.0008660800000000001 0 0.00086618 3.3 0.0008661000000000001 3.3 0.0008662 0 0.0008661200000000001 0 0.00086622 3.3 0.00086614 3.3 0.00086624 0 0.00086616 0 0.00086626 3.3 0.00086618 3.3 0.00086628 0 0.0008662 0 0.0008663 3.3 0.00086622 3.3 0.00086632 0 0.00086624 0 0.00086634 3.3 0.00086626 3.3 0.0008663599999999999 0 0.0008662800000000001 0 0.00086638 3.3 0.0008663000000000001 3.3 0.0008664 0 0.0008663200000000001 0 0.00086642 3.3 0.0008663400000000001 3.3 0.00086644 0 0.00086636 0 0.00086646 3.3 0.00086638 3.3 0.00086648 0 0.0008664 0 0.0008665 3.3 0.00086642 3.3 0.00086652 0 0.00086644 0 0.00086654 3.3 0.00086646 3.3 0.0008665599999999999 0 0.00086648 0 0.0008665799999999999 3.3 0.0008665000000000001 3.3 0.0008666 0 0.0008665200000000001 0 0.00086662 3.3 0.0008665400000000001 3.3 0.00086664 0 0.00086656 0 0.00086666 3.3 0.00086658 3.3 0.00086668 0 0.0008666 0 0.0008667 3.3 0.00086662 3.3 0.00086672 0 0.00086664 0 0.00086674 3.3 0.00086666 3.3 0.00086676 0 0.00086668 0 0.0008667799999999999 3.3 0.0008667000000000001 3.3 0.0008668 0 0.0008667200000000001 0 0.00086682 3.3 0.0008667400000000001 3.3 0.00086684 0 0.0008667600000000001 0 0.00086686 3.3 0.00086678 3.3 0.00086688 0 0.0008668 0 0.0008669 3.3 0.00086682 3.3 0.00086692 0 0.00086684 0 0.00086694 3.3 0.00086686 3.3 0.00086696 0 0.00086688 0 0.0008669799999999999 3.3 0.0008669 3.3 0.0008669999999999999 0 0.0008669200000000001 0 0.00086702 3.3 0.0008669400000000001 3.3 0.00086704 0 0.0008669600000000001 0 0.00086706 3.3 0.00086698 3.3 0.00086708 0 0.000867 0 0.0008671 3.3 0.00086702 3.3 0.00086712 0 0.00086704 0 0.00086714 3.3 0.00086706 3.3 0.00086716 0 0.00086708 0 0.00086718 3.3 0.0008671 3.3 0.0008671999999999999 0 0.0008671200000000001 0 0.00086722 3.3 0.0008671400000000001 3.3 0.00086724 0 0.0008671600000000001 0 0.00086726 3.3 0.0008671800000000001 3.3 0.00086728 0 0.0008672 0 0.0008673 3.3 0.00086722 3.3 0.00086732 0 0.00086724 0 0.00086734 3.3 0.00086726 3.3 0.00086736 0 0.00086728 0 0.00086738 3.3 0.0008673 3.3 0.0008673999999999999 0 0.00086732 0 0.0008674199999999999 3.3 0.0008673400000000001 3.3 0.00086744 0 0.0008673600000000001 0 0.00086746 3.3 0.0008673800000000001 3.3 0.00086748 0 0.0008674 0 0.0008675 3.3 0.00086742 3.3 0.00086752 0 0.00086744 0 0.00086754 3.3 0.00086746 3.3 0.00086756 0 0.00086748 0 0.00086758 3.3 0.0008675 3.3 0.0008676 0 0.00086752 0 0.0008676199999999999 3.3 0.0008675400000000001 3.3 0.00086764 0 0.0008675600000000001 0 0.00086766 3.3 0.0008675800000000001 3.3 0.00086768 0 0.0008676000000000001 0 0.0008677 3.3 0.00086762 3.3 0.00086772 0 0.00086764 0 0.00086774 3.3 0.00086766 3.3 0.00086776 0 0.00086768 0 0.00086778 3.3 0.0008677 3.3 0.0008678 0 0.00086772 0 0.0008678199999999999 3.3 0.00086774 3.3 0.0008678399999999999 0 0.0008677600000000001 0 0.00086786 3.3 0.0008677800000000001 3.3 0.00086788 0 0.0008678000000000001 0 0.0008679 3.3 0.00086782 3.3 0.00086792 0 0.00086784 0 0.00086794 3.3 0.00086786 3.3 0.00086796 0 0.00086788 0 0.00086798 3.3 0.0008679 3.3 0.000868 0 0.00086792 0 0.00086802 3.3 0.00086794 3.3 0.0008680399999999999 0 0.0008679600000000001 0 0.00086806 3.3 0.0008679800000000001 3.3 0.00086808 0 0.0008680000000000001 0 0.0008681 3.3 0.0008680200000000001 3.3 0.00086812 0 0.00086804 0 0.00086814 3.3 0.00086806 3.3 0.00086816 0 0.00086808 0 0.00086818 3.3 0.0008681 3.3 0.0008682 0 0.00086812 0 0.00086822 3.3 0.00086814 3.3 0.0008682399999999999 0 0.00086816 0 0.0008682599999999999 3.3 0.0008681800000000001 3.3 0.00086828 0 0.0008682000000000001 0 0.0008683 3.3 0.0008682200000000001 3.3 0.00086832 0 0.00086824 0 0.00086834 3.3 0.00086826 3.3 0.00086836 0 0.00086828 0 0.00086838 3.3 0.0008683 3.3 0.0008684 0 0.00086832 0 0.00086842 3.3 0.00086834 3.3 0.0008684399999999999 0 0.00086836 0 0.0008684599999999999 3.3 0.0008683800000000001 3.3 0.00086848 0 0.0008684000000000001 0 0.0008685 3.3 0.0008684200000000001 3.3 0.00086852 0 0.00086844 0 0.00086854 3.3 0.00086846 3.3 0.00086856 0 0.00086848 0 0.00086858 3.3 0.0008685 3.3 0.0008686 0 0.00086852 0 0.00086862 3.3 0.00086854 3.3 0.00086864 0 0.00086856 0 0.0008686599999999999 3.3 0.00086858 3.3 0.0008686799999999999 0 0.0008686000000000001 0 0.0008687 3.3 0.0008686200000000001 3.3 0.00086872 0 0.0008686400000000001 0 0.00086874 3.3 0.00086866 3.3 0.00086876 0 0.00086868 0 0.00086878 3.3 0.0008687 3.3 0.0008688 0 0.00086872 0 0.00086882 3.3 0.00086874 3.3 0.00086884 0 0.00086876 0 0.0008688599999999999 3.3 0.00086878 3.3 0.0008688799999999999 0 0.0008688000000000001 0 0.0008689 3.3 0.0008688200000000001 3.3 0.00086892 0 0.0008688400000000001 0 0.00086894 3.3 0.00086886 3.3 0.00086896 0 0.00086888 0 0.00086898 3.3 0.0008689 3.3 0.000869 0 0.00086892 0 0.00086902 3.3 0.00086894 3.3 0.00086904 0 0.00086896 0 0.00086906 3.3 0.00086898 3.3 0.0008690799999999999 0 0.000869 0 0.0008690999999999999 3.3 0.0008690200000000001 3.3 0.00086912 0 0.0008690400000000001 0 0.00086914 3.3 0.0008690600000000001 3.3 0.00086916 0 0.00086908 0 0.00086918 3.3 0.0008691 3.3 0.0008692 0 0.00086912 0 0.00086922 3.3 0.00086914 3.3 0.00086924 0 0.00086916 0 0.00086926 3.3 0.00086918 3.3 0.0008692799999999999 0 0.0008692 0 0.0008692999999999999 3.3 0.0008692200000000001 3.3 0.00086932 0 0.0008692400000000001 0 0.00086934 3.3 0.0008692600000000001 3.3 0.00086936 0 0.00086928 0 0.00086938 3.3 0.0008693 3.3 0.0008694 0 0.00086932 0 0.00086942 3.3 0.00086934 3.3 0.00086944 0 0.00086936 0 0.00086946 3.3 0.00086938 3.3 0.00086948 0 0.0008694 0 0.0008694999999999999 3.3 0.00086942 3.3 0.0008695199999999999 0 0.0008694400000000001 0 0.00086954 3.3 0.0008694600000000001 3.3 0.00086956 0 0.0008694800000000001 0 0.00086958 3.3 0.0008695 3.3 0.0008696 0 0.00086952 0 0.00086962 3.3 0.00086954 3.3 0.00086964 0 0.00086956 0 0.00086966 3.3 0.00086958 3.3 0.00086968 0 0.0008696 0 0.0008696999999999999 3.3 0.00086962 3.3 0.0008697199999999999 0 0.0008696400000000001 0 0.00086974 3.3 0.0008696600000000001 3.3 0.00086976 0 0.0008696800000000001 0 0.00086978 3.3 0.0008697 3.3 0.0008698 0 0.00086972 0 0.00086982 3.3 0.00086974 3.3 0.00086984 0 0.00086976 0 0.00086986 3.3 0.00086978 3.3 0.00086988 0 0.0008698 0 0.0008699 3.3 0.00086982 3.3 0.0008699199999999999 0 0.0008698400000000001 0 0.00086994 3.3 0.0008698600000000001 3.3 0.00086996 0 0.0008698800000000001 0 0.00086998 3.3 0.0008699000000000001 3.3 0.00087 0 0.00086992 0 0.00087002 3.3 0.00086994 3.3 0.00087004 0 0.00086996 0 0.00087006 3.3 0.00086998 3.3 0.00087008 0 0.00087 0 0.0008701 3.3 0.00087002 3.3 0.0008701199999999999 0 0.00087004 0 0.0008701399999999999 3.3 0.0008700600000000001 3.3 0.00087016 0 0.0008700800000000001 0 0.00087018 3.3 0.0008701000000000001 3.3 0.0008702 0 0.00087012 0 0.00087022 3.3 0.00087014 3.3 0.00087024 0 0.00087016 0 0.00087026 3.3 0.00087018 3.3 0.00087028 0 0.0008702 0 0.0008703 3.3 0.00087022 3.3 0.00087032 0 0.00087024 0 0.0008703399999999999 3.3 0.0008702600000000001 3.3 0.00087036 0 0.0008702800000000001 0 0.00087038 3.3 0.0008703000000000001 3.3 0.0008704 0 0.0008703200000000001 0 0.00087042 3.3 0.00087034 3.3 0.00087044 0 0.00087036 0 0.00087046 3.3 0.00087038 3.3 0.00087048 0 0.0008704 0 0.0008705 3.3 0.00087042 3.3 0.00087052 0 0.00087044 0 0.0008705399999999999 3.3 0.00087046 3.3 0.0008705599999999999 0 0.0008704800000000001 0 0.00087058 3.3 0.0008705000000000001 3.3 0.0008706 0 0.0008705200000000001 0 0.00087062 3.3 0.00087054 3.3 0.00087064 0 0.00087056 0 0.00087066 3.3 0.00087058 3.3 0.00087068 0 0.0008706 0 0.0008707 3.3 0.00087062 3.3 0.00087072 0 0.00087064 0 0.00087074 3.3 0.00087066 3.3 0.0008707599999999999 0 0.0008706800000000001 0 0.00087078 3.3 0.0008707000000000001 3.3 0.0008708 0 0.0008707200000000001 0 0.00087082 3.3 0.0008707400000000001 3.3 0.00087084 0 0.00087076 0 0.00087086 3.3 0.00087078 3.3 0.00087088 0 0.0008708 0 0.0008709 3.3 0.00087082 3.3 0.00087092 0 0.00087084 0 0.00087094 3.3 0.00087086 3.3 0.0008709599999999999 0 0.00087088 0 0.0008709799999999999 3.3 0.0008709000000000001 3.3 0.000871 0 0.0008709200000000001 0 0.00087102 3.3 0.0008709400000000001 3.3 0.00087104 0 0.00087096 0 0.00087106 3.3 0.00087098 3.3 0.00087108 0 0.000871 0 0.0008711 3.3 0.00087102 3.3 0.00087112 0 0.00087104 0 0.00087114 3.3 0.00087106 3.3 0.00087116 0 0.00087108 0 0.0008711799999999999 3.3 0.0008711000000000001 3.3 0.0008712 0 0.0008711200000000001 0 0.00087122 3.3 0.0008711400000000001 3.3 0.00087124 0 0.0008711600000000001 0 0.00087126 3.3 0.00087118 3.3 0.00087128 0 0.0008712 0 0.0008713 3.3 0.00087122 3.3 0.00087132 0 0.00087124 0 0.00087134 3.3 0.00087126 3.3 0.00087136 0 0.00087128 0 0.0008713799999999999 3.3 0.0008713 3.3 0.0008713999999999999 0 0.0008713200000000001 0 0.00087142 3.3 0.0008713400000000001 3.3 0.00087144 0 0.0008713600000000001 0 0.00087146 3.3 0.00087138 3.3 0.00087148 0 0.0008714 0 0.0008715 3.3 0.00087142 3.3 0.00087152 0 0.00087144 0 0.00087154 3.3 0.00087146 3.3 0.00087156 0 0.00087148 0 0.00087158 3.3 0.0008715 3.3 0.0008715999999999999 0 0.0008715200000000001 0 0.00087162 3.3 0.0008715400000000001 3.3 0.00087164 0 0.0008715600000000001 0 0.00087166 3.3 0.0008715800000000001 3.3 0.00087168 0 0.0008716 0 0.0008717 3.3 0.00087162 3.3 0.00087172 0 0.00087164 0 0.00087174 3.3 0.00087166 3.3 0.00087176 0 0.00087168 0 0.00087178 3.3 0.0008717 3.3 0.0008717999999999999 0 0.00087172 0 0.0008718199999999999 3.3 0.0008717400000000001 3.3 0.00087184 0 0.0008717600000000001 0 0.00087186 3.3 0.0008717800000000001 3.3 0.00087188 0 0.0008718 0 0.0008719 3.3 0.00087182 3.3 0.00087192 0 0.00087184 0 0.00087194 3.3 0.00087186 3.3 0.00087196 0 0.00087188 0 0.00087198 3.3 0.0008719 3.3 0.0008719999999999999 0 0.00087192 0 0.0008720199999999999 3.3 0.0008719400000000001 3.3 0.00087204 0 0.0008719600000000001 0 0.00087206 3.3 0.0008719800000000001 3.3 0.00087208 0 0.000872 0 0.0008721 3.3 0.00087202 3.3 0.00087212 0 0.00087204 0 0.00087214 3.3 0.00087206 3.3 0.00087216 0 0.00087208 0 0.00087218 3.3 0.0008721 3.3 0.0008722 0 0.00087212 0 0.0008722199999999999 3.3 0.00087214 3.3 0.0008722399999999999 0 0.0008721600000000001 0 0.00087226 3.3 0.0008721800000000001 3.3 0.00087228 0 0.0008722000000000001 0 0.0008723 3.3 0.00087222 3.3 0.00087232 0 0.00087224 0 0.00087234 3.3 0.00087226 3.3 0.00087236 0 0.00087228 0 0.00087238 3.3 0.0008723 3.3 0.0008724 0 0.00087232 0 0.0008724199999999999 3.3 0.00087234 3.3 0.0008724399999999999 0 0.0008723600000000001 0 0.00087246 3.3 0.0008723800000000001 3.3 0.00087248 0 0.0008724000000000001 0 0.0008725 3.3 0.00087242 3.3 0.00087252 0 0.00087244 0 0.00087254 3.3 0.00087246 3.3 0.00087256 0 0.00087248 0 0.00087258 3.3 0.0008725 3.3 0.0008726 0 0.00087252 0 0.00087262 3.3 0.00087254 3.3 0.0008726399999999999 0 0.00087256 0 0.0008726599999999999 3.3 0.0008725800000000001 3.3 0.00087268 0 0.0008726000000000001 0 0.0008727 3.3 0.0008726200000000001 3.3 0.00087272 0 0.00087264 0 0.00087274 3.3 0.00087266 3.3 0.00087276 0 0.00087268 0 0.00087278 3.3 0.0008727 3.3 0.0008728 0 0.00087272 0 0.00087282 3.3 0.00087274 3.3 0.0008728399999999999 0 0.00087276 0 0.0008728599999999999 3.3 0.0008727800000000001 3.3 0.00087288 0 0.0008728000000000001 0 0.0008729 3.3 0.0008728200000000001 3.3 0.00087292 0 0.00087284 0 0.00087294 3.3 0.00087286 3.3 0.00087296 0 0.00087288 0 0.00087298 3.3 0.0008729 3.3 0.000873 0 0.00087292 0 0.00087302 3.3 0.00087294 3.3 0.00087304 0 0.00087296 0 0.0008730599999999999 3.3 0.0008729800000000001 3.3 0.00087308 0 0.0008730000000000001 0 0.0008731 3.3 0.0008730200000000001 3.3 0.00087312 0 0.0008730400000000001 0 0.00087314 3.3 0.00087306 3.3 0.00087316 0 0.00087308 0 0.00087318 3.3 0.0008731 3.3 0.0008732 0 0.00087312 0 0.00087322 3.3 0.00087314 3.3 0.00087324 0 0.00087316 0 0.0008732599999999999 3.3 0.00087318 3.3 0.0008732799999999999 0 0.0008732000000000001 0 0.0008733 3.3 0.0008732200000000001 3.3 0.00087332 0 0.0008732400000000001 0 0.00087334 3.3 0.00087326 3.3 0.00087336 0 0.00087328 0 0.00087338 3.3 0.0008733 3.3 0.0008734 0 0.00087332 0 0.00087342 3.3 0.00087334 3.3 0.00087344 0 0.00087336 0 0.00087346 3.3 0.00087338 3.3 0.0008734799999999999 0 0.0008734000000000001 0 0.0008735 3.3 0.0008734200000000001 3.3 0.00087352 0 0.0008734400000000001 0 0.00087354 3.3 0.0008734600000000001 3.3 0.00087356 0 0.00087348 0 0.00087358 3.3 0.0008735 3.3 0.0008736 0 0.00087352 0 0.00087362 3.3 0.00087354 3.3 0.00087364 0 0.00087356 0 0.00087366 3.3 0.00087358 3.3 0.0008736799999999999 0 0.0008736 0 0.0008736999999999999 3.3 0.0008736200000000001 3.3 0.00087372 0 0.0008736400000000001 0 0.00087374 3.3 0.0008736600000000001 3.3 0.00087376 0 0.00087368 0 0.00087378 3.3 0.0008737 3.3 0.0008738 0 0.00087372 0 0.00087382 3.3 0.00087374 3.3 0.00087384 0 0.00087376 0 0.00087386 3.3 0.00087378 3.3 0.00087388 0 0.0008738 0 0.0008738999999999999 3.3 0.0008738200000000001 3.3 0.00087392 0 0.0008738400000000001 0 0.00087394 3.3 0.0008738600000000001 3.3 0.00087396 0 0.0008738800000000001 0 0.00087398 3.3 0.0008739 3.3 0.000874 0 0.00087392 0 0.00087402 3.3 0.00087394 3.3 0.00087404 0 0.00087396 0 0.00087406 3.3 0.00087398 3.3 0.00087408 0 0.000874 0 0.0008740999999999999 3.3 0.00087402 3.3 0.0008741199999999999 0 0.0008740400000000001 0 0.00087414 3.3 0.0008740600000000001 3.3 0.00087416 0 0.0008740800000000001 0 0.00087418 3.3 0.0008741 3.3 0.0008742 0 0.00087412 0 0.00087422 3.3 0.00087414 3.3 0.00087424 0 0.00087416 0 0.00087426 3.3 0.00087418 3.3 0.00087428 0 0.0008742 0 0.0008743 3.3 0.00087422 3.3 0.0008743199999999999 0 0.0008742400000000001 0 0.00087434 3.3 0.0008742600000000001 3.3 0.00087436 0 0.0008742800000000001 0 0.00087438 3.3 0.0008743000000000001 3.3 0.0008744 0 0.00087432 0 0.00087442 3.3 0.00087434 3.3 0.00087444 0 0.00087436 0 0.00087446 3.3 0.00087438 3.3 0.00087448 0 0.0008744 0 0.0008745 3.3 0.00087442 3.3 0.0008745199999999999 0 0.00087444 0 0.0008745399999999999 3.3 0.0008744600000000001 3.3 0.00087456 0 0.0008744800000000001 0 0.00087458 3.3 0.0008745000000000001 3.3 0.0008746 0 0.00087452 0 0.00087462 3.3 0.00087454 3.3 0.00087464 0 0.00087456 0 0.00087466 3.3 0.00087458 3.3 0.00087468 0 0.0008746 0 0.0008747 3.3 0.00087462 3.3 0.00087472 0 0.00087464 0 0.0008747399999999999 3.3 0.0008746600000000001 3.3 0.00087476 0 0.0008746800000000001 0 0.00087478 3.3 0.0008747000000000001 3.3 0.0008748 0 0.0008747200000000001 0 0.00087482 3.3 0.00087474 3.3 0.00087484 0 0.00087476 0 0.00087486 3.3 0.00087478 3.3 0.00087488 0 0.0008748 0 0.0008749 3.3 0.00087482 3.3 0.00087492 0 0.00087484 0 0.0008749399999999999 3.3 0.00087486 3.3 0.0008749599999999999 0 0.0008748800000000001 0 0.00087498 3.3 0.0008749000000000001 3.3 0.000875 0 0.0008749200000000001 0 0.00087502 3.3 0.00087494 3.3 0.00087504 0 0.00087496 0 0.00087506 3.3 0.00087498 3.3 0.00087508 0 0.000875 0 0.0008751 3.3 0.00087502 3.3 0.00087512 0 0.00087504 0 0.0008751399999999999 3.3 0.00087506 3.3 0.0008751599999999999 0 0.0008750800000000001 0 0.00087518 3.3 0.0008751000000000001 3.3 0.0008752 0 0.0008751200000000001 0 0.00087522 3.3 0.00087514 3.3 0.00087524 0 0.00087516 0 0.00087526 3.3 0.00087518 3.3 0.00087528 0 0.0008752 0 0.0008753 3.3 0.00087522 3.3 0.00087532 0 0.00087524 0 0.00087534 3.3 0.00087526 3.3 0.0008753599999999999 0 0.00087528 0 0.0008753799999999999 3.3 0.0008753000000000001 3.3 0.0008754 0 0.0008753200000000001 0 0.00087542 3.3 0.0008753400000000001 3.3 0.00087544 0 0.00087536 0 0.00087546 3.3 0.00087538 3.3 0.00087548 0 0.0008754 0 0.0008755 3.3 0.00087542 3.3 0.00087552 0 0.00087544 0 0.00087554 3.3 0.00087546 3.3 0.0008755599999999999 0 0.00087548 0 0.0008755799999999999 3.3 0.0008755000000000001 3.3 0.0008756 0 0.0008755200000000001 0 0.00087562 3.3 0.0008755400000000001 3.3 0.00087564 0 0.00087556 0 0.00087566 3.3 0.00087558 3.3 0.00087568 0 0.0008756 0 0.0008757 3.3 0.00087562 3.3 0.00087572 0 0.00087564 0 0.00087574 3.3 0.00087566 3.3 0.00087576 0 0.00087568 0 0.0008757799999999999 3.3 0.0008757 3.3 0.0008757999999999999 0 0.0008757200000000001 0 0.00087582 3.3 0.0008757400000000001 3.3 0.00087584 0 0.0008757600000000001 0 0.00087586 3.3 0.00087578 3.3 0.00087588 0 0.0008758 0 0.0008759 3.3 0.00087582 3.3 0.00087592 0 0.00087584 0 0.00087594 3.3 0.00087586 3.3 0.00087596 0 0.00087588 0 0.0008759799999999999 3.3 0.0008759 3.3 0.0008759999999999999 0 0.0008759200000000001 0 0.00087602 3.3 0.0008759400000000001 3.3 0.00087604 0 0.0008759600000000001 0 0.00087606 3.3 0.00087598 3.3 0.00087608 0 0.000876 0 0.0008761 3.3 0.00087602 3.3 0.00087612 0 0.00087604 0 0.00087614 3.3 0.00087606 3.3 0.00087616 0 0.00087608 0 0.00087618 3.3 0.0008761 3.3 0.0008761999999999999 0 0.00087612 0 0.0008762199999999999 3.3 0.0008761400000000001 3.3 0.00087624 0 0.0008761600000000001 0 0.00087626 3.3 0.0008761800000000001 3.3 0.00087628 0 0.0008762 0 0.0008763 3.3 0.00087622 3.3 0.00087632 0 0.00087624 0 0.00087634 3.3 0.00087626 3.3 0.00087636 0 0.00087628 0 0.00087638 3.3 0.0008763 3.3 0.0008763999999999999 0 0.00087632 0 0.0008764199999999999 3.3 0.0008763400000000001 3.3 0.00087644 0 0.0008763600000000001 0 0.00087646 3.3 0.0008763800000000001 3.3 0.00087648 0 0.0008764 0 0.0008765 3.3 0.00087642 3.3 0.00087652 0 0.00087644 0 0.00087654 3.3 0.00087646 3.3 0.00087656 0 0.00087648 0 0.00087658 3.3 0.0008765 3.3 0.0008766 0 0.00087652 0 0.0008766199999999999 3.3 0.0008765400000000001 3.3 0.00087664 0 0.0008765600000000001 0 0.00087666 3.3 0.0008765800000000001 3.3 0.00087668 0 0.0008766000000000001 0 0.0008767 3.3 0.00087662 3.3 0.00087672 0 0.00087664 0 0.00087674 3.3 0.00087666 3.3 0.00087676 0 0.00087668 0 0.00087678 3.3 0.0008767 3.3 0.0008768 0 0.00087672 0 0.0008768199999999999 3.3 0.00087674 3.3 0.0008768399999999999 0 0.0008767600000000001 0 0.00087686 3.3 0.0008767800000000001 3.3 0.00087688 0 0.0008768000000000001 0 0.0008769 3.3 0.00087682 3.3 0.00087692 0 0.00087684 0 0.00087694 3.3 0.00087686 3.3 0.00087696 0 0.00087688 0 0.00087698 3.3 0.0008769 3.3 0.000877 0 0.00087692 0 0.00087702 3.3 0.00087694 3.3 0.0008770399999999999 0 0.0008769600000000001 0 0.00087706 3.3 0.0008769800000000001 3.3 0.00087708 0 0.0008770000000000001 0 0.0008771 3.3 0.0008770200000000001 3.3 0.00087712 0 0.00087704 0 0.00087714 3.3 0.00087706 3.3 0.00087716 0 0.00087708 0 0.00087718 3.3 0.0008771 3.3 0.0008772 0 0.00087712 0 0.00087722 3.3 0.00087714 3.3 0.0008772399999999999 0 0.00087716 0 0.0008772599999999999 3.3 0.0008771800000000001 3.3 0.00087728 0 0.0008772000000000001 0 0.0008773 3.3 0.0008772200000000001 3.3 0.00087732 0 0.00087724 0 0.00087734 3.3 0.00087726 3.3 0.00087736 0 0.00087728 0 0.00087738 3.3 0.0008773 3.3 0.0008774 0 0.00087732 0 0.00087742 3.3 0.00087734 3.3 0.00087744 0 0.00087736 0 0.0008774599999999999 3.3 0.0008773800000000001 3.3 0.00087748 0 0.0008774000000000001 0 0.0008775 3.3 0.0008774200000000001 3.3 0.00087752 0 0.0008774400000000001 0 0.00087754 3.3 0.00087746 3.3 0.00087756 0 0.00087748 0 0.00087758 3.3 0.0008775 3.3 0.0008776 0 0.00087752 0 0.00087762 3.3 0.00087754 3.3 0.00087764 0 0.00087756 0 0.0008776599999999999 3.3 0.00087758 3.3 0.0008776799999999999 0 0.0008776000000000001 0 0.0008777 3.3 0.0008776200000000001 3.3 0.00087772 0 0.0008776400000000001 0 0.00087774 3.3 0.00087766 3.3 0.00087776 0 0.00087768 0 0.00087778 3.3 0.0008777 3.3 0.0008778 0 0.00087772 0 0.00087782 3.3 0.00087774 3.3 0.00087784 0 0.00087776 0 0.00087786 3.3 0.00087778 3.3 0.0008778799999999999 0 0.0008778000000000001 0 0.0008779 3.3 0.0008778200000000001 3.3 0.00087792 0 0.0008778400000000001 0 0.00087794 3.3 0.0008778600000000001 3.3 0.00087796 0 0.00087788 0 0.00087798 3.3 0.0008779 3.3 0.000878 0 0.00087792 0 0.00087802 3.3 0.00087794 3.3 0.00087804 0 0.00087796 0 0.00087806 3.3 0.00087798 3.3 0.0008780799999999999 0 0.000878 0 0.0008780999999999999 3.3 0.0008780200000000001 3.3 0.00087812 0 0.0008780400000000001 0 0.00087814 3.3 0.0008780600000000001 3.3 0.00087816 0 0.00087808 0 0.00087818 3.3 0.0008781 3.3 0.0008782 0 0.00087812 0 0.00087822 3.3 0.00087814 3.3 0.00087824 0 0.00087816 0 0.00087826 3.3 0.00087818 3.3 0.00087828 0 0.0008782 0 0.0008782999999999999 3.3 0.0008782200000000001 3.3 0.00087832 0 0.0008782400000000001 0 0.00087834 3.3 0.0008782600000000001 3.3 0.00087836 0 0.0008782800000000001 0 0.00087838 3.3 0.0008783 3.3 0.0008784 0 0.00087832 0 0.00087842 3.3 0.00087834 3.3 0.00087844 0 0.00087836 0 0.00087846 3.3 0.00087838 3.3 0.00087848 0 0.0008784 0 0.0008784999999999999 3.3 0.00087842 3.3 0.0008785199999999999 0 0.0008784400000000001 0 0.00087854 3.3 0.0008784600000000001 3.3 0.00087856 0 0.0008784800000000001 0 0.00087858 3.3 0.0008785 3.3 0.0008786 0 0.00087852 0 0.00087862 3.3 0.00087854 3.3 0.00087864 0 0.00087856 0 0.00087866 3.3 0.00087858 3.3 0.00087868 0 0.0008786 0 0.0008786999999999999 3.3 0.00087862 3.3 0.0008787199999999999 0 0.0008786400000000001 0 0.00087874 3.3 0.0008786600000000001 3.3 0.00087876 0 0.0008786800000000001 0 0.00087878 3.3 0.0008787 3.3 0.0008788 0 0.00087872 0 0.00087882 3.3 0.00087874 3.3 0.00087884 0 0.00087876 0 0.00087886 3.3 0.00087878 3.3 0.00087888 0 0.0008788 0 0.0008789 3.3 0.00087882 3.3 0.0008789199999999999 0 0.00087884 0 0.0008789399999999999 3.3 0.0008788600000000001 3.3 0.00087896 0 0.0008788800000000001 0 0.00087898 3.3 0.0008789000000000001 3.3 0.000879 0 0.00087892 0 0.00087902 3.3 0.00087894 3.3 0.00087904 0 0.00087896 0 0.00087906 3.3 0.00087898 3.3 0.00087908 0 0.000879 0 0.0008791 3.3 0.00087902 3.3 0.0008791199999999999 0 0.00087904 0 0.0008791399999999999 3.3 0.0008790600000000001 3.3 0.00087916 0 0.0008790800000000001 0 0.00087918 3.3 0.0008791000000000001 3.3 0.0008792 0 0.00087912 0 0.00087922 3.3 0.00087914 3.3 0.00087924 0 0.00087916 0 0.00087926 3.3 0.00087918 3.3 0.00087928 0 0.0008792 0 0.0008793 3.3 0.00087922 3.3 0.00087932 0 0.00087924 0 0.0008793399999999999 3.3 0.00087926 3.3 0.0008793599999999999 0 0.0008792800000000001 0 0.00087938 3.3 0.0008793000000000001 3.3 0.0008794 0 0.0008793200000000001 0 0.00087942 3.3 0.00087934 3.3 0.00087944 0 0.00087936 0 0.00087946 3.3 0.00087938 3.3 0.00087948 0 0.0008794 0 0.0008795 3.3 0.00087942 3.3 0.00087952 0 0.00087944 0 0.0008795399999999999 3.3 0.00087946 3.3 0.0008795599999999999 0 0.0008794800000000001 0 0.00087958 3.3 0.0008795000000000001 3.3 0.0008796 0 0.0008795200000000001 0 0.00087962 3.3 0.00087954 3.3 0.00087964 0 0.00087956 0 0.00087966 3.3 0.00087958 3.3 0.00087968 0 0.0008796 0 0.0008797 3.3 0.00087962 3.3 0.00087972 0 0.00087964 0 0.00087974 3.3 0.00087966 3.3 0.0008797599999999999 0 0.00087968 0 0.0008797799999999999 3.3 0.0008797000000000001 3.3 0.0008798 0 0.0008797200000000001 0 0.00087982 3.3 0.0008797400000000001 3.3 0.00087984 0 0.00087976 0 0.00087986 3.3 0.00087978 3.3 0.00087988 0 0.0008798 0 0.0008799 3.3 0.00087982 3.3 0.00087992 0 0.00087984 0 0.00087994 3.3 0.00087986 3.3 0.0008799599999999999 0 0.00087988 0 0.0008799799999999999 3.3 0.0008799000000000001 3.3 0.00088 0 0.0008799200000000001 0 0.00088002 3.3 0.0008799400000000001 3.3 0.00088004 0 0.00087996 0 0.00088006 3.3 0.00087998 3.3 0.00088008 0 0.00088 0 0.0008801 3.3 0.00088002 3.3 0.00088012 0 0.00088004 0 0.00088014 3.3 0.00088006 3.3 0.00088016 0 0.00088008 0 0.0008801799999999999 3.3 0.0008801000000000001 3.3 0.0008802 0 0.0008801200000000001 0 0.00088022 3.3 0.0008801400000000001 3.3 0.00088024 0 0.0008801600000000001 0 0.00088026 3.3 0.00088018 3.3 0.00088028 0 0.0008802 0 0.0008803 3.3 0.00088022 3.3 0.00088032 0 0.00088024 0 0.00088034 3.3 0.00088026 3.3 0.00088036 0 0.00088028 0 0.0008803799999999999 3.3 0.0008803 3.3 0.0008803999999999999 0 0.0008803200000000001 0 0.00088042 3.3 0.0008803400000000001 3.3 0.00088044 0 0.0008803600000000001 0 0.00088046 3.3 0.00088038 3.3 0.00088048 0 0.0008804 0 0.0008805 3.3 0.00088042 3.3 0.00088052 0 0.00088044 0 0.00088054 3.3 0.00088046 3.3 0.00088056 0 0.00088048 0 0.00088058 3.3 0.0008805 3.3 0.0008805999999999999 0 0.0008805200000000001 0 0.00088062 3.3 0.0008805400000000001 3.3 0.00088064 0 0.0008805600000000001 0 0.00088066 3.3 0.0008805800000000001 3.3 0.00088068 0 0.0008806 0 0.0008807 3.3 0.00088062 3.3 0.00088072 0 0.00088064 0 0.00088074 3.3 0.00088066 3.3 0.00088076 0 0.00088068 0 0.00088078 3.3 0.0008807 3.3 0.0008807999999999999 0 0.00088072 0 0.0008808199999999999 3.3 0.0008807400000000001 3.3 0.00088084 0 0.0008807600000000001 0 0.00088086 3.3 0.0008807800000000001 3.3 0.00088088 0 0.0008808 0 0.0008809 3.3 0.00088082 3.3 0.00088092 0 0.00088084 0 0.00088094 3.3 0.00088086 3.3 0.00088096 0 0.00088088 0 0.00088098 3.3 0.0008809 3.3 0.000881 0 0.00088092 0 0.0008810199999999999 3.3 0.0008809400000000001 3.3 0.00088104 0 0.0008809600000000001 0 0.00088106 3.3 0.0008809800000000001 3.3 0.00088108 0 0.0008810000000000001 0 0.0008811 3.3 0.00088102 3.3 0.00088112 0 0.00088104 0 0.00088114 3.3 0.00088106 3.3 0.00088116 0 0.00088108 0 0.00088118 3.3 0.0008811 3.3 0.0008812 0 0.00088112 0 0.0008812199999999999 3.3 0.00088114 3.3 0.0008812399999999999 0 0.0008811600000000001 0 0.00088126 3.3 0.0008811800000000001 3.3 0.00088128 0 0.0008812000000000001 0 0.0008813 3.3 0.00088122 3.3 0.00088132 0 0.00088124 0 0.00088134 3.3 0.00088126 3.3 0.00088136 0 0.00088128 0 0.00088138 3.3 0.0008813 3.3 0.0008814 0 0.00088132 0 0.00088142 3.3 0.00088134 3.3 0.0008814399999999999 0 0.0008813600000000001 0 0.00088146 3.3 0.0008813800000000001 3.3 0.00088148 0 0.0008814000000000001 0 0.0008815 3.3 0.0008814200000000001 3.3 0.00088152 0 0.00088144 0 0.00088154 3.3 0.00088146 3.3 0.00088156 0 0.00088148 0 0.00088158 3.3 0.0008815 3.3 0.0008816 0 0.00088152 0 0.00088162 3.3 0.00088154 3.3 0.0008816399999999999 0 0.00088156 0 0.0008816599999999999 3.3 0.0008815800000000001 3.3 0.00088168 0 0.0008816000000000001 0 0.0008817 3.3 0.0008816200000000001 3.3 0.00088172 0 0.00088164 0 0.00088174 3.3 0.00088166 3.3 0.00088176 0 0.00088168 0 0.00088178 3.3 0.0008817 3.3 0.0008818 0 0.00088172 0 0.00088182 3.3 0.00088174 3.3 0.00088184 0 0.00088176 0 0.0008818599999999999 3.3 0.0008817800000000001 3.3 0.00088188 0 0.0008818000000000001 0 0.0008819 3.3 0.0008818200000000001 3.3 0.00088192 0 0.0008818400000000001 0 0.00088194 3.3 0.00088186 3.3 0.00088196 0 0.00088188 0 0.00088198 3.3 0.0008819 3.3 0.000882 0 0.00088192 0 0.00088202 3.3 0.00088194 3.3 0.00088204 0 0.00088196 0 0.0008820599999999999 3.3 0.00088198 3.3 0.0008820799999999999 0 0.0008820000000000001 0 0.0008821 3.3 0.0008820200000000001 3.3 0.00088212 0 0.0008820400000000001 0 0.00088214 3.3 0.00088206 3.3 0.00088216 0 0.00088208 0 0.00088218 3.3 0.0008821 3.3 0.0008822 0 0.00088212 0 0.00088222 3.3 0.00088214 3.3 0.00088224 0 0.00088216 0 0.0008822599999999999 3.3 0.00088218 3.3 0.0008822799999999999 0 0.0008822000000000001 0 0.0008823 3.3 0.0008822200000000001 3.3 0.00088232 0 0.0008822400000000001 0 0.00088234 3.3 0.00088226 3.3 0.00088236 0 0.00088228 0 0.00088238 3.3 0.0008823 3.3 0.0008824 0 0.00088232 0 0.00088242 3.3 0.00088234 3.3 0.00088244 0 0.00088236 0 0.00088246 3.3 0.00088238 3.3 0.0008824799999999999 0 0.0008824 0 0.0008824999999999999 3.3 0.0008824200000000001 3.3 0.00088252 0 0.0008824400000000001 0 0.00088254 3.3 0.0008824600000000001 3.3 0.00088256 0 0.00088248 0 0.00088258 3.3 0.0008825 3.3 0.0008826 0 0.00088252 0 0.00088262 3.3 0.00088254 3.3 0.00088264 0 0.00088256 0 0.00088266 3.3 0.00088258 3.3 0.0008826799999999999 0 0.0008826 0 0.0008826999999999999 3.3 0.0008826200000000001 3.3 0.00088272 0 0.0008826400000000001 0 0.00088274 3.3 0.0008826600000000001 3.3 0.00088276 0 0.00088268 0 0.00088278 3.3 0.0008827 3.3 0.0008828 0 0.00088272 0 0.00088282 3.3 0.00088274 3.3 0.00088284 0 0.00088276 0 0.00088286 3.3 0.00088278 3.3 0.00088288 0 0.0008828 0 0.0008828999999999999 3.3 0.00088282 3.3 0.0008829199999999999 0 0.0008828400000000001 0 0.00088294 3.3 0.0008828600000000001 3.3 0.00088296 0 0.0008828800000000001 0 0.00088298 3.3 0.0008829 3.3 0.000883 0 0.00088292 0 0.00088302 3.3 0.00088294 3.3 0.00088304 0 0.00088296 0 0.00088306 3.3 0.00088298 3.3 0.00088308 0 0.000883 0 0.0008830999999999999 3.3 0.00088302 3.3 0.0008831199999999999 0 0.0008830400000000001 0 0.00088314 3.3 0.0008830600000000001 3.3 0.00088316 0 0.0008830800000000001 0 0.00088318 3.3 0.0008831 3.3 0.0008832 0 0.00088312 0 0.00088322 3.3 0.00088314 3.3 0.00088324 0 0.00088316 0 0.00088326 3.3 0.00088318 3.3 0.00088328 0 0.0008832 0 0.0008833 3.3 0.00088322 3.3 0.0008833199999999999 0 0.00088324 0 0.0008833399999999999 3.3 0.0008832600000000001 3.3 0.00088336 0 0.0008832800000000001 0 0.00088338 3.3 0.0008833000000000001 3.3 0.0008834 0 0.00088332 0 0.00088342 3.3 0.00088334 3.3 0.00088344 0 0.00088336 0 0.00088346 3.3 0.00088338 3.3 0.00088348 0 0.0008834 0 0.0008835 3.3 0.00088342 3.3 0.0008835199999999999 0 0.00088344 0 0.0008835399999999999 3.3 0.0008834600000000001 3.3 0.00088356 0 0.0008834800000000001 0 0.00088358 3.3 0.0008835000000000001 3.3 0.0008836 0 0.00088352 0 0.00088362 3.3 0.00088354 3.3 0.00088364 0 0.00088356 0 0.00088366 3.3 0.00088358 3.3 0.00088368 0 0.0008836 0 0.0008837 3.3 0.00088362 3.3 0.00088372 0 0.00088364 0 0.0008837399999999999 3.3 0.0008836600000000001 3.3 0.00088376 0 0.0008836800000000001 0 0.00088378 3.3 0.0008837000000000001 3.3 0.0008838 0 0.0008837200000000001 0 0.00088382 3.3 0.00088374 3.3 0.00088384 0 0.00088376 0 0.00088386 3.3 0.00088378 3.3 0.00088388 0 0.0008838 0 0.0008839 3.3 0.00088382 3.3 0.00088392 0 0.00088384 0 0.0008839399999999999 3.3 0.00088386 3.3 0.0008839599999999999 0 0.0008838800000000001 0 0.00088398 3.3 0.0008839000000000001 3.3 0.000884 0 0.0008839200000000001 0 0.00088402 3.3 0.00088394 3.3 0.00088404 0 0.00088396 0 0.00088406 3.3 0.00088398 3.3 0.00088408 0 0.000884 0 0.0008841 3.3 0.00088402 3.3 0.00088412 0 0.00088404 0 0.00088414 3.3 0.00088406 3.3 0.0008841599999999999 0 0.0008840800000000001 0 0.00088418 3.3 0.0008841000000000001 3.3 0.0008842 0 0.0008841200000000001 0 0.00088422 3.3 0.0008841400000000001 3.3 0.00088424 0 0.00088416 0 0.00088426 3.3 0.00088418 3.3 0.00088428 0 0.0008842 0 0.0008843 3.3 0.00088422 3.3 0.00088432 0 0.00088424 0 0.00088434 3.3 0.00088426 3.3 0.0008843599999999999 0 0.00088428 0 0.0008843799999999999 3.3 0.0008843000000000001 3.3 0.0008844 0 0.0008843200000000001 0 0.00088442 3.3 0.0008843400000000001 3.3 0.00088444 0 0.00088436 0 0.00088446 3.3 0.00088438 3.3 0.00088448 0 0.0008844 0 0.0008845 3.3 0.00088442 3.3 0.00088452 0 0.00088444 0 0.00088454 3.3 0.00088446 3.3 0.00088456 0 0.00088448 0 0.0008845799999999999 3.3 0.0008845000000000001 3.3 0.0008846 0 0.0008845200000000001 0 0.00088462 3.3 0.0008845400000000001 3.3 0.00088464 0 0.0008845600000000001 0 0.00088466 3.3 0.00088458 3.3 0.00088468 0 0.0008846 0 0.0008847 3.3 0.00088462 3.3 0.00088472 0 0.00088464 0 0.00088474 3.3 0.00088466 3.3 0.00088476 0 0.00088468 0 0.0008847799999999999 3.3 0.0008847 3.3 0.0008847999999999999 0 0.0008847200000000001 0 0.00088482 3.3 0.0008847400000000001 3.3 0.00088484 0 0.0008847600000000001 0 0.00088486 3.3 0.00088478 3.3 0.00088488 0 0.0008848 0 0.0008849 3.3 0.00088482 3.3 0.00088492 0 0.00088484 0 0.00088494 3.3 0.00088486 3.3 0.00088496 0 0.00088488 0 0.00088498 3.3 0.0008849 3.3 0.0008849999999999999 0 0.0008849200000000001 0 0.00088502 3.3 0.0008849400000000001 3.3 0.00088504 0 0.0008849600000000001 0 0.00088506 3.3 0.0008849800000000001 3.3 0.00088508 0 0.000885 0 0.0008851 3.3 0.00088502 3.3 0.00088512 0 0.00088504 0 0.00088514 3.3 0.00088506 3.3 0.00088516 0 0.00088508 0 0.00088518 3.3 0.0008851 3.3 0.0008851999999999999 0 0.00088512 0 0.0008852199999999999 3.3 0.0008851400000000001 3.3 0.00088524 0 0.0008851600000000001 0 0.00088526 3.3 0.0008851800000000001 3.3 0.00088528 0 0.0008852 0 0.0008853 3.3 0.00088522 3.3 0.00088532 0 0.00088524 0 0.00088534 3.3 0.00088526 3.3 0.00088536 0 0.00088528 0 0.00088538 3.3 0.0008853 3.3 0.0008853999999999999 0 0.00088532 0 0.0008854199999999999 3.3 0.0008853400000000001 3.3 0.00088544 0 0.0008853600000000001 0 0.00088546 3.3 0.0008853800000000001 3.3 0.00088548 0 0.0008854 0 0.0008855 3.3 0.00088542 3.3 0.00088552 0 0.00088544 0 0.00088554 3.3 0.00088546 3.3 0.00088556 0 0.00088548 0 0.00088558 3.3 0.0008855 3.3 0.0008856 0 0.00088552 0 0.0008856199999999999 3.3 0.00088554 3.3 0.0008856399999999999 0 0.0008855600000000001 0 0.00088566 3.3 0.0008855800000000001 3.3 0.00088568 0 0.0008856000000000001 0 0.0008857 3.3 0.00088562 3.3 0.00088572 0 0.00088564 0 0.00088574 3.3 0.00088566 3.3 0.00088576 0 0.00088568 0 0.00088578 3.3 0.0008857 3.3 0.0008858 0 0.00088572 0 0.0008858199999999999 3.3 0.00088574 3.3 0.0008858399999999999 0 0.0008857600000000001 0 0.00088586 3.3 0.0008857800000000001 3.3 0.00088588 0 0.0008858000000000001 0 0.0008859 3.3 0.00088582 3.3 0.00088592 0 0.00088584 0 0.00088594 3.3 0.00088586 3.3 0.00088596 0 0.00088588 0 0.00088598 3.3 0.0008859 3.3 0.000886 0 0.00088592 0 0.00088602 3.3 0.00088594 3.3 0.0008860399999999999 0 0.00088596 0 0.0008860599999999999 3.3 0.0008859800000000001 3.3 0.00088608 0 0.0008860000000000001 0 0.0008861 3.3 0.0008860200000000001 3.3 0.00088612 0 0.00088604 0 0.00088614 3.3 0.00088606 3.3 0.00088616 0 0.00088608 0 0.00088618 3.3 0.0008861 3.3 0.0008862 0 0.00088612 0 0.00088622 3.3 0.00088614 3.3 0.0008862399999999999 0 0.00088616 0 0.0008862599999999999 3.3 0.0008861800000000001 3.3 0.00088628 0 0.0008862000000000001 0 0.0008863 3.3 0.0008862200000000001 3.3 0.00088632 0 0.00088624 0 0.00088634 3.3 0.00088626 3.3 0.00088636 0 0.00088628 0 0.00088638 3.3 0.0008863 3.3 0.0008864 0 0.00088632 0 0.00088642 3.3 0.00088634 3.3 0.00088644 0 0.00088636 0 0.0008864599999999999 3.3 0.00088638 3.3 0.0008864799999999999 0 0.0008864000000000001 0 0.0008865 3.3 0.0008864200000000001 3.3 0.00088652 0 0.0008864400000000001 0 0.00088654 3.3 0.00088646 3.3 0.00088656 0 0.00088648 0 0.00088658 3.3 0.0008865 3.3 0.0008866 0 0.00088652 0 0.00088662 3.3 0.00088654 3.3 0.00088664 0 0.00088656 0 0.0008866599999999999 3.3 0.00088658 3.3 0.0008866799999999999 0 0.0008866000000000001 0 0.0008867 3.3 0.0008866200000000001 3.3 0.00088672 0 0.0008866400000000001 0 0.00088674 3.3 0.00088666 3.3 0.00088676 0 0.00088668 0 0.00088678 3.3 0.0008867 3.3 0.0008868 0 0.00088672 0 0.00088682 3.3 0.00088674 3.3 0.00088684 0 0.00088676 0 0.00088686 3.3 0.00088678 3.3 0.0008868799999999999 0 0.0008868 0 0.0008868999999999999 3.3 0.0008868200000000001 3.3 0.00088692 0 0.0008868400000000001 0 0.00088694 3.3 0.0008868600000000001 3.3 0.00088696 0 0.00088688 0 0.00088698 3.3 0.0008869 3.3 0.000887 0 0.00088692 0 0.00088702 3.3 0.00088694 3.3 0.00088704 0 0.00088696 0 0.00088706 3.3 0.00088698 3.3 0.0008870799999999999 0 0.000887 0 0.0008870999999999999 3.3 0.0008870200000000001 3.3 0.00088712 0 0.0008870400000000001 0 0.00088714 3.3 0.0008870600000000001 3.3 0.00088716 0 0.00088708 0 0.00088718 3.3 0.0008871 3.3 0.0008872 0 0.00088712 0 0.00088722 3.3 0.00088714 3.3 0.00088724 0 0.00088716 0 0.00088726 3.3 0.00088718 3.3 0.00088728 0 0.0008872 0 0.0008872999999999999 3.3 0.0008872200000000001 3.3 0.00088732 0 0.0008872400000000001 0 0.00088734 3.3 0.0008872600000000001 3.3 0.00088736 0 0.0008872800000000001 0 0.00088738 3.3 0.0008873 3.3 0.0008874 0 0.00088732 0 0.00088742 3.3 0.00088734 3.3 0.00088744 0 0.00088736 0 0.00088746 3.3 0.00088738 3.3 0.00088748 0 0.0008874 0 0.0008874999999999999 3.3 0.00088742 3.3 0.0008875199999999999 0 0.0008874400000000001 0 0.00088754 3.3 0.0008874600000000001 3.3 0.00088756 0 0.0008874800000000001 0 0.00088758 3.3 0.0008875 3.3 0.0008876 0 0.00088752 0 0.00088762 3.3 0.00088754 3.3 0.00088764 0 0.00088756 0 0.00088766 3.3 0.00088758 3.3 0.00088768 0 0.0008876 0 0.0008877 3.3 0.00088762 3.3 0.0008877199999999999 0 0.0008876400000000001 0 0.00088774 3.3 0.0008876600000000001 3.3 0.00088776 0 0.0008876800000000001 0 0.00088778 3.3 0.0008877000000000001 3.3 0.0008878 0 0.00088772 0 0.00088782 3.3 0.00088774 3.3 0.00088784 0 0.00088776 0 0.00088786 3.3 0.00088778 3.3 0.00088788 0 0.0008878 0 0.0008879 3.3 0.00088782 3.3 0.0008879199999999999 0 0.00088784 0 0.0008879399999999999 3.3 0.0008878600000000001 3.3 0.00088796 0 0.0008878800000000001 0 0.00088798 3.3 0.0008879000000000001 3.3 0.000888 0 0.00088792 0 0.00088802 3.3 0.00088794 3.3 0.00088804 0 0.00088796 0 0.00088806 3.3 0.00088798 3.3 0.00088808 0 0.000888 0 0.0008881 3.3 0.00088802 3.3 0.00088812 0 0.00088804 0 0.0008881399999999999 3.3 0.0008880600000000001 3.3 0.00088816 0 0.0008880800000000001 0 0.00088818 3.3 0.0008881000000000001 3.3 0.0008882 0 0.0008881200000000001 0 0.00088822 3.3 0.00088814 3.3 0.00088824 0 0.00088816 0 0.00088826 3.3 0.00088818 3.3 0.00088828 0 0.0008882 0 0.0008883 3.3 0.00088822 3.3 0.00088832 0 0.00088824 0 0.0008883399999999999 3.3 0.00088826 3.3 0.0008883599999999999 0 0.0008882800000000001 0 0.00088838 3.3 0.0008883000000000001 3.3 0.0008884 0 0.0008883200000000001 0 0.00088842 3.3 0.00088834 3.3 0.00088844 0 0.00088836 0 0.00088846 3.3 0.00088838 3.3 0.00088848 0 0.0008884 0 0.0008885 3.3 0.00088842 3.3 0.00088852 0 0.00088844 0 0.00088854 3.3 0.00088846 3.3 0.0008885599999999999 0 0.0008884800000000001 0 0.00088858 3.3 0.0008885000000000001 3.3 0.0008886 0 0.0008885200000000001 0 0.00088862 3.3 0.0008885400000000001 3.3 0.00088864 0 0.00088856 0 0.00088866 3.3 0.00088858 3.3 0.00088868 0 0.0008886 0 0.0008887 3.3 0.00088862 3.3 0.00088872 0 0.00088864 0 0.00088874 3.3 0.00088866 3.3 0.0008887599999999999 0 0.00088868 0 0.0008887799999999999 3.3 0.0008887000000000001 3.3 0.0008888 0 0.0008887200000000001 0 0.00088882 3.3 0.0008887400000000001 3.3 0.00088884 0 0.00088876 0 0.00088886 3.3 0.00088878 3.3 0.00088888 0 0.0008888 0 0.0008889 3.3 0.00088882 3.3 0.00088892 0 0.00088884 0 0.00088894 3.3 0.00088886 3.3 0.0008889599999999999 0 0.00088888 0 0.0008889799999999999 3.3 0.0008889000000000001 3.3 0.000889 0 0.0008889200000000001 0 0.00088902 3.3 0.0008889400000000001 3.3 0.00088904 0 0.00088896 0 0.00088906 3.3 0.00088898 3.3 0.00088908 0 0.000889 0 0.0008891 3.3 0.00088902 3.3 0.00088912 0 0.00088904 0 0.00088914 3.3 0.00088906 3.3 0.00088916 0 0.00088908 0 0.0008891799999999999 3.3 0.0008891 3.3 0.0008891999999999999 0 0.0008891200000000001 0 0.00088922 3.3 0.0008891400000000001 3.3 0.00088924 0 0.0008891600000000001 0 0.00088926 3.3 0.00088918 3.3 0.00088928 0 0.0008892 0 0.0008893 3.3 0.00088922 3.3 0.00088932 0 0.00088924 0 0.00088934 3.3 0.00088926 3.3 0.00088936 0 0.00088928 0 0.0008893799999999999 3.3 0.0008893 3.3 0.0008893999999999999 0 0.0008893200000000001 0 0.00088942 3.3 0.0008893400000000001 3.3 0.00088944 0 0.0008893600000000001 0 0.00088946 3.3 0.00088938 3.3 0.00088948 0 0.0008894 0 0.0008895 3.3 0.00088942 3.3 0.00088952 0 0.00088944 0 0.00088954 3.3 0.00088946 3.3 0.00088956 0 0.00088948 0 0.00088958 3.3 0.0008895 3.3 0.0008895999999999999 0 0.00088952 0 0.0008896199999999999 3.3 0.0008895400000000001 3.3 0.00088964 0 0.0008895600000000001 0 0.00088966 3.3 0.0008895800000000001 3.3 0.00088968 0 0.0008896 0 0.0008897 3.3 0.00088962 3.3 0.00088972 0 0.00088964 0 0.00088974 3.3 0.00088966 3.3 0.00088976 0 0.00088968 0 0.00088978 3.3 0.0008897 3.3 0.0008897999999999999 0 0.00088972 0 0.0008898199999999999 3.3 0.0008897400000000001 3.3 0.00088984 0 0.0008897600000000001 0 0.00088986 3.3 0.0008897800000000001 3.3 0.00088988 0 0.0008898 0 0.0008899 3.3 0.00088982 3.3 0.00088992 0 0.00088984 0 0.00088994 3.3 0.00088986 3.3 0.00088996 0 0.00088988 0 0.00088998 3.3 0.0008899 3.3 0.00089 0 0.00088992 0 0.0008900199999999999 3.3 0.00088994 3.3 0.0008900399999999999 0 0.0008899600000000001 0 0.00089006 3.3 0.0008899800000000001 3.3 0.00089008 0 0.0008900000000000001 0 0.0008901 3.3 0.00089002 3.3 0.00089012 0 0.00089004 0 0.00089014 3.3 0.00089006 3.3 0.00089016 0 0.00089008 0 0.00089018 3.3 0.0008901 3.3 0.0008902 0 0.00089012 0 0.0008902199999999999 3.3 0.00089014 3.3 0.0008902399999999999 0 0.0008901600000000001 0 0.00089026 3.3 0.0008901800000000001 3.3 0.00089028 0 0.0008902000000000001 0 0.0008903 3.3 0.00089022 3.3 0.00089032 0 0.00089024 0 0.00089034 3.3 0.00089026 3.3 0.00089036 0 0.00089028 0 0.00089038 3.3 0.0008903 3.3 0.0008904 0 0.00089032 0 0.00089042 3.3 0.00089034 3.3 0.0008904399999999999 0 0.0008903600000000001 0 0.00089046 3.3 0.0008903800000000001 3.3 0.00089048 0 0.0008904000000000001 0 0.0008905 3.3 0.0008904200000000001 3.3 0.00089052 0 0.00089044 0 0.00089054 3.3 0.00089046 3.3 0.00089056 0 0.00089048 0 0.00089058 3.3 0.0008905 3.3 0.0008906 0 0.00089052 0 0.00089062 3.3 0.00089054 3.3 0.0008906399999999999 0 0.00089056 0 0.0008906599999999999 3.3 0.0008905800000000001 3.3 0.00089068 0 0.0008906000000000001 0 0.0008907 3.3 0.0008906200000000001 3.3 0.00089072 0 0.00089064 0 0.00089074 3.3 0.00089066 3.3 0.00089076 0 0.00089068 0 0.00089078 3.3 0.0008907 3.3 0.0008908 0 0.00089072 0 0.00089082 3.3 0.00089074 3.3 0.00089084 0 0.00089076 0 0.0008908599999999999 3.3 0.0008907800000000001 3.3 0.00089088 0 0.0008908000000000001 0 0.0008909 3.3 0.0008908200000000001 3.3 0.00089092 0 0.0008908400000000001 0 0.00089094 3.3 0.00089086 3.3 0.00089096 0 0.00089088 0 0.00089098 3.3 0.0008909 3.3 0.000891 0 0.00089092 0 0.00089102 3.3 0.00089094 3.3 0.00089104 0 0.00089096 0 0.0008910599999999999 3.3 0.00089098 3.3 0.0008910799999999999 0 0.0008910000000000001 0 0.0008911 3.3 0.0008910200000000001 3.3 0.00089112 0 0.0008910400000000001 0 0.00089114 3.3 0.00089106 3.3 0.00089116 0 0.00089108 0 0.00089118 3.3 0.0008911 3.3 0.0008912 0 0.00089112 0 0.00089122 3.3 0.00089114 3.3 0.00089124 0 0.00089116 0 0.00089126 3.3 0.00089118 3.3 0.0008912799999999999 0 0.0008912000000000001 0 0.0008913 3.3 0.0008912200000000001 3.3 0.00089132 0 0.0008912400000000001 0 0.00089134 3.3 0.0008912600000000001 3.3 0.00089136 0 0.00089128 0 0.00089138 3.3 0.0008913 3.3 0.0008914 0 0.00089132 0 0.00089142 3.3 0.00089134 3.3 0.00089144 0 0.00089136 0 0.00089146 3.3 0.00089138 3.3 0.0008914799999999999 0 0.0008914 0 0.0008914999999999999 3.3 0.0008914200000000001 3.3 0.00089152 0 0.0008914400000000001 0 0.00089154 3.3 0.0008914600000000001 3.3 0.00089156 0 0.00089148 0 0.00089158 3.3 0.0008915 3.3 0.0008916 0 0.00089152 0 0.00089162 3.3 0.00089154 3.3 0.00089164 0 0.00089156 0 0.00089166 3.3 0.00089158 3.3 0.00089168 0 0.0008916 0 0.0008916999999999999 3.3 0.0008916200000000001 3.3 0.00089172 0 0.0008916400000000001 0 0.00089174 3.3 0.0008916600000000001 3.3 0.00089176 0 0.0008916800000000001 0 0.00089178 3.3 0.0008917 3.3 0.0008918 0 0.00089172 0 0.00089182 3.3 0.00089174 3.3 0.00089184 0 0.00089176 0 0.00089186 3.3 0.00089178 3.3 0.00089188 0 0.0008918 0 0.0008918999999999999 3.3 0.00089182 3.3 0.0008919199999999999 0 0.0008918400000000001 0 0.00089194 3.3 0.0008918600000000001 3.3 0.00089196 0 0.0008918800000000001 0 0.00089198 3.3 0.0008919 3.3 0.000892 0 0.00089192 0 0.00089202 3.3 0.00089194 3.3 0.00089204 0 0.00089196 0 0.00089206 3.3 0.00089198 3.3 0.00089208 0 0.000892 0 0.0008921 3.3 0.00089202 3.3 0.0008921199999999999 0 0.0008920400000000001 0 0.00089214 3.3 0.0008920600000000001 3.3 0.00089216 0 0.0008920800000000001 0 0.00089218 3.3 0.0008921000000000001 3.3 0.0008922 0 0.00089212 0 0.00089222 3.3 0.00089214 3.3 0.00089224 0 0.00089216 0 0.00089226 3.3 0.00089218 3.3 0.00089228 0 0.0008922 0 0.0008923 3.3 0.00089222 3.3 0.0008923199999999999 0 0.00089224 0 0.0008923399999999999 3.3 0.0008922600000000001 3.3 0.00089236 0 0.0008922800000000001 0 0.00089238 3.3 0.0008923000000000001 3.3 0.0008924 0 0.00089232 0 0.00089242 3.3 0.00089234 3.3 0.00089244 0 0.00089236 0 0.00089246 3.3 0.00089238 3.3 0.00089248 0 0.0008924 0 0.0008925 3.3 0.00089242 3.3 0.0008925199999999999 0 0.00089244 0 0.0008925399999999999 3.3 0.0008924600000000001 3.3 0.00089256 0 0.0008924800000000001 0 0.00089258 3.3 0.0008925000000000001 3.3 0.0008926 0 0.00089252 0 0.00089262 3.3 0.00089254 3.3 0.00089264 0 0.00089256 0 0.00089266 3.3 0.00089258 3.3 0.00089268 0 0.0008926 0 0.0008927 3.3 0.00089262 3.3 0.00089272 0 0.00089264 0 0.0008927399999999999 3.3 0.00089266 3.3 0.0008927599999999999 0 0.0008926800000000001 0 0.00089278 3.3 0.0008927000000000001 3.3 0.0008928 0 0.0008927200000000001 0 0.00089282 3.3 0.00089274 3.3 0.00089284 0 0.00089276 0 0.00089286 3.3 0.00089278 3.3 0.00089288 0 0.0008928 0 0.0008929 3.3 0.00089282 3.3 0.00089292 0 0.00089284 0 0.0008929399999999999 3.3 0.00089286 3.3 0.0008929599999999999 0 0.0008928800000000001 0 0.00089298 3.3 0.0008929000000000001 3.3 0.000893 0 0.0008929200000000001 0 0.00089302 3.3 0.00089294 3.3 0.00089304 0 0.00089296 0 0.00089306 3.3 0.00089298 3.3 0.00089308 0 0.000893 0 0.0008931 3.3 0.00089302 3.3 0.00089312 0 0.00089304 0 0.00089314 3.3 0.00089306 3.3 0.0008931599999999999 0 0.00089308 0 0.0008931799999999999 3.3 0.0008931000000000001 3.3 0.0008932 0 0.0008931200000000001 0 0.00089322 3.3 0.0008931400000000001 3.3 0.00089324 0 0.00089316 0 0.00089326 3.3 0.00089318 3.3 0.00089328 0 0.0008932 0 0.0008933 3.3 0.00089322 3.3 0.00089332 0 0.00089324 0 0.00089334 3.3 0.00089326 3.3 0.0008933599999999999 0 0.00089328 0 0.0008933799999999999 3.3 0.0008933000000000001 3.3 0.0008934 0 0.0008933200000000001 0 0.00089342 3.3 0.0008933400000000001 3.3 0.00089344 0 0.00089336 0 0.00089346 3.3 0.00089338 3.3 0.00089348 0 0.0008934 0 0.0008935 3.3 0.00089342 3.3 0.00089352 0 0.00089344 0 0.00089354 3.3 0.00089346 3.3 0.00089356 0 0.00089348 0 0.0008935799999999999 3.3 0.0008935 3.3 0.0008935999999999999 0 0.0008935200000000001 0 0.00089362 3.3 0.0008935400000000001 3.3 0.00089364 0 0.0008935600000000001 0 0.00089366 3.3 0.00089358 3.3 0.00089368 0 0.0008936 0 0.0008937 3.3 0.00089362 3.3 0.00089372 0 0.00089364 0 0.00089374 3.3 0.00089366 3.3 0.00089376 0 0.00089368 0 0.0008937799999999999 3.3 0.0008937 3.3 0.0008937999999999999 0 0.0008937200000000001 0 0.00089382 3.3 0.0008937400000000001 3.3 0.00089384 0 0.0008937600000000001 0 0.00089386 3.3 0.00089378 3.3 0.00089388 0 0.0008938 0 0.0008939 3.3 0.00089382 3.3 0.00089392 0 0.00089384 0 0.00089394 3.3 0.00089386 3.3 0.00089396 0 0.00089388 0 0.00089398 3.3 0.0008939 3.3 0.0008939999999999999 0 0.0008939200000000001 0 0.00089402 3.3 0.0008939400000000001 3.3 0.00089404 0 0.0008939600000000001 0 0.00089406 3.3 0.0008939800000000001 3.3 0.00089408 0 0.000894 0 0.0008941 3.3 0.00089402 3.3 0.00089412 0 0.00089404 0 0.00089414 3.3 0.00089406 3.3 0.00089416 0 0.00089408 0 0.00089418 3.3 0.0008941 3.3 0.0008941999999999999 0 0.00089412 0 0.0008942199999999999 3.3 0.0008941400000000001 3.3 0.00089424 0 0.0008941600000000001 0 0.00089426 3.3 0.0008941800000000001 3.3 0.00089428 0 0.0008942 0 0.0008943 3.3 0.00089422 3.3 0.00089432 0 0.00089424 0 0.00089434 3.3 0.00089426 3.3 0.00089436 0 0.00089428 0 0.00089438 3.3 0.0008943 3.3 0.0008944 0 0.00089432 0 0.0008944199999999999 3.3 0.0008943400000000001 3.3 0.00089444 0 0.0008943600000000001 0 0.00089446 3.3 0.0008943800000000001 3.3 0.00089448 0 0.0008944000000000001 0 0.0008945 3.3 0.00089442 3.3 0.00089452 0 0.00089444 0 0.00089454 3.3 0.00089446 3.3 0.00089456 0 0.00089448 0 0.00089458 3.3 0.0008945 3.3 0.0008946 0 0.00089452 0 0.0008946199999999999 3.3 0.00089454 3.3 0.0008946399999999999 0 0.0008945600000000001 0 0.00089466 3.3 0.0008945800000000001 3.3 0.00089468 0 0.0008946000000000001 0 0.0008947 3.3 0.00089462 3.3 0.00089472 0 0.00089464 0 0.00089474 3.3 0.00089466 3.3 0.00089476 0 0.00089468 0 0.00089478 3.3 0.0008947 3.3 0.0008948 0 0.00089472 0 0.00089482 3.3 0.00089474 3.3 0.0008948399999999999 0 0.0008947600000000001 0 0.00089486 3.3 0.0008947800000000001 3.3 0.00089488 0 0.0008948000000000001 0 0.0008949 3.3 0.0008948200000000001 3.3 0.00089492 0 0.00089484 0 0.00089494 3.3 0.00089486 3.3 0.00089496 0 0.00089488 0 0.00089498 3.3 0.0008949 3.3 0.000895 0 0.00089492 0 0.00089502 3.3 0.00089494 3.3 0.0008950399999999999 0 0.00089496 0 0.0008950599999999999 3.3 0.0008949800000000001 3.3 0.00089508 0 0.0008950000000000001 0 0.0008951 3.3 0.0008950200000000001 3.3 0.00089512 0 0.00089504 0 0.00089514 3.3 0.00089506 3.3 0.00089516 0 0.00089508 0 0.00089518 3.3 0.0008951 3.3 0.0008952 0 0.00089512 0 0.00089522 3.3 0.00089514 3.3 0.00089524 0 0.00089516 0 0.0008952599999999999 3.3 0.0008951800000000001 3.3 0.00089528 0 0.0008952000000000001 0 0.0008953 3.3 0.0008952200000000001 3.3 0.00089532 0 0.0008952400000000001 0 0.00089534 3.3 0.00089526 3.3 0.00089536 0 0.00089528 0 0.00089538 3.3 0.0008953 3.3 0.0008954 0 0.00089532 0 0.00089542 3.3 0.00089534 3.3 0.00089544 0 0.00089536 0 0.0008954599999999999 3.3 0.00089538 3.3 0.0008954799999999999 0 0.0008954000000000001 0 0.0008955 3.3 0.0008954200000000001 3.3 0.00089552 0 0.0008954400000000001 0 0.00089554 3.3 0.00089546 3.3 0.00089556 0 0.00089548 0 0.00089558 3.3 0.0008955 3.3 0.0008956 0 0.00089552 0 0.00089562 3.3 0.00089554 3.3 0.00089564 0 0.00089556 0 0.0008956599999999999 3.3 0.00089558 3.3 0.0008956799999999999 0 0.0008956000000000001 0 0.0008957 3.3 0.0008956200000000001 3.3 0.00089572 0 0.0008956400000000001 0 0.00089574 3.3 0.00089566 3.3 0.00089576 0 0.00089568 0 0.00089578 3.3 0.0008957 3.3 0.0008958 0 0.00089572 0 0.00089582 3.3 0.00089574 3.3 0.00089584 0 0.00089576 0 0.00089586 3.3 0.00089578 3.3 0.0008958799999999999 0 0.0008958 0 0.0008958999999999999 3.3 0.0008958200000000001 3.3 0.00089592 0 0.0008958400000000001 0 0.00089594 3.3 0.0008958600000000001 3.3 0.00089596 0 0.00089588 0 0.00089598 3.3 0.0008959 3.3 0.000896 0 0.00089592 0 0.00089602 3.3 0.00089594 3.3 0.00089604 0 0.00089596 0 0.00089606 3.3 0.00089598 3.3 0.0008960799999999999 0 0.000896 0 0.0008960999999999999 3.3 0.0008960200000000001 3.3 0.00089612 0 0.0008960400000000001 0 0.00089614 3.3 0.0008960600000000001 3.3 0.00089616 0 0.00089608 0 0.00089618 3.3 0.0008961 3.3 0.0008962 0 0.00089612 0 0.00089622 3.3 0.00089614 3.3 0.00089624 0 0.00089616 0 0.00089626 3.3 0.00089618 3.3 0.00089628 0 0.0008962 0 0.0008962999999999999 3.3 0.00089622 3.3 0.0008963199999999999 0 0.0008962400000000001 0 0.00089634 3.3 0.0008962600000000001 3.3 0.00089636 0 0.0008962800000000001 0 0.00089638 3.3 0.0008963 3.3 0.0008964 0 0.00089632 0 0.00089642 3.3 0.00089634 3.3 0.00089644 0 0.00089636 0 0.00089646 3.3 0.00089638 3.3 0.00089648 0 0.0008964 0 0.0008964999999999999 3.3 0.00089642 3.3 0.0008965199999999999 0 0.0008964400000000001 0 0.00089654 3.3 0.0008964600000000001 3.3 0.00089656 0 0.0008964800000000001 0 0.00089658 3.3 0.0008965 3.3 0.0008966 0 0.00089652 0 0.00089662 3.3 0.00089654 3.3 0.00089664 0 0.00089656 0 0.00089666 3.3 0.00089658 3.3 0.00089668 0 0.0008966 0 0.0008967 3.3 0.00089662 3.3 0.0008967199999999999 0 0.00089664 0 0.0008967399999999999 3.3 0.0008966600000000001 3.3 0.00089676 0 0.0008966800000000001 0 0.00089678 3.3 0.0008967000000000001 3.3 0.0008968 0 0.00089672 0 0.00089682 3.3 0.00089674 3.3 0.00089684 0 0.00089676 0 0.00089686 3.3 0.00089678 3.3 0.00089688 0 0.0008968 0 0.0008969 3.3 0.00089682 3.3 0.0008969199999999999 0 0.00089684 0 0.0008969399999999999 3.3 0.0008968600000000001 3.3 0.00089696 0 0.0008968800000000001 0 0.00089698 3.3 0.0008969000000000001 3.3 0.000897 0 0.00089692 0 0.00089702 3.3 0.00089694 3.3 0.00089704 0 0.00089696 0 0.00089706 3.3 0.00089698 3.3 0.00089708 0 0.000897 0 0.0008971 3.3 0.00089702 3.3 0.00089712 0 0.00089704 0 0.0008971399999999999 3.3 0.00089706 3.3 0.0008971599999999999 0 0.0008970800000000001 0 0.00089718 3.3 0.0008971000000000001 3.3 0.0008972 0 0.0008971200000000001 0 0.00089722 3.3 0.00089714 3.3 0.00089724 0 0.00089716 0 0.00089726 3.3 0.00089718 3.3 0.00089728 0 0.0008972 0 0.0008973 3.3 0.00089722 3.3 0.00089732 0 0.00089724 0 0.0008973399999999999 3.3 0.00089726 3.3 0.0008973599999999999 0 0.0008972800000000001 0 0.00089738 3.3 0.0008973000000000001 3.3 0.0008974 0 0.0008973200000000001 0 0.00089742 3.3 0.00089734 3.3 0.00089744 0 0.00089736 0 0.00089746 3.3 0.00089738 3.3 0.00089748 0 0.0008974 0 0.0008975 3.3 0.00089742 3.3 0.00089752 0 0.00089744 0 0.00089754 3.3 0.00089746 3.3 0.0008975599999999999 0 0.0008974800000000001 0 0.00089758 3.3 0.0008975000000000001 3.3 0.0008976 0 0.0008975200000000001 0 0.00089762 3.3 0.0008975400000000001 3.3 0.00089764 0 0.00089756 0 0.00089766 3.3 0.00089758 3.3 0.00089768 0 0.0008976 0 0.0008977 3.3 0.00089762 3.3 0.00089772 0 0.00089764 0 0.00089774 3.3 0.00089766 3.3 0.0008977599999999999 0 0.00089768 0 0.0008977799999999999 3.3 0.0008977000000000001 3.3 0.0008978 0 0.0008977200000000001 0 0.00089782 3.3 0.0008977400000000001 3.3 0.00089784 0 0.00089776 0 0.00089786 3.3 0.00089778 3.3 0.00089788 0 0.0008978 0 0.0008979 3.3 0.00089782 3.3 0.00089792 0 0.00089784 0 0.00089794 3.3 0.00089786 3.3 0.00089796 0 0.00089788 0 0.0008979799999999999 3.3 0.0008979000000000001 3.3 0.000898 0 0.0008979200000000001 0 0.00089802 3.3 0.0008979400000000001 3.3 0.00089804 0 0.0008979600000000001 0 0.00089806 3.3 0.00089798 3.3 0.00089808 0 0.000898 0 0.0008981 3.3 0.00089802 3.3 0.00089812 0 0.00089804 0 0.00089814 3.3 0.00089806 3.3 0.00089816 0 0.00089808 0 0.0008981799999999999 3.3 0.0008981 3.3 0.0008981999999999999 0 0.0008981200000000001 0 0.00089822 3.3 0.0008981400000000001 3.3 0.00089824 0 0.0008981600000000001 0 0.00089826 3.3 0.00089818 3.3 0.00089828 0 0.0008982 0 0.0008983 3.3 0.00089822 3.3 0.00089832 0 0.00089824 0 0.00089834 3.3 0.00089826 3.3 0.00089836 0 0.00089828 0 0.00089838 3.3 0.0008983 3.3 0.0008983999999999999 0 0.0008983200000000001 0 0.00089842 3.3 0.0008983400000000001 3.3 0.00089844 0 0.0008983600000000001 0 0.00089846 3.3 0.0008983800000000001 3.3 0.00089848 0 0.0008984 0 0.0008985 3.3 0.00089842 3.3 0.00089852 0 0.00089844 0 0.00089854 3.3 0.00089846 3.3 0.00089856 0 0.00089848 0 0.00089858 3.3 0.0008985 3.3 0.0008985999999999999 0 0.00089852 0 0.0008986199999999999 3.3 0.0008985400000000001 3.3 0.00089864 0 0.0008985600000000001 0 0.00089866 3.3 0.0008985800000000001 3.3 0.00089868 0 0.0008986 0 0.0008987 3.3 0.00089862 3.3 0.00089872 0 0.00089864 0 0.00089874 3.3 0.00089866 3.3 0.00089876 0 0.00089868 0 0.00089878 3.3 0.0008987 3.3 0.0008988 0 0.00089872 0 0.0008988199999999999 3.3 0.0008987400000000001 3.3 0.00089884 0 0.0008987600000000001 0 0.00089886 3.3 0.0008987800000000001 3.3 0.00089888 0 0.0008988000000000001 0 0.0008989 3.3 0.00089882 3.3 0.00089892 0 0.00089884 0 0.00089894 3.3 0.00089886 3.3 0.00089896 0 0.00089888 0 0.00089898 3.3 0.0008989 3.3 0.000899 0 0.00089892 0 0.0008990199999999999 3.3 0.00089894 3.3 0.0008990399999999999 0 0.0008989600000000001 0 0.00089906 3.3 0.0008989800000000001 3.3 0.00089908 0 0.0008990000000000001 0 0.0008991 3.3 0.00089902 3.3 0.00089912 0 0.00089904 0 0.00089914 3.3 0.00089906 3.3 0.00089916 0 0.00089908 0 0.00089918 3.3 0.0008991 3.3 0.0008992 0 0.00089912 0 0.0008992199999999999 3.3 0.00089914 3.3 0.0008992399999999999 0 0.0008991600000000001 0 0.00089926 3.3 0.0008991800000000001 3.3 0.00089928 0 0.0008992000000000001 0 0.0008993 3.3 0.00089922 3.3 0.00089932 0 0.00089924 0 0.00089934 3.3 0.00089926 3.3 0.00089936 0 0.00089928 0 0.00089938 3.3 0.0008993 3.3 0.0008994 0 0.00089932 0 0.00089942 3.3 0.00089934 3.3 0.0008994399999999999 0 0.00089936 0 0.0008994599999999999 3.3 0.0008993800000000001 3.3 0.00089948 0 0.0008994000000000001 0 0.0008995 3.3 0.0008994200000000001 3.3 0.00089952 0 0.00089944 0 0.00089954 3.3 0.00089946 3.3 0.00089956 0 0.00089948 0 0.00089958 3.3 0.0008995 3.3 0.0008996 0 0.00089952 0 0.00089962 3.3 0.00089954 3.3 0.0008996399999999999 0 0.00089956 0 0.0008996599999999999 3.3 0.0008995800000000001 3.3 0.00089968 0 0.0008996000000000001 0 0.0008997 3.3 0.0008996200000000001 3.3 0.00089972 0 0.00089964 0 0.00089974 3.3 0.00089966 3.3 0.00089976 0 0.00089968 0 0.00089978 3.3 0.0008997 3.3 0.0008998 0 0.00089972 0 0.00089982 3.3 0.00089974 3.3 0.00089984 0 0.00089976 0 0.0008998599999999999 3.3 0.00089978 3.3 0.0008998799999999999 0 0.0008998000000000001 0 0.0008999 3.3 0.0008998200000000001 3.3 0.00089992 0 0.0008998400000000001 0 0.00089994 3.3 0.00089986 3.3 0.00089996 0 0.00089988 0 0.00089998 3.3 0.0008999 3.3 0.0009 0 0.00089992 0 0.00090002 3.3 0.00089994 3.3 0.00090004 0 0.00089996 0 0.0009000599999999999 3.3 0.00089998 3.3 0.0009000799999999999 0 0.0009000000000000001 0 0.0009001 3.3 0.0009000200000000001 3.3 0.00090012 0 0.0009000400000000001 0 0.00090014 3.3 0.00090006 3.3 0.00090016 0 0.00090008 0 0.00090018 3.3 0.0009001 3.3 0.0009002 0 0.00090012 0 0.00090022 3.3 0.00090014 3.3 0.00090024 0 0.00090016 0 0.00090026 3.3 0.00090018 3.3 0.0009002799999999999 0 0.0009002 0 0.0009002999999999999 3.3 0.0009002200000000001 3.3 0.00090032 0 0.0009002400000000001 0 0.00090034 3.3 0.0009002600000000001 3.3 0.00090036 0 0.00090028 0 0.00090038 3.3 0.0009003 3.3 0.0009004 0 0.00090032 0 0.00090042 3.3 0.00090034 3.3 0.00090044 0 0.00090036 0 0.00090046 3.3 0.00090038 3.3 0.0009004799999999999 0 0.0009004 0 0.0009004999999999999 3.3 0.0009004200000000001 3.3 0.00090052 0 0.0009004400000000001 0 0.00090054 3.3 0.0009004600000000001 3.3 0.00090056 0 0.00090048 0 0.00090058 3.3 0.0009005 3.3 0.0009006 0 0.00090052 0 0.00090062 3.3 0.00090054 3.3 0.00090064 0 0.00090056 0 0.00090066 3.3 0.00090058 3.3 0.00090068 0 0.0009006 0 0.0009006999999999999 3.3 0.00090062 3.3 0.0009007199999999999 0 0.0009006400000000001 0 0.00090074 3.3 0.0009006600000000001 3.3 0.00090076 0 0.0009006800000000001 0 0.00090078 3.3 0.0009007 3.3 0.0009008 0 0.00090072 0 0.00090082 3.3 0.00090074 3.3 0.00090084 0 0.00090076 0 0.00090086 3.3 0.00090078 3.3 0.00090088 0 0.0009008 0 0.0009008999999999999 3.3 0.00090082 3.3 0.0009009199999999999 0 0.0009008400000000001 0 0.00090094 3.3 0.0009008600000000001 3.3 0.00090096 0 0.0009008800000000001 0 0.00090098 3.3 0.0009009 3.3 0.000901 0 0.00090092 0 0.00090102 3.3 0.00090094 3.3 0.00090104 0 0.00090096 0 0.00090106 3.3 0.00090098 3.3 0.00090108 0 0.000901 0 0.0009011 3.3 0.00090102 3.3 0.0009011199999999999 0 0.0009010400000000001 0 0.00090114 3.3 0.0009010600000000001 3.3 0.00090116 0 0.0009010800000000001 0 0.00090118 3.3 0.0009011000000000001 3.3 0.0009012 0 0.00090112 0 0.00090122 3.3 0.00090114 3.3 0.00090124 0 0.00090116 0 0.00090126 3.3 0.00090118 3.3 0.00090128 0 0.0009012 0 0.0009013 3.3 0.00090122 3.3 0.0009013199999999999 0 0.00090124 0 0.0009013399999999999 3.3 0.0009012600000000001 3.3 0.00090136 0 0.0009012800000000001 0 0.00090138 3.3 0.0009013000000000001 3.3 0.0009014 0 0.00090132 0 0.00090142 3.3 0.00090134 3.3 0.00090144 0 0.00090136 0 0.00090146 3.3 0.00090138 3.3 0.00090148 0 0.0009014 0 0.0009015 3.3 0.00090142 3.3 0.00090152 0 0.00090144 0 0.0009015399999999999 3.3 0.0009014600000000001 3.3 0.00090156 0 0.0009014800000000001 0 0.00090158 3.3 0.0009015000000000001 3.3 0.0009016 0 0.0009015200000000001 0 0.00090162 3.3 0.00090154 3.3 0.00090164 0 0.00090156 0 0.00090166 3.3 0.00090158 3.3 0.00090168 0 0.0009016 0 0.0009017 3.3 0.00090162 3.3 0.00090172 0 0.00090164 0 0.0009017399999999999 3.3 0.00090166 3.3 0.0009017599999999999 0 0.0009016800000000001 0 0.00090178 3.3 0.0009017000000000001 3.3 0.0009018 0 0.0009017200000000001 0 0.00090182 3.3 0.00090174 3.3 0.00090184 0 0.00090176 0 0.00090186 3.3 0.00090178 3.3 0.00090188 0 0.0009018 0 0.0009019 3.3 0.00090182 3.3 0.00090192 0 0.00090184 0 0.00090194 3.3 0.00090186 3.3 0.0009019599999999999 0 0.0009018800000000001 0 0.00090198 3.3 0.0009019000000000001 3.3 0.000902 0 0.0009019200000000001 0 0.00090202 3.3 0.0009019400000000001 3.3 0.00090204 0 0.00090196 0 0.00090206 3.3 0.00090198 3.3 0.00090208 0 0.000902 0 0.0009021 3.3 0.00090202 3.3 0.00090212 0 0.00090204 0 0.00090214 3.3 0.00090206 3.3 0.0009021599999999999 0 0.00090208 0 0.0009021799999999999 3.3 0.0009021000000000001 3.3 0.0009022 0 0.0009021200000000001 0 0.00090222 3.3 0.0009021400000000001 3.3 0.00090224 0 0.00090216 0 0.00090226 3.3 0.00090218 3.3 0.00090228 0 0.0009022 0 0.0009023 3.3 0.00090222 3.3 0.00090232 0 0.00090224 0 0.00090234 3.3 0.00090226 3.3 0.00090236 0 0.00090228 0 0.0009023799999999999 3.3 0.0009023000000000001 3.3 0.0009024 0 0.0009023200000000001 0 0.00090242 3.3 0.0009023400000000001 3.3 0.00090244 0 0.0009023600000000001 0 0.00090246 3.3 0.00090238 3.3 0.00090248 0 0.0009024 0 0.0009025 3.3 0.00090242 3.3 0.00090252 0 0.00090244 0 0.00090254 3.3 0.00090246 3.3 0.00090256 0 0.00090248 0 0.0009025799999999999 3.3 0.0009025 3.3 0.0009025999999999999 0 0.0009025200000000001 0 0.00090262 3.3 0.0009025400000000001 3.3 0.00090264 0 0.0009025600000000001 0 0.00090266 3.3 0.00090258 3.3 0.00090268 0 0.0009026 0 0.0009027 3.3 0.00090262 3.3 0.00090272 0 0.00090264 0 0.00090274 3.3 0.00090266 3.3 0.00090276 0 0.00090268 0 0.0009027799999999999 3.3 0.0009027 3.3 0.0009027999999999999 0 0.0009027200000000001 0 0.00090282 3.3 0.0009027400000000001 3.3 0.00090284 0 0.0009027600000000001 0 0.00090286 3.3 0.00090278 3.3 0.00090288 0 0.0009028 0 0.0009029 3.3 0.00090282 3.3 0.00090292 0 0.00090284 0 0.00090294 3.3 0.00090286 3.3 0.00090296 0 0.00090288 0 0.00090298 3.3 0.0009029 3.3 0.0009029999999999999 0 0.00090292 0 0.0009030199999999999 3.3 0.0009029400000000001 3.3 0.00090304 0 0.0009029600000000001 0 0.00090306 3.3 0.0009029800000000001 3.3 0.00090308 0 0.000903 0 0.0009031 3.3 0.00090302 3.3 0.00090312 0 0.00090304 0 0.00090314 3.3 0.00090306 3.3 0.00090316 0 0.00090308 0 0.00090318 3.3 0.0009031 3.3 0.0009031999999999999 0 0.00090312 0 0.0009032199999999999 3.3 0.0009031400000000001 3.3 0.00090324 0 0.0009031600000000001 0 0.00090326 3.3 0.0009031800000000001 3.3 0.00090328 0 0.0009032 0 0.0009033 3.3 0.00090322 3.3 0.00090332 0 0.00090324 0 0.00090334 3.3 0.00090326 3.3 0.00090336 0 0.00090328 0 0.00090338 3.3 0.0009033 3.3 0.0009034 0 0.00090332 0 0.0009034199999999999 3.3 0.00090334 3.3 0.0009034399999999999 0 0.0009033600000000001 0 0.00090346 3.3 0.0009033800000000001 3.3 0.00090348 0 0.0009034000000000001 0 0.0009035 3.3 0.00090342 3.3 0.00090352 0 0.00090344 0 0.00090354 3.3 0.00090346 3.3 0.00090356 0 0.00090348 0 0.00090358 3.3 0.0009035 3.3 0.0009036 0 0.00090352 0 0.0009036199999999999 3.3 0.00090354 3.3 0.0009036399999999999 0 0.0009035600000000001 0 0.00090366 3.3 0.0009035800000000001 3.3 0.00090368 0 0.0009036000000000001 0 0.0009037 3.3 0.00090362 3.3 0.00090372 0 0.00090364 0 0.00090374 3.3 0.00090366 3.3 0.00090376 0 0.00090368 0 0.00090378 3.3 0.0009037 3.3 0.0009038 0 0.00090372 0 0.00090382 3.3 0.00090374 3.3 0.0009038399999999999 0 0.00090376 0 0.0009038599999999999 3.3 0.0009037800000000001 3.3 0.00090388 0 0.0009038000000000001 0 0.0009039 3.3 0.0009038200000000001 3.3 0.00090392 0 0.00090384 0 0.00090394 3.3 0.00090386 3.3 0.00090396 0 0.00090388 0 0.00090398 3.3 0.0009039 3.3 0.000904 0 0.00090392 0 0.00090402 3.3 0.00090394 3.3 0.0009040399999999999 0 0.00090396 0 0.0009040599999999999 3.3 0.0009039800000000001 3.3 0.00090408 0 0.0009040000000000001 0 0.0009041 3.3 0.0009040200000000001 3.3 0.00090412 0 0.00090404 0 0.00090414 3.3 0.00090406 3.3 0.00090416 0 0.00090408 0 0.00090418 3.3 0.0009041 3.3 0.0009042 0 0.00090412 0 0.00090422 3.3 0.00090414 3.3 0.00090424 0 0.00090416 0 0.0009042599999999999 3.3 0.00090418 3.3 0.0009042799999999999 0 0.0009042000000000001 0 0.0009043 3.3 0.0009042200000000001 3.3 0.00090432 0 0.0009042400000000001 0 0.00090434 3.3 0.00090426 3.3 0.00090436 0 0.00090428 0 0.00090438 3.3 0.0009043 3.3 0.0009044 0 0.00090432 0 0.00090442 3.3 0.00090434 3.3 0.00090444 0 0.00090436 0 0.0009044599999999999 3.3 0.00090438 3.3 0.0009044799999999999 0 0.0009044000000000001 0 0.0009045 3.3 0.0009044200000000001 3.3 0.00090452 0 0.0009044400000000001 0 0.00090454 3.3 0.00090446 3.3 0.00090456 0 0.00090448 0 0.00090458 3.3 0.0009045 3.3 0.0009046 0 0.00090452 0 0.00090462 3.3 0.00090454 3.3 0.00090464 0 0.00090456 0 0.00090466 3.3 0.00090458 3.3 0.0009046799999999999 0 0.0009046000000000001 0 0.0009047 3.3 0.0009046200000000001 3.3 0.00090472 0 0.0009046400000000001 0 0.00090474 3.3 0.0009046600000000001 3.3 0.00090476 0 0.00090468 0 0.00090478 3.3 0.0009047 3.3 0.0009048 0 0.00090472 0 0.00090482 3.3 0.00090474 3.3 0.00090484 0 0.00090476 0 0.00090486 3.3 0.00090478 3.3 0.0009048799999999999 0 0.0009048 0 0.0009048999999999999 3.3 0.0009048200000000001 3.3 0.00090492 0 0.0009048400000000001 0 0.00090494 3.3 0.0009048600000000001 3.3 0.00090496 0 0.00090488 0 0.00090498 3.3 0.0009049 3.3 0.000905 0 0.00090492 0 0.00090502 3.3 0.00090494 3.3 0.00090504 0 0.00090496 0 0.00090506 3.3 0.00090498 3.3 0.00090508 0 0.000905 0 0.0009050999999999999 3.3 0.0009050200000000001 3.3 0.00090512 0 0.0009050400000000001 0 0.00090514 3.3 0.0009050600000000001 3.3 0.00090516 0 0.0009050800000000001 0 0.00090518 3.3 0.0009051 3.3 0.0009052 0 0.00090512 0 0.00090522 3.3 0.00090514 3.3 0.00090524 0 0.00090516 0 0.00090526 3.3 0.00090518 3.3 0.00090528 0 0.0009052 0 0.0009052999999999999 3.3 0.00090522 3.3 0.0009053199999999999 0 0.0009052400000000001 0 0.00090534 3.3 0.0009052600000000001 3.3 0.00090536 0 0.0009052800000000001 0 0.00090538 3.3 0.0009053 3.3 0.0009054 0 0.00090532 0 0.00090542 3.3 0.00090534 3.3 0.00090544 0 0.00090536 0 0.00090546 3.3 0.00090538 3.3 0.00090548 0 0.0009054 0 0.0009055 3.3 0.00090542 3.3 0.0009055199999999999 0 0.0009054400000000001 0 0.00090554 3.3 0.0009054600000000001 3.3 0.00090556 0 0.0009054800000000001 0 0.00090558 3.3 0.0009055000000000001 3.3 0.0009056 0 0.00090552 0 0.00090562 3.3 0.00090554 3.3 0.00090564 0 0.00090556 0 0.00090566 3.3 0.00090558 3.3 0.00090568 0 0.0009056 0 0.0009057 3.3 0.00090562 3.3 0.0009057199999999999 0 0.00090564 0 0.0009057399999999999 3.3 0.0009056600000000001 3.3 0.00090576 0 0.0009056800000000001 0 0.00090578 3.3 0.0009057000000000001 3.3 0.0009058 0 0.00090572 0 0.00090582 3.3 0.00090574 3.3 0.00090584 0 0.00090576 0 0.00090586 3.3 0.00090578 3.3 0.00090588 0 0.0009058 0 0.0009059 3.3 0.00090582 3.3 0.00090592 0 0.00090584 0 0.0009059399999999999 3.3 0.0009058600000000001 3.3 0.00090596 0 0.0009058800000000001 0 0.00090598 3.3 0.0009059000000000001 3.3 0.000906 0 0.0009059200000000001 0 0.00090602 3.3 0.00090594 3.3 0.00090604 0 0.00090596 0 0.00090606 3.3 0.00090598 3.3 0.00090608 0 0.000906 0 0.0009061 3.3 0.00090602 3.3 0.00090612 0 0.00090604 0 0.0009061399999999999 3.3 0.00090606 3.3 0.0009061599999999999 0 0.0009060800000000001 0 0.00090618 3.3 0.0009061000000000001 3.3 0.0009062 0 0.0009061200000000001 0 0.00090622 3.3 0.00090614 3.3 0.00090624 0 0.00090616 0 0.00090626 3.3 0.00090618 3.3 0.00090628 0 0.0009062 0 0.0009063 3.3 0.00090622 3.3 0.00090632 0 0.00090624 0 0.0009063399999999999 3.3 0.00090626 3.3 0.0009063599999999999 0 0.0009062800000000001 0 0.00090638 3.3 0.0009063000000000001 3.3 0.0009064 0 0.0009063200000000001 0 0.00090642 3.3 0.00090634 3.3 0.00090644 0 0.00090636 0 0.00090646 3.3 0.00090638 3.3 0.00090648 0 0.0009064 0 0.0009065 3.3 0.00090642 3.3 0.00090652 0 0.00090644 0 0.00090654 3.3 0.00090646 3.3 0.0009065599999999999 0 0.00090648 0 0.0009065799999999999 3.3 0.0009065000000000001 3.3 0.0009066 0 0.0009065200000000001 0 0.00090662 3.3 0.0009065400000000001 3.3 0.00090664 0 0.00090656 0 0.00090666 3.3 0.00090658 3.3 0.00090668 0 0.0009066 0 0.0009067 3.3 0.00090662 3.3 0.00090672 0 0.00090664 0 0.00090674 3.3 0.00090666 3.3 0.0009067599999999999 0 0.00090668 0 0.0009067799999999999 3.3 0.0009067000000000001 3.3 0.0009068 0 0.0009067200000000001 0 0.00090682 3.3 0.0009067400000000001 3.3 0.00090684 0 0.00090676 0 0.00090686 3.3 0.00090678 3.3 0.00090688 0 0.0009068 0 0.0009069 3.3 0.00090682 3.3 0.00090692 0 0.00090684 0 0.00090694 3.3 0.00090686 3.3 0.00090696 0 0.00090688 0 0.0009069799999999999 3.3 0.0009069 3.3 0.0009069999999999999 0 0.0009069200000000001 0 0.00090702 3.3 0.0009069400000000001 3.3 0.00090704 0 0.0009069600000000001 0 0.00090706 3.3 0.00090698 3.3 0.00090708 0 0.000907 0 0.0009071 3.3 0.00090702 3.3 0.00090712 0 0.00090704 0 0.00090714 3.3 0.00090706 3.3 0.00090716 0 0.00090708 0 0.0009071799999999999 3.3 0.0009071 3.3 0.0009071999999999999 0 0.0009071200000000001 0 0.00090722 3.3 0.0009071400000000001 3.3 0.00090724 0 0.0009071600000000001 0 0.00090726 3.3 0.00090718 3.3 0.00090728 0 0.0009072 0 0.0009073 3.3 0.00090722 3.3 0.00090732 0 0.00090724 0 0.00090734 3.3 0.00090726 3.3 0.00090736 0 0.00090728 0 0.00090738 3.3 0.0009073 3.3 0.0009073999999999999 0 0.00090732 0 0.0009074199999999999 3.3 0.0009073400000000001 3.3 0.00090744 0 0.0009073600000000001 0 0.00090746 3.3 0.0009073800000000001 3.3 0.00090748 0 0.0009074 0 0.0009075 3.3 0.00090742 3.3 0.00090752 0 0.00090744 0 0.00090754 3.3 0.00090746 3.3 0.00090756 0 0.00090748 0 0.00090758 3.3 0.0009075 3.3 0.0009075999999999999 0 0.00090752 0 0.0009076199999999999 3.3 0.0009075400000000001 3.3 0.00090764 0 0.0009075600000000001 0 0.00090766 3.3 0.0009075800000000001 3.3 0.00090768 0 0.0009076 0 0.0009077 3.3 0.00090762 3.3 0.00090772 0 0.00090764 0 0.00090774 3.3 0.00090766 3.3 0.00090776 0 0.00090768 0 0.00090778 3.3 0.0009077 3.3 0.0009078 0 0.00090772 0 0.0009078199999999999 3.3 0.0009077400000000001 3.3 0.00090784 0 0.0009077600000000001 0 0.00090786 3.3 0.0009077800000000001 3.3 0.00090788 0 0.0009078000000000001 0 0.0009079 3.3 0.00090782 3.3 0.00090792 0 0.00090784 0 0.00090794 3.3 0.00090786 3.3 0.00090796 0 0.00090788 0 0.00090798 3.3 0.0009079 3.3 0.000908 0 0.00090792 0 0.0009080199999999999 3.3 0.00090794 3.3 0.0009080399999999999 0 0.0009079600000000001 0 0.00090806 3.3 0.0009079800000000001 3.3 0.00090808 0 0.0009080000000000001 0 0.0009081 3.3 0.00090802 3.3 0.00090812 0 0.00090804 0 0.00090814 3.3 0.00090806 3.3 0.00090816 0 0.00090808 0 0.00090818 3.3 0.0009081 3.3 0.0009082 0 0.00090812 0 0.00090822 3.3 0.00090814 3.3 0.0009082399999999999 0 0.0009081600000000001 0 0.00090826 3.3 0.0009081800000000001 3.3 0.00090828 0 0.0009082000000000001 0 0.0009083 3.3 0.0009082200000000001 3.3 0.00090832 0 0.00090824 0 0.00090834 3.3 0.00090826 3.3 0.00090836 0 0.00090828 0 0.00090838 3.3 0.0009083 3.3 0.0009084 0 0.00090832 0 0.00090842 3.3 0.00090834 3.3 0.0009084399999999999 0 0.00090836 0 0.0009084599999999999 3.3 0.0009083800000000001 3.3 0.00090848 0 0.0009084000000000001 0 0.0009085 3.3 0.0009084200000000001 3.3 0.00090852 0 0.00090844 0 0.00090854 3.3 0.00090846 3.3 0.00090856 0 0.00090848 0 0.00090858 3.3 0.0009085 3.3 0.0009086 0 0.00090852 0 0.00090862 3.3 0.00090854 3.3 0.00090864 0 0.00090856 0 0.0009086599999999999 3.3 0.0009085800000000001 3.3 0.00090868 0 0.0009086000000000001 0 0.0009087 3.3 0.0009086200000000001 3.3 0.00090872 0 0.0009086400000000001 0 0.00090874 3.3 0.00090866 3.3 0.00090876 0 0.00090868 0 0.00090878 3.3 0.0009087 3.3 0.0009088 0 0.00090872 0 0.00090882 3.3 0.00090874 3.3 0.00090884 0 0.00090876 0 0.0009088599999999999 3.3 0.00090878 3.3 0.0009088799999999999 0 0.0009088000000000001 0 0.0009089 3.3 0.0009088200000000001 3.3 0.00090892 0 0.0009088400000000001 0 0.00090894 3.3 0.00090886 3.3 0.00090896 0 0.00090888 0 0.00090898 3.3 0.0009089 3.3 0.000909 0 0.00090892 0 0.00090902 3.3 0.00090894 3.3 0.00090904 0 0.00090896 0 0.00090906 3.3 0.00090898 3.3 0.0009090799999999999 0 0.0009090000000000001 0 0.0009091 3.3 0.0009090200000000001 3.3 0.00090912 0 0.0009090400000000001 0 0.00090914 3.3 0.0009090600000000001 3.3 0.00090916 0 0.00090908 0 0.00090918 3.3 0.0009091 3.3 0.0009092 0 0.00090912 0 0.00090922 3.3 0.00090914 3.3 0.00090924 0 0.00090916 0 0.00090926 3.3 0.00090918 3.3 0.0009092799999999999 0 0.0009092 0 0.0009092999999999999 3.3 0.0009092200000000001 3.3 0.00090932 0 0.0009092400000000001 0 0.00090934 3.3 0.0009092600000000001 3.3 0.00090936 0 0.00090928 0 0.00090938 3.3 0.0009093 3.3 0.0009094 0 0.00090932 0 0.00090942 3.3 0.00090934 3.3 0.00090944 0 0.00090936 0 0.00090946 3.3 0.00090938 3.3 0.0009094799999999999 0 0.0009094 0 0.0009094999999999999 3.3 0.0009094200000000001 3.3 0.00090952 0 0.0009094400000000001 0 0.00090954 3.3 0.0009094600000000001 3.3 0.00090956 0 0.00090948 0 0.00090958 3.3 0.0009095 3.3 0.0009096 0 0.00090952 0 0.00090962 3.3 0.00090954 3.3 0.00090964 0 0.00090956 0 0.00090966 3.3 0.00090958 3.3 0.00090968 0 0.0009096 0 0.0009096999999999999 3.3 0.00090962 3.3 0.0009097199999999999 0 0.0009096400000000001 0 0.00090974 3.3 0.0009096600000000001 3.3 0.00090976 0 0.0009096800000000001 0 0.00090978 3.3 0.0009097 3.3 0.0009098 0 0.00090972 0 0.00090982 3.3 0.00090974 3.3 0.00090984 0 0.00090976 0 0.00090986 3.3 0.00090978 3.3 0.00090988 0 0.0009098 0 0.0009098999999999999 3.3 0.00090982 3.3 0.0009099199999999999 0 0.0009098400000000001 0 0.00090994 3.3 0.0009098600000000001 3.3 0.00090996 0 0.0009098800000000001 0 0.00090998 3.3 0.0009099 3.3 0.00091 0 0.00090992 0 0.00091002 3.3 0.00090994 3.3 0.00091004 0 0.00090996 0 0.00091006 3.3 0.00090998 3.3 0.00091008 0 0.00091 0 0.0009101 3.3 0.00091002 3.3 0.0009101199999999999 0 0.00091004 0 0.0009101399999999999 3.3 0.0009100600000000001 3.3 0.00091016 0 0.0009100800000000001 0 0.00091018 3.3 0.0009101000000000001 3.3 0.0009102 0 0.00091012 0 0.00091022 3.3 0.00091014 3.3 0.00091024 0 0.00091016 0 0.00091026 3.3 0.00091018 3.3 0.00091028 0 0.0009102 0 0.0009103 3.3 0.00091022 3.3 0.0009103199999999999 0 0.00091024 0 0.0009103399999999999 3.3 0.0009102600000000001 3.3 0.00091036 0 0.0009102800000000001 0 0.00091038 3.3 0.0009103000000000001 3.3 0.0009104 0 0.00091032 0 0.00091042 3.3 0.00091034 3.3 0.00091044 0 0.00091036 0 0.00091046 3.3 0.00091038 3.3 0.00091048 0 0.0009104 0 0.0009105 3.3 0.00091042 3.3 0.00091052 0 0.00091044 0 0.0009105399999999999 3.3 0.00091046 3.3 0.0009105599999999999 0 0.0009104800000000001 0 0.00091058 3.3 0.0009105000000000001 3.3 0.0009106 0 0.0009105200000000001 0 0.00091062 3.3 0.00091054 3.3 0.00091064 0 0.00091056 0 0.00091066 3.3 0.00091058 3.3 0.00091068 0 0.0009106 0 0.0009107 3.3 0.00091062 3.3 0.00091072 0 0.00091064 0 0.0009107399999999999 3.3 0.00091066 3.3 0.0009107599999999999 0 0.0009106800000000001 0 0.00091078 3.3 0.0009107000000000001 3.3 0.0009108 0 0.0009107200000000001 0 0.00091082 3.3 0.00091074 3.3 0.00091084 0 0.00091076 0 0.00091086 3.3 0.00091078 3.3 0.00091088 0 0.0009108 0 0.0009109 3.3 0.00091082 3.3 0.00091092 0 0.00091084 0 0.00091094 3.3 0.00091086 3.3 0.0009109599999999999 0 0.00091088 0 0.0009109799999999999 3.3 0.0009109000000000001 3.3 0.000911 0 0.0009109200000000001 0 0.00091102 3.3 0.0009109400000000001 3.3 0.00091104 0 0.00091096 0 0.00091106 3.3 0.00091098 3.3 0.00091108 0 0.000911 0 0.0009111 3.3 0.00091102 3.3 0.00091112 0 0.00091104 0 0.00091114 3.3 0.00091106 3.3 0.0009111599999999999 0 0.00091108 0 0.0009111799999999999 3.3 0.0009111000000000001 3.3 0.0009112 0 0.0009111200000000001 0 0.00091122 3.3 0.0009111400000000001 3.3 0.00091124 0 0.00091116 0 0.00091126 3.3 0.00091118 3.3 0.00091128 0 0.0009112 0 0.0009113 3.3 0.00091122 3.3 0.00091132 0 0.00091124 0 0.00091134 3.3 0.00091126 3.3 0.00091136 0 0.00091128 0 0.0009113799999999999 3.3 0.0009113000000000001 3.3 0.0009114 0 0.0009113200000000001 0 0.00091142 3.3 0.0009113400000000001 3.3 0.00091144 0 0.0009113600000000001 0 0.00091146 3.3 0.00091138 3.3 0.00091148 0 0.0009114 0 0.0009115 3.3 0.00091142 3.3 0.00091152 0 0.00091144 0 0.00091154 3.3 0.00091146 3.3 0.00091156 0 0.00091148 0 0.0009115799999999999 3.3 0.0009115 3.3 0.0009115999999999999 0 0.0009115200000000001 0 0.00091162 3.3 0.0009115400000000001 3.3 0.00091164 0 0.0009115600000000001 0 0.00091166 3.3 0.00091158 3.3 0.00091168 0 0.0009116 0 0.0009117 3.3 0.00091162 3.3 0.00091172 0 0.00091164 0 0.00091174 3.3 0.00091166 3.3 0.00091176 0 0.00091168 0 0.00091178 3.3 0.0009117 3.3 0.0009117999999999999 0 0.0009117200000000001 0 0.00091182 3.3 0.0009117400000000001 3.3 0.00091184 0 0.0009117600000000001 0 0.00091186 3.3 0.0009117800000000001 3.3 0.00091188 0 0.0009118 0 0.0009119 3.3 0.00091182 3.3 0.00091192 0 0.00091184 0 0.00091194 3.3 0.00091186 3.3 0.00091196 0 0.00091188 0 0.00091198 3.3 0.0009119 3.3 0.0009119999999999999 0 0.00091192 0 0.0009120199999999999 3.3 0.0009119400000000001 3.3 0.00091204 0 0.0009119600000000001 0 0.00091206 3.3 0.0009119800000000001 3.3 0.00091208 0 0.000912 0 0.0009121 3.3 0.00091202 3.3 0.00091212 0 0.00091204 0 0.00091214 3.3 0.00091206 3.3 0.00091216 0 0.00091208 0 0.00091218 3.3 0.0009121 3.3 0.0009122 0 0.00091212 0 0.0009122199999999999 3.3 0.0009121400000000001 3.3 0.00091224 0 0.0009121600000000001 0 0.00091226 3.3 0.0009121800000000001 3.3 0.00091228 0 0.0009122000000000001 0 0.0009123 3.3 0.00091222 3.3 0.00091232 0 0.00091224 0 0.00091234 3.3 0.00091226 3.3 0.00091236 0 0.00091228 0 0.00091238 3.3 0.0009123 3.3 0.0009124 0 0.00091232 0 0.0009124199999999999 3.3 0.00091234 3.3 0.0009124399999999999 0 0.0009123600000000001 0 0.00091246 3.3 0.0009123800000000001 3.3 0.00091248 0 0.0009124000000000001 0 0.0009125 3.3 0.00091242 3.3 0.00091252 0 0.00091244 0 0.00091254 3.3 0.00091246 3.3 0.00091256 0 0.00091248 0 0.00091258 3.3 0.0009125 3.3 0.0009126 0 0.00091252 0 0.00091262 3.3 0.00091254 3.3 0.0009126399999999999 0 0.0009125600000000001 0 0.00091266 3.3 0.0009125800000000001 3.3 0.00091268 0 0.0009126000000000001 0 0.0009127 3.3 0.0009126200000000001 3.3 0.00091272 0 0.00091264 0 0.00091274 3.3 0.00091266 3.3 0.00091276 0 0.00091268 0 0.00091278 3.3 0.0009127 3.3 0.0009128 0 0.00091272 0 0.00091282 3.3 0.00091274 3.3 0.0009128399999999999 0 0.00091276 0 0.0009128599999999999 3.3 0.0009127800000000001 3.3 0.00091288 0 0.0009128000000000001 0 0.0009129 3.3 0.0009128200000000001 3.3 0.00091292 0 0.00091284 0 0.00091294 3.3 0.00091286 3.3 0.00091296 0 0.00091288 0 0.00091298 3.3 0.0009129 3.3 0.000913 0 0.00091292 0 0.00091302 3.3 0.00091294 3.3 0.0009130399999999999 0 0.00091296 0 0.0009130599999999999 3.3 0.0009129800000000001 3.3 0.00091308 0 0.0009130000000000001 0 0.0009131 3.3 0.0009130200000000001 3.3 0.00091312 0 0.00091304 0 0.00091314 3.3 0.00091306 3.3 0.00091316 0 0.00091308 0 0.00091318 3.3 0.0009131 3.3 0.0009132 0 0.00091312 0 0.00091322 3.3 0.00091314 3.3 0.00091324 0 0.00091316 0 0.0009132599999999999 3.3 0.00091318 3.3 0.0009132799999999999 0 0.0009132000000000001 0 0.0009133 3.3 0.0009132200000000001 3.3 0.00091332 0 0.0009132400000000001 0 0.00091334 3.3 0.00091326 3.3 0.00091336 0 0.00091328 0 0.00091338 3.3 0.0009133 3.3 0.0009134 0 0.00091332 0 0.00091342 3.3 0.00091334 3.3 0.00091344 0 0.00091336 0 0.0009134599999999999 3.3 0.00091338 3.3 0.0009134799999999999 0 0.0009134000000000001 0 0.0009135 3.3 0.0009134200000000001 3.3 0.00091352 0 0.0009134400000000001 0 0.00091354 3.3 0.00091346 3.3 0.00091356 0 0.00091348 0 0.00091358 3.3 0.0009135 3.3 0.0009136 0 0.00091352 0 0.00091362 3.3 0.00091354 3.3 0.00091364 0 0.00091356 0 0.00091366 3.3 0.00091358 3.3 0.0009136799999999999 0 0.0009136 0 0.0009136999999999999 3.3 0.0009136200000000001 3.3 0.00091372 0 0.0009136400000000001 0 0.00091374 3.3 0.0009136600000000001 3.3 0.00091376 0 0.00091368 0 0.00091378 3.3 0.0009137 3.3 0.0009138 0 0.00091372 0 0.00091382 3.3 0.00091374 3.3 0.00091384 0 0.00091376 0 0.00091386 3.3 0.00091378 3.3 0.0009138799999999999 0 0.0009138 0 0.0009138999999999999 3.3 0.0009138200000000001 3.3 0.00091392 0 0.0009138400000000001 0 0.00091394 3.3 0.0009138600000000001 3.3 0.00091396 0 0.00091388 0 0.00091398 3.3 0.0009139 3.3 0.000914 0 0.00091392 0 0.00091402 3.3 0.00091394 3.3 0.00091404 0 0.00091396 0 0.00091406 3.3 0.00091398 3.3 0.00091408 0 0.000914 0 0.0009140999999999999 3.3 0.00091402 3.3 0.0009141199999999999 0 0.0009140400000000001 0 0.00091414 3.3 0.0009140600000000001 3.3 0.00091416 0 0.0009140800000000001 0 0.00091418 3.3 0.0009141 3.3 0.0009142 0 0.00091412 0 0.00091422 3.3 0.00091414 3.3 0.00091424 0 0.00091416 0 0.00091426 3.3 0.00091418 3.3 0.00091428 0 0.0009142 0 0.0009142999999999999 3.3 0.00091422 3.3 0.0009143199999999999 0 0.0009142400000000001 0 0.00091434 3.3 0.0009142600000000001 3.3 0.00091436 0 0.0009142800000000001 0 0.00091438 3.3 0.0009143 3.3 0.0009144 0 0.00091432 0 0.00091442 3.3 0.00091434 3.3 0.00091444 0 0.00091436 0 0.00091446 3.3 0.00091438 3.3 0.00091448 0 0.0009144 0 0.0009145 3.3 0.00091442 3.3 0.0009145199999999999 0 0.00091444 0 0.0009145399999999999 3.3 0.0009144600000000001 3.3 0.00091456 0 0.0009144800000000001 0 0.00091458 3.3 0.0009145000000000001 3.3 0.0009146 0 0.00091452 0 0.00091462 3.3 0.00091454 3.3 0.00091464 0 0.00091456 0 0.00091466 3.3 0.00091458 3.3 0.00091468 0 0.0009146 0 0.0009147 3.3 0.00091462 3.3 0.0009147199999999999 0 0.00091464 0 0.0009147399999999999 3.3 0.0009146600000000001 3.3 0.00091476 0 0.0009146800000000001 0 0.00091478 3.3 0.0009147000000000001 3.3 0.0009148 0 0.00091472 0 0.00091482 3.3 0.00091474 3.3 0.00091484 0 0.00091476 0 0.00091486 3.3 0.00091478 3.3 0.00091488 0 0.0009148 0 0.0009149 3.3 0.00091482 3.3 0.00091492 0 0.00091484 0 0.0009149399999999999 3.3 0.0009148600000000001 3.3 0.00091496 0 0.0009148800000000001 0 0.00091498 3.3 0.0009149000000000001 3.3 0.000915 0 0.0009149200000000001 0 0.00091502 3.3 0.00091494 3.3 0.00091504 0 0.00091496 0 0.00091506 3.3 0.00091498 3.3 0.00091508 0 0.000915 0 0.0009151 3.3 0.00091502 3.3 0.00091512 0 0.00091504 0 0.0009151399999999999 3.3 0.00091506 3.3 0.0009151599999999999 0 0.0009150800000000001 0 0.00091518 3.3 0.0009151000000000001 3.3 0.0009152 0 0.0009151200000000001 0 0.00091522 3.3 0.00091514 3.3 0.00091524 0 0.00091516 0 0.00091526 3.3 0.00091518 3.3 0.00091528 0 0.0009152 0 0.0009153 3.3 0.00091522 3.3 0.00091532 0 0.00091524 0 0.00091534 3.3 0.00091526 3.3 0.0009153599999999999 0 0.0009152800000000001 0 0.00091538 3.3 0.0009153000000000001 3.3 0.0009154 0 0.0009153200000000001 0 0.00091542 3.3 0.0009153400000000001 3.3 0.00091544 0 0.00091536 0 0.00091546 3.3 0.00091538 3.3 0.00091548 0 0.0009154 0 0.0009155 3.3 0.00091542 3.3 0.00091552 0 0.00091544 0 0.00091554 3.3 0.00091546 3.3 0.0009155599999999999 0 0.00091548 0 0.0009155799999999999 3.3 0.0009155000000000001 3.3 0.0009156 0 0.0009155200000000001 0 0.00091562 3.3 0.0009155400000000001 3.3 0.00091564 0 0.00091556 0 0.00091566 3.3 0.00091558 3.3 0.00091568 0 0.0009156 0 0.0009157 3.3 0.00091562 3.3 0.00091572 0 0.00091564 0 0.00091574 3.3 0.00091566 3.3 0.00091576 0 0.00091568 0 0.0009157799999999999 3.3 0.0009157000000000001 3.3 0.0009158 0 0.0009157200000000001 0 0.00091582 3.3 0.0009157400000000001 3.3 0.00091584 0 0.0009157600000000001 0 0.00091586 3.3 0.00091578 3.3 0.00091588 0 0.0009158 0 0.0009159 3.3 0.00091582 3.3 0.00091592 0 0.00091584 0 0.00091594 3.3 0.00091586 3.3 0.00091596 0 0.00091588 0 0.0009159799999999999 3.3 0.0009159 3.3 0.0009159999999999999 0 0.0009159200000000001 0 0.00091602 3.3 0.0009159400000000001 3.3 0.00091604 0 0.0009159600000000001 0 0.00091606 3.3 0.00091598 3.3 0.00091608 0 0.000916 0 0.0009161 3.3 0.00091602 3.3 0.00091612 0 0.00091604 0 0.00091614 3.3 0.00091606 3.3 0.00091616 0 0.00091608 0 0.00091618 3.3 0.0009161 3.3 0.0009161999999999999 0 0.0009161200000000001 0 0.00091622 3.3 0.0009161400000000001 3.3 0.00091624 0 0.0009161600000000001 0 0.00091626 3.3 0.0009161800000000001 3.3 0.00091628 0 0.0009162 0 0.0009163 3.3 0.00091622 3.3 0.00091632 0 0.00091624 0 0.00091634 3.3 0.00091626 3.3 0.00091636 0 0.00091628 0 0.00091638 3.3 0.0009163 3.3 0.0009163999999999999 0 0.00091632 0 0.0009164199999999999 3.3 0.0009163400000000001 3.3 0.00091644 0 0.0009163600000000001 0 0.00091646 3.3 0.0009163800000000001 3.3 0.00091648 0 0.0009164 0 0.0009165 3.3 0.00091642 3.3 0.00091652 0 0.00091644 0 0.00091654 3.3 0.00091646 3.3 0.00091656 0 0.00091648 0 0.00091658 3.3 0.0009165 3.3 0.0009165999999999999 0 0.00091652 0 0.0009166199999999999 3.3 0.0009165400000000001 3.3 0.00091664 0 0.0009165600000000001 0 0.00091666 3.3 0.0009165800000000001 3.3 0.00091668 0 0.0009166 0 0.0009167 3.3 0.00091662 3.3 0.00091672 0 0.00091664 0 0.00091674 3.3 0.00091666 3.3 0.00091676 0 0.00091668 0 0.00091678 3.3 0.0009167 3.3 0.0009168 0 0.00091672 0 0.0009168199999999999 3.3 0.00091674 3.3 0.0009168399999999999 0 0.0009167600000000001 0 0.00091686 3.3 0.0009167800000000001 3.3 0.00091688 0 0.0009168000000000001 0 0.0009169 3.3 0.00091682 3.3 0.00091692 0 0.00091684 0 0.00091694 3.3 0.00091686 3.3 0.00091696 0 0.00091688 0 0.00091698 3.3 0.0009169 3.3 0.000917 0 0.00091692 0 0.0009170199999999999 3.3 0.00091694 3.3 0.0009170399999999999 0 0.0009169600000000001 0 0.00091706 3.3 0.0009169800000000001 3.3 0.00091708 0 0.0009170000000000001 0 0.0009171 3.3 0.00091702 3.3 0.00091712 0 0.00091704 0 0.00091714 3.3 0.00091706 3.3 0.00091716 0 0.00091708 0 0.00091718 3.3 0.0009171 3.3 0.0009172 0 0.00091712 0 0.00091722 3.3 0.00091714 3.3 0.0009172399999999999 0 0.00091716 0 0.0009172599999999999 3.3 0.0009171800000000001 3.3 0.00091728 0 0.0009172000000000001 0 0.0009173 3.3 0.0009172200000000001 3.3 0.00091732 0 0.00091724 0 0.00091734 3.3 0.00091726 3.3 0.00091736 0 0.00091728 0 0.00091738 3.3 0.0009173 3.3 0.0009174 0 0.00091732 0 0.00091742 3.3 0.00091734 3.3 0.0009174399999999999 0 0.00091736 0 0.0009174599999999999 3.3 0.0009173800000000001 3.3 0.00091748 0 0.0009174000000000001 0 0.0009175 3.3 0.0009174200000000001 3.3 0.00091752 0 0.00091744 0 0.00091754 3.3 0.00091746 3.3 0.00091756 0 0.00091748 0 0.00091758 3.3 0.0009175 3.3 0.0009176 0 0.00091752 0 0.00091762 3.3 0.00091754 3.3 0.00091764 0 0.00091756 0 0.0009176599999999999 3.3 0.00091758 3.3 0.0009176799999999999 0 0.0009176000000000001 0 0.0009177 3.3 0.0009176200000000001 3.3 0.00091772 0 0.0009176400000000001 0 0.00091774 3.3 0.00091766 3.3 0.00091776 0 0.00091768 0 0.00091778 3.3 0.0009177 3.3 0.0009178 0 0.00091772 0 0.00091782 3.3 0.00091774 3.3 0.00091784 0 0.00091776 0 0.0009178599999999999 3.3 0.00091778 3.3 0.0009178799999999999 0 0.0009178000000000001 0 0.0009179 3.3 0.0009178200000000001 3.3 0.00091792 0 0.0009178400000000001 0 0.00091794 3.3 0.00091786 3.3 0.00091796 0 0.00091788 0 0.00091798 3.3 0.0009179 3.3 0.000918 0 0.00091792 0 0.00091802 3.3 0.00091794 3.3 0.00091804 0 0.00091796 0 0.00091806 3.3 0.00091798 3.3 0.0009180799999999999 0 0.000918 0 0.0009180999999999999 3.3 0.0009180200000000001 3.3 0.00091812 0 0.0009180400000000001 0 0.00091814 3.3 0.0009180600000000001 3.3 0.00091816 0 0.00091808 0 0.00091818 3.3 0.0009181 3.3 0.0009182 0 0.00091812 0 0.00091822 3.3 0.00091814 3.3 0.00091824 0 0.00091816 0 0.00091826 3.3 0.00091818 3.3 0.0009182799999999999 0 0.0009182 0 0.0009182999999999999 3.3 0.0009182200000000001 3.3 0.00091832 0 0.0009182400000000001 0 0.00091834 3.3 0.0009182600000000001 3.3 0.00091836 0 0.00091828 0 0.00091838 3.3 0.0009183 3.3 0.0009184 0 0.00091832 0 0.00091842 3.3 0.00091834 3.3 0.00091844 0 0.00091836 0 0.00091846 3.3 0.00091838 3.3 0.00091848 0 0.0009184 0 0.0009184999999999999 3.3 0.0009184200000000001 3.3 0.00091852 0 0.0009184400000000001 0 0.00091854 3.3 0.0009184600000000001 3.3 0.00091856 0 0.0009184800000000001 0 0.00091858 3.3 0.0009185 3.3 0.0009186 0 0.00091852 0 0.00091862 3.3 0.00091854 3.3 0.00091864 0 0.00091856 0 0.00091866 3.3 0.00091858 3.3 0.00091868 0 0.0009186 0 0.0009186999999999999 3.3 0.00091862 3.3 0.0009187199999999999 0 0.0009186400000000001 0 0.00091874 3.3 0.0009186600000000001 3.3 0.00091876 0 0.0009186800000000001 0 0.00091878 3.3 0.0009187 3.3 0.0009188 0 0.00091872 0 0.00091882 3.3 0.00091874 3.3 0.00091884 0 0.00091876 0 0.00091886 3.3 0.00091878 3.3 0.00091888 0 0.0009188 0 0.0009189 3.3 0.00091882 3.3 0.0009189199999999999 0 0.0009188400000000001 0 0.00091894 3.3 0.0009188600000000001 3.3 0.00091896 0 0.0009188800000000001 0 0.00091898 3.3 0.0009189000000000001 3.3 0.000919 0 0.00091892 0 0.00091902 3.3 0.00091894 3.3 0.00091904 0 0.00091896 0 0.00091906 3.3 0.00091898 3.3 0.00091908 0 0.000919 0 0.0009191 3.3 0.00091902 3.3 0.0009191199999999999 0 0.00091904 0 0.0009191399999999999 3.3 0.0009190600000000001 3.3 0.00091916 0 0.0009190800000000001 0 0.00091918 3.3 0.0009191000000000001 3.3 0.0009192 0 0.00091912 0 0.00091922 3.3 0.00091914 3.3 0.00091924 0 0.00091916 0 0.00091926 3.3 0.00091918 3.3 0.00091928 0 0.0009192 0 0.0009193 3.3 0.00091922 3.3 0.00091932 0 0.00091924 0 0.0009193399999999999 3.3 0.0009192600000000001 3.3 0.00091936 0 0.0009192800000000001 0 0.00091938 3.3 0.0009193000000000001 3.3 0.0009194 0 0.0009193200000000001 0 0.00091942 3.3 0.00091934 3.3 0.00091944 0 0.00091936 0 0.00091946 3.3 0.00091938 3.3 0.00091948 0 0.0009194 0 0.0009195 3.3 0.00091942 3.3 0.00091952 0 0.00091944 0 0.0009195399999999999 3.3 0.00091946 3.3 0.0009195599999999999 0 0.0009194800000000001 0 0.00091958 3.3 0.0009195000000000001 3.3 0.0009196 0 0.0009195200000000001 0 0.00091962 3.3 0.00091954 3.3 0.00091964 0 0.00091956 0 0.00091966 3.3 0.00091958 3.3 0.00091968 0 0.0009196 0 0.0009197 3.3 0.00091962 3.3 0.00091972 0 0.00091964 0 0.0009197399999999999 3.3 0.00091966 3.3 0.0009197599999999999 0 0.0009196800000000001 0 0.00091978 3.3 0.0009197000000000001 3.3 0.0009198 0 0.0009197200000000001 0 0.00091982 3.3 0.00091974 3.3 0.00091984 0 0.00091976 0 0.00091986 3.3 0.00091978 3.3 0.00091988 0 0.0009198 0 0.0009199 3.3 0.00091982 3.3 0.00091992 0 0.00091984 0 0.00091994 3.3 0.00091986 3.3 0.0009199599999999999 0 0.00091988 0 0.0009199799999999999 3.3 0.0009199000000000001 3.3 0.00092 0 0.0009199200000000001 0 0.00092002 3.3 0.0009199400000000001 3.3 0.00092004 0 0.00091996 0 0.00092006 3.3 0.00091998 3.3 0.00092008 0 0.00092 0 0.0009201 3.3 0.00092002 3.3 0.00092012 0 0.00092004 0 0.00092014 3.3 0.00092006 3.3 0.0009201599999999999 0 0.00092008 0 0.0009201799999999999 3.3 0.0009201000000000001 3.3 0.0009202 0 0.0009201200000000001 0 0.00092022 3.3 0.0009201400000000001 3.3 0.00092024 0 0.00092016 0 0.00092026 3.3 0.00092018 3.3 0.00092028 0 0.0009202 0 0.0009203 3.3 0.00092022 3.3 0.00092032 0 0.00092024 0 0.00092034 3.3 0.00092026 3.3 0.00092036 0 0.00092028 0 0.0009203799999999999 3.3 0.0009203 3.3 0.0009203999999999999 0 0.0009203200000000001 0 0.00092042 3.3 0.0009203400000000001 3.3 0.00092044 0 0.0009203600000000001 0 0.00092046 3.3 0.00092038 3.3 0.00092048 0 0.0009204 0 0.0009205 3.3 0.00092042 3.3 0.00092052 0 0.00092044 0 0.00092054 3.3 0.00092046 3.3 0.00092056 0 0.00092048 0 0.0009205799999999999 3.3 0.0009205 3.3 0.0009205999999999999 0 0.0009205200000000001 0 0.00092062 3.3 0.0009205400000000001 3.3 0.00092064 0 0.0009205600000000001 0 0.00092066 3.3 0.00092058 3.3 0.00092068 0 0.0009206 0 0.0009207 3.3 0.00092062 3.3 0.00092072 0 0.00092064 0 0.00092074 3.3 0.00092066 3.3 0.00092076 0 0.00092068 0 0.00092078 3.3 0.0009207 3.3 0.0009207999999999999 0 0.00092072 0 0.0009208199999999999 3.3 0.0009207400000000001 3.3 0.00092084 0 0.0009207600000000001 0 0.00092086 3.3 0.0009207800000000001 3.3 0.00092088 0 0.0009208 0 0.0009209 3.3 0.00092082 3.3 0.00092092 0 0.00092084 0 0.00092094 3.3 0.00092086 3.3 0.00092096 0 0.00092088 0 0.00092098 3.3 0.0009209 3.3 0.0009209999999999999 0 0.00092092 0 0.0009210199999999999 3.3 0.0009209400000000001 3.3 0.00092104 0 0.0009209600000000001 0 0.00092106 3.3 0.0009209800000000001 3.3 0.00092108 0 0.000921 0 0.0009211 3.3 0.00092102 3.3 0.00092112 0 0.00092104 0 0.00092114 3.3 0.00092106 3.3 0.00092116 0 0.00092108 0 0.00092118 3.3 0.0009211 3.3 0.0009212 0 0.00092112 0 0.0009212199999999999 3.3 0.00092114 3.3 0.0009212399999999999 0 0.0009211600000000001 0 0.00092126 3.3 0.0009211800000000001 3.3 0.00092128 0 0.0009212000000000001 0 0.0009213 3.3 0.00092122 3.3 0.00092132 0 0.00092124 0 0.00092134 3.3 0.00092126 3.3 0.00092136 0 0.00092128 0 0.00092138 3.3 0.0009213 3.3 0.0009214 0 0.00092132 0 0.0009214199999999999 3.3 0.00092134 3.3 0.0009214399999999999 0 0.0009213600000000001 0 0.00092146 3.3 0.0009213800000000001 3.3 0.00092148 0 0.0009214000000000001 0 0.0009215 3.3 0.00092142 3.3 0.00092152 0 0.00092144 0 0.00092154 3.3 0.00092146 3.3 0.00092156 0 0.00092148 0 0.00092158 3.3 0.0009215 3.3 0.0009216 0 0.00092152 0 0.00092162 3.3 0.00092154 3.3 0.0009216399999999999 0 0.0009215600000000001 0 0.00092166 3.3 0.0009215800000000001 3.3 0.00092168 0 0.0009216000000000001 0 0.0009217 3.3 0.0009216200000000001 3.3 0.00092172 0 0.00092164 0 0.00092174 3.3 0.00092166 3.3 0.00092176 0 0.00092168 0 0.00092178 3.3 0.0009217 3.3 0.0009218 0 0.00092172 0 0.00092182 3.3 0.00092174 3.3 0.0009218399999999999 0 0.00092176 0 0.0009218599999999999 3.3 0.0009217800000000001 3.3 0.00092188 0 0.0009218000000000001 0 0.0009219 3.3 0.0009218200000000001 3.3 0.00092192 0 0.00092184 0 0.00092194 3.3 0.00092186 3.3 0.00092196 0 0.00092188 0 0.00092198 3.3 0.0009219 3.3 0.000922 0 0.00092192 0 0.00092202 3.3 0.00092194 3.3 0.00092204 0 0.00092196 0 0.0009220599999999999 3.3 0.0009219800000000001 3.3 0.00092208 0 0.0009220000000000001 0 0.0009221 3.3 0.0009220200000000001 3.3 0.00092212 0 0.0009220400000000001 0 0.00092214 3.3 0.00092206 3.3 0.00092216 0 0.00092208 0 0.00092218 3.3 0.0009221 3.3 0.0009222 0 0.00092212 0 0.00092222 3.3 0.00092214 3.3 0.00092224 0 0.00092216 0 0.0009222599999999999 3.3 0.00092218 3.3 0.0009222799999999999 0 0.0009222000000000001 0 0.0009223 3.3 0.0009222200000000001 3.3 0.00092232 0 0.0009222400000000001 0 0.00092234 3.3 0.00092226 3.3 0.00092236 0 0.00092228 0 0.00092238 3.3 0.0009223 3.3 0.0009224 0 0.00092232 0 0.00092242 3.3 0.00092234 3.3 0.00092244 0 0.00092236 0 0.00092246 3.3 0.00092238 3.3 0.0009224799999999999 0 0.0009224000000000001 0 0.0009225 3.3 0.0009224200000000001 3.3 0.00092252 0 0.0009224400000000001 0 0.00092254 3.3 0.0009224600000000001 3.3 0.00092256 0 0.00092248 0 0.00092258 3.3 0.0009225 3.3 0.0009226 0 0.00092252 0 0.00092262 3.3 0.00092254 3.3 0.00092264 0 0.00092256 0 0.00092266 3.3 0.00092258 3.3 0.0009226799999999999 0 0.0009226 0 0.0009226999999999999 3.3 0.0009226200000000001 3.3 0.00092272 0 0.0009226400000000001 0 0.00092274 3.3 0.0009226600000000001 3.3 0.00092276 0 0.00092268 0 0.00092278 3.3 0.0009227 3.3 0.0009228 0 0.00092272 0 0.00092282 3.3 0.00092274 3.3 0.00092284 0 0.00092276 0 0.00092286 3.3 0.00092278 3.3 0.00092288 0 0.0009228 0 0.0009228999999999999 3.3 0.0009228200000000001 3.3 0.00092292 0 0.0009228400000000001 0 0.00092294 3.3 0.0009228600000000001 3.3 0.00092296 0 0.0009228800000000001 0 0.00092298 3.3 0.0009229 3.3 0.000923 0 0.00092292 0 0.00092302 3.3 0.00092294 3.3 0.00092304 0 0.00092296 0 0.00092306 3.3 0.00092298 3.3 0.00092308 0 0.000923 0 0.0009230999999999999 3.3 0.00092302 3.3 0.0009231199999999999 0 0.0009230400000000001 0 0.00092314 3.3 0.0009230600000000001 3.3 0.00092316 0 0.0009230800000000001 0 0.00092318 3.3 0.0009231 3.3 0.0009232 0 0.00092312 0 0.00092322 3.3 0.00092314 3.3 0.00092324 0 0.00092316 0 0.00092326 3.3 0.00092318 3.3 0.00092328 0 0.0009232 0 0.0009232999999999999 3.3 0.00092322 3.3 0.0009233199999999999 0 0.0009232400000000001 0 0.00092334 3.3 0.0009232600000000001 3.3 0.00092336 0 0.0009232800000000001 0 0.00092338 3.3 0.0009233 3.3 0.0009234 0 0.00092332 0 0.00092342 3.3 0.00092334 3.3 0.00092344 0 0.00092336 0 0.00092346 3.3 0.00092338 3.3 0.00092348 0 0.0009234 0 0.0009235 3.3 0.00092342 3.3 0.0009235199999999999 0 0.00092344 0 0.0009235399999999999 3.3 0.0009234600000000001 3.3 0.00092356 0 0.0009234800000000001 0 0.00092358 3.3 0.0009235000000000001 3.3 0.0009236 0 0.00092352 0 0.00092362 3.3 0.00092354 3.3 0.00092364 0 0.00092356 0 0.00092366 3.3 0.00092358 3.3 0.00092368 0 0.0009236 0 0.0009237 3.3 0.00092362 3.3 0.0009237199999999999 0 0.00092364 0 0.0009237399999999999 3.3 0.0009236600000000001 3.3 0.00092376 0 0.0009236800000000001 0 0.00092378 3.3 0.0009237000000000001 3.3 0.0009238 0 0.00092372 0 0.00092382 3.3 0.00092374 3.3 0.00092384 0 0.00092376 0 0.00092386 3.3 0.00092378 3.3 0.00092388 0 0.0009238 0 0.0009239 3.3 0.00092382 3.3 0.00092392 0 0.00092384 0 0.0009239399999999999 3.3 0.00092386 3.3 0.0009239599999999999 0 0.0009238800000000001 0 0.00092398 3.3 0.0009239000000000001 3.3 0.000924 0 0.0009239200000000001 0 0.00092402 3.3 0.00092394 3.3 0.00092404 0 0.00092396 0 0.00092406 3.3 0.00092398 3.3 0.00092408 0 0.000924 0 0.0009241 3.3 0.00092402 3.3 0.00092412 0 0.00092404 0 0.0009241399999999999 3.3 0.00092406 3.3 0.0009241599999999999 0 0.0009240800000000001 0 0.00092418 3.3 0.0009241000000000001 3.3 0.0009242 0 0.0009241200000000001 0 0.00092422 3.3 0.00092414 3.3 0.00092424 0 0.00092416 0 0.00092426 3.3 0.00092418 3.3 0.00092428 0 0.0009242 0 0.0009243 3.3 0.00092422 3.3 0.00092432 0 0.00092424 0 0.00092434 3.3 0.00092426 3.3 0.0009243599999999999 0 0.00092428 0 0.0009243799999999999 3.3 0.0009243000000000001 3.3 0.0009244 0 0.0009243200000000001 0 0.00092442 3.3 0.0009243400000000001 3.3 0.00092444 0 0.00092436 0 0.00092446 3.3 0.00092438 3.3 0.00092448 0 0.0009244 0 0.0009245 3.3 0.00092442 3.3 0.00092452 0 0.00092444 0 0.00092454 3.3 0.00092446 3.3 0.0009245599999999999 0 0.00092448 0 0.0009245799999999999 3.3 0.0009245000000000001 3.3 0.0009246 0 0.0009245200000000001 0 0.00092462 3.3 0.0009245400000000001 3.3 0.00092464 0 0.00092456 0 0.00092466 3.3 0.00092458 3.3 0.00092468 0 0.0009246 0 0.0009247 3.3 0.00092462 3.3 0.00092472 0 0.00092464 0 0.00092474 3.3 0.00092466 3.3 0.00092476 0 0.00092468 0 0.0009247799999999999 3.3 0.0009247 3.3 0.0009247999999999999 0 0.0009247200000000001 0 0.00092482 3.3 0.0009247400000000001 3.3 0.00092484 0 0.0009247600000000001 0 0.00092486 3.3 0.00092478 3.3 0.00092488 0 0.0009248 0 0.0009249 3.3 0.00092482 3.3 0.00092492 0 0.00092484 0 0.00092494 3.3 0.00092486 3.3 0.00092496 0 0.00092488 0 0.0009249799999999999 3.3 0.0009249 3.3 0.0009249999999999999 0 0.0009249200000000001 0 0.00092502 3.3 0.0009249400000000001 3.3 0.00092504 0 0.0009249600000000001 0 0.00092506 3.3 0.00092498 3.3 0.00092508 0 0.000925 0 0.0009251 3.3 0.00092502 3.3 0.00092512 0 0.00092504 0 0.00092514 3.3 0.00092506 3.3 0.00092516 0 0.00092508 0 0.00092518 3.3 0.0009251 3.3 0.0009251999999999999 0 0.0009251200000000001 0 0.00092522 3.3 0.0009251400000000001 3.3 0.00092524 0 0.0009251600000000001 0 0.00092526 3.3 0.0009251800000000001 3.3 0.00092528 0 0.0009252 0 0.0009253 3.3 0.00092522 3.3 0.00092532 0 0.00092524 0 0.00092534 3.3 0.00092526 3.3 0.00092536 0 0.00092528 0 0.00092538 3.3 0.0009253 3.3 0.0009253999999999999 0 0.00092532 0 0.0009254199999999999 3.3 0.0009253400000000001 3.3 0.00092544 0 0.0009253600000000001 0 0.00092546 3.3 0.0009253800000000001 3.3 0.00092548 0 0.0009254 0 0.0009255 3.3 0.00092542 3.3 0.00092552 0 0.00092544 0 0.00092554 3.3 0.00092546 3.3 0.00092556 0 0.00092548 0 0.00092558 3.3 0.0009255 3.3 0.0009256 0 0.00092552 0 0.0009256199999999999 3.3 0.0009255400000000001 3.3 0.00092564 0 0.0009255600000000001 0 0.00092566 3.3 0.0009255800000000001 3.3 0.00092568 0 0.0009256000000000001 0 0.0009257 3.3 0.00092562 3.3 0.00092572 0 0.00092564 0 0.00092574 3.3 0.00092566 3.3 0.00092576 0 0.00092568 0 0.00092578 3.3 0.0009257 3.3 0.0009258 0 0.00092572 0 0.0009258199999999999 3.3 0.00092574 3.3 0.0009258399999999999 0 0.0009257600000000001 0 0.00092586 3.3 0.0009257800000000001 3.3 0.00092588 0 0.0009258000000000001 0 0.0009259 3.3 0.00092582 3.3 0.00092592 0 0.00092584 0 0.00092594 3.3 0.00092586 3.3 0.00092596 0 0.00092588 0 0.00092598 3.3 0.0009259 3.3 0.000926 0 0.00092592 0 0.00092602 3.3 0.00092594 3.3 0.0009260399999999999 0 0.0009259600000000001 0 0.00092606 3.3 0.0009259800000000001 3.3 0.00092608 0 0.0009260000000000001 0 0.0009261 3.3 0.0009260200000000001 3.3 0.00092612 0 0.00092604 0 0.00092614 3.3 0.00092606 3.3 0.00092616 0 0.00092608 0 0.00092618 3.3 0.0009261 3.3 0.0009262 0 0.00092612 0 0.00092622 3.3 0.00092614 3.3 0.0009262399999999999 0 0.00092616 0 0.0009262599999999999 3.3 0.0009261800000000001 3.3 0.00092628 0 0.0009262000000000001 0 0.0009263 3.3 0.0009262200000000001 3.3 0.00092632 0 0.00092624 0 0.00092634 3.3 0.00092626 3.3 0.00092636 0 0.00092628 0 0.00092638 3.3 0.0009263 3.3 0.0009264 0 0.00092632 0 0.00092642 3.3 0.00092634 3.3 0.00092644 0 0.00092636 0 0.0009264599999999999 3.3 0.0009263800000000001 3.3 0.00092648 0 0.0009264000000000001 0 0.0009265 3.3 0.0009264200000000001 3.3 0.00092652 0 0.0009264400000000001 0 0.00092654 3.3 0.00092646 3.3 0.00092656 0 0.00092648 0 0.00092658 3.3 0.0009265 3.3 0.0009266 0 0.00092652 0 0.00092662 3.3 0.00092654 3.3 0.00092664 0 0.00092656 0 0.0009266599999999999 3.3 0.00092658 3.3 0.0009266799999999999 0 0.0009266000000000001 0 0.0009267 3.3 0.0009266200000000001 3.3 0.00092672 0 0.0009266400000000001 0 0.00092674 3.3 0.00092666 3.3 0.00092676 0 0.00092668 0 0.00092678 3.3 0.0009267 3.3 0.0009268 0 0.00092672 0 0.00092682 3.3 0.00092674 3.3 0.00092684 0 0.00092676 0 0.0009268599999999999 3.3 0.00092678 3.3 0.0009268799999999999 0 0.0009268000000000001 0 0.0009269 3.3 0.0009268200000000001 3.3 0.00092692 0 0.0009268400000000001 0 0.00092694 3.3 0.00092686 3.3 0.00092696 0 0.00092688 0 0.00092698 3.3 0.0009269 3.3 0.000927 0 0.00092692 0 0.00092702 3.3 0.00092694 3.3 0.00092704 0 0.00092696 0 0.00092706 3.3 0.00092698 3.3 0.0009270799999999999 0 0.000927 0 0.0009270999999999999 3.3 0.0009270200000000001 3.3 0.00092712 0 0.0009270400000000001 0 0.00092714 3.3 0.0009270600000000001 3.3 0.00092716 0 0.00092708 0 0.00092718 3.3 0.0009271 3.3 0.0009272 0 0.00092712 0 0.00092722 3.3 0.00092714 3.3 0.00092724 0 0.00092716 0 0.00092726 3.3 0.00092718 3.3 0.0009272799999999999 0 0.0009272 0 0.0009272999999999999 3.3 0.0009272200000000001 3.3 0.00092732 0 0.0009272400000000001 0 0.00092734 3.3 0.0009272600000000001 3.3 0.00092736 0 0.00092728 0 0.00092738 3.3 0.0009273 3.3 0.0009274 0 0.00092732 0 0.00092742 3.3 0.00092734 3.3 0.00092744 0 0.00092736 0 0.00092746 3.3 0.00092738 3.3 0.00092748 0 0.0009274 0 0.0009274999999999999 3.3 0.00092742 3.3 0.0009275199999999999 0 0.0009274400000000001 0 0.00092754 3.3 0.0009274600000000001 3.3 0.00092756 0 0.0009274800000000001 0 0.00092758 3.3 0.0009275 3.3 0.0009276 0 0.00092752 0 0.00092762 3.3 0.00092754 3.3 0.00092764 0 0.00092756 0 0.00092766 3.3 0.00092758 3.3 0.00092768 0 0.0009276 0 0.0009276999999999999 3.3 0.00092762 3.3 0.0009277199999999999 0 0.0009276400000000001 0 0.00092774 3.3 0.0009276600000000001 3.3 0.00092776 0 0.0009276800000000001 0 0.00092778 3.3 0.0009277 3.3 0.0009278 0 0.00092772 0 0.00092782 3.3 0.00092774 3.3 0.00092784 0 0.00092776 0 0.00092786 3.3 0.00092778 3.3 0.00092788 0 0.0009278 0 0.0009279 3.3 0.00092782 3.3 0.0009279199999999999 0 0.00092784 0 0.0009279399999999999 3.3 0.0009278600000000001 3.3 0.00092796 0 0.0009278800000000001 0 0.00092798 3.3 0.0009279000000000001 3.3 0.000928 0 0.00092792 0 0.00092802 3.3 0.00092794 3.3 0.00092804 0 0.00092796 0 0.00092806 3.3 0.00092798 3.3 0.00092808 0 0.000928 0 0.0009281 3.3 0.00092802 3.3 0.0009281199999999999 0 0.00092804 0 0.0009281399999999999 3.3 0.0009280600000000001 3.3 0.00092816 0 0.0009280800000000001 0 0.00092818 3.3 0.0009281000000000001 3.3 0.0009282 0 0.00092812 0 0.00092822 3.3 0.00092814 3.3 0.00092824 0 0.00092816 0 0.00092826 3.3 0.00092818 3.3 0.00092828 0 0.0009282 0 0.0009283 3.3 0.00092822 3.3 0.00092832 0 0.00092824 0 0.0009283399999999999 3.3 0.00092826 3.3 0.0009283599999999999 0 0.0009282800000000001 0 0.00092838 3.3 0.0009283000000000001 3.3 0.0009284 0 0.0009283200000000001 0 0.00092842 3.3 0.00092834 3.3 0.00092844 0 0.00092836 0 0.00092846 3.3 0.00092838 3.3 0.00092848 0 0.0009284 0 0.0009285 3.3 0.00092842 3.3 0.00092852 0 0.00092844 0 0.0009285399999999999 3.3 0.00092846 3.3 0.0009285599999999999 0 0.0009284800000000001 0 0.00092858 3.3 0.0009285000000000001 3.3 0.0009286 0 0.0009285200000000001 0 0.00092862 3.3 0.00092854 3.3 0.00092864 0 0.00092856 0 0.00092866 3.3 0.00092858 3.3 0.00092868 0 0.0009286 0 0.0009287 3.3 0.00092862 3.3 0.00092872 0 0.00092864 0 0.00092874 3.3 0.00092866 3.3 0.0009287599999999999 0 0.0009286800000000001 0 0.00092878 3.3 0.0009287000000000001 3.3 0.0009288 0 0.0009287200000000001 0 0.00092882 3.3 0.0009287400000000001 3.3 0.00092884 0 0.00092876 0 0.00092886 3.3 0.00092878 3.3 0.00092888 0 0.0009288 0 0.0009289 3.3 0.00092882 3.3 0.00092892 0 0.00092884 0 0.00092894 3.3 0.00092886 3.3 0.0009289599999999999 0 0.00092888 0 0.0009289799999999999 3.3 0.0009289000000000001 3.3 0.000929 0 0.0009289200000000001 0 0.00092902 3.3 0.0009289400000000001 3.3 0.00092904 0 0.00092896 0 0.00092906 3.3 0.00092898 3.3 0.00092908 0 0.000929 0 0.0009291 3.3 0.00092902 3.3 0.00092912 0 0.00092904 0 0.00092914 3.3 0.00092906 3.3 0.00092916 0 0.00092908 0 0.0009291799999999999 3.3 0.0009291000000000001 3.3 0.0009292 0 0.0009291200000000001 0 0.00092922 3.3 0.0009291400000000001 3.3 0.00092924 0 0.0009291600000000001 0 0.00092926 3.3 0.00092918 3.3 0.00092928 0 0.0009292 0 0.0009293 3.3 0.00092922 3.3 0.00092932 0 0.00092924 0 0.00092934 3.3 0.00092926 3.3 0.00092936 0 0.00092928 0 0.0009293799999999999 3.3 0.0009293 3.3 0.0009293999999999999 0 0.0009293200000000001 0 0.00092942 3.3 0.0009293400000000001 3.3 0.00092944 0 0.0009293600000000001 0 0.00092946 3.3 0.00092938 3.3 0.00092948 0 0.0009294 0 0.0009295 3.3 0.00092942 3.3 0.00092952 0 0.00092944 0 0.00092954 3.3 0.00092946 3.3 0.00092956 0 0.00092948 0 0.00092958 3.3 0.0009295 3.3 0.0009295999999999999 0 0.0009295200000000001 0 0.00092962 3.3 0.0009295400000000001 3.3 0.00092964 0 0.0009295600000000001 0 0.00092966 3.3 0.0009295800000000001 3.3 0.00092968 0 0.0009296 0 0.0009297 3.3 0.00092962 3.3 0.00092972 0 0.00092964 0 0.00092974 3.3 0.00092966 3.3 0.00092976 0 0.00092968 0 0.00092978 3.3 0.0009297 3.3 0.0009297999999999999 0 0.00092972 0 0.0009298199999999999 3.3 0.0009297400000000001 3.3 0.00092984 0 0.0009297600000000001 0 0.00092986 3.3 0.0009297800000000001 3.3 0.00092988 0 0.0009298 0 0.0009299 3.3 0.00092982 3.3 0.00092992 0 0.00092984 0 0.00092994 3.3 0.00092986 3.3 0.00092996 0 0.00092988 0 0.00092998 3.3 0.0009299 3.3 0.0009299999999999999 0 0.00092992 0 0.0009300199999999999 3.3 0.0009299400000000001 3.3 0.00093004 0 0.0009299600000000001 0 0.00093006 3.3 0.0009299800000000001 3.3 0.00093008 0 0.00093 0 0.0009301 3.3 0.00093002 3.3 0.00093012 0 0.00093004 0 0.00093014 3.3 0.00093006 3.3 0.00093016 0 0.00093008 0 0.00093018 3.3 0.0009301 3.3 0.0009302 0 0.00093012 0 0.0009302199999999999 3.3 0.00093014 3.3 0.0009302399999999999 0 0.0009301600000000001 0 0.00093026 3.3 0.0009301800000000001 3.3 0.00093028 0 0.0009302000000000001 0 0.0009303 3.3 0.00093022 3.3 0.00093032 0 0.00093024 0 0.00093034 3.3 0.00093026 3.3 0.00093036 0 0.00093028 0 0.00093038 3.3 0.0009303 3.3 0.0009304 0 0.00093032 0 0.0009304199999999999 3.3 0.00093034 3.3 0.0009304399999999999 0 0.0009303600000000001 0 0.00093046 3.3 0.0009303800000000001 3.3 0.00093048 0 0.0009304000000000001 0 0.0009305 3.3 0.00093042 3.3 0.00093052 0 0.00093044 0 0.00093054 3.3 0.00093046 3.3 0.00093056 0 0.00093048 0 0.00093058 3.3 0.0009305 3.3 0.0009306 0 0.00093052 0 0.00093062 3.3 0.00093054 3.3 0.0009306399999999999 0 0.00093056 0 0.0009306599999999999 3.3 0.0009305800000000001 3.3 0.00093068 0 0.0009306000000000001 0 0.0009307 3.3 0.0009306200000000001 3.3 0.00093072 0 0.00093064 0 0.00093074 3.3 0.00093066 3.3 0.00093076 0 0.00093068 0 0.00093078 3.3 0.0009307 3.3 0.0009308 0 0.00093072 0 0.00093082 3.3 0.00093074 3.3 0.0009308399999999999 0 0.00093076 0 0.0009308599999999999 3.3 0.0009307800000000001 3.3 0.00093088 0 0.0009308000000000001 0 0.0009309 3.3 0.0009308200000000001 3.3 0.00093092 0 0.00093084 0 0.00093094 3.3 0.00093086 3.3 0.00093096 0 0.00093088 0 0.00093098 3.3 0.0009309 3.3 0.000931 0 0.00093092 0 0.00093102 3.3 0.00093094 3.3 0.00093104 0 0.00093096 0 0.0009310599999999999 3.3 0.00093098 3.3 0.0009310799999999999 0 0.0009310000000000001 0 0.0009311 3.3 0.0009310200000000001 3.3 0.00093112 0 0.0009310400000000001 0 0.00093114 3.3 0.00093106 3.3 0.00093116 0 0.00093108 0 0.00093118 3.3 0.0009311 3.3 0.0009312 0 0.00093112 0 0.00093122 3.3 0.00093114 3.3 0.00093124 0 0.00093116 0 0.0009312599999999999 3.3 0.00093118 3.3 0.0009312799999999999 0 0.0009312000000000001 0 0.0009313 3.3 0.0009312200000000001 3.3 0.00093132 0 0.0009312400000000001 0 0.00093134 3.3 0.00093126 3.3 0.00093136 0 0.00093128 0 0.00093138 3.3 0.0009313 3.3 0.0009314 0 0.00093132 0 0.00093142 3.3 0.00093134 3.3 0.00093144 0 0.00093136 0 0.00093146 3.3 0.00093138 3.3 0.0009314799999999999 0 0.0009314 0 0.0009314999999999999 3.3 0.0009314200000000001 3.3 0.00093152 0 0.0009314400000000001 0 0.00093154 3.3 0.0009314600000000001 3.3 0.00093156 0 0.00093148 0 0.00093158 3.3 0.0009315 3.3 0.0009316 0 0.00093152 0 0.00093162 3.3 0.00093154 3.3 0.00093164 0 0.00093156 0 0.00093166 3.3 0.00093158 3.3 0.0009316799999999999 0 0.0009316 0 0.0009316999999999999 3.3 0.0009316200000000001 3.3 0.00093172 0 0.0009316400000000001 0 0.00093174 3.3 0.0009316600000000001 3.3 0.00093176 0 0.00093168 0 0.00093178 3.3 0.0009317 3.3 0.0009318 0 0.00093172 0 0.00093182 3.3 0.00093174 3.3 0.00093184 0 0.00093176 0 0.00093186 3.3 0.00093178 3.3 0.00093188 0 0.0009318 0 0.0009318999999999999 3.3 0.00093182 3.3 0.0009319199999999999 0 0.0009318400000000001 0 0.00093194 3.3 0.0009318600000000001 3.3 0.00093196 0 0.0009318800000000001 0 0.00093198 3.3 0.0009319 3.3 0.000932 0 0.00093192 0 0.00093202 3.3 0.00093194 3.3 0.00093204 0 0.00093196 0 0.00093206 3.3 0.00093198 3.3 0.00093208 0 0.000932 0 0.0009320999999999999 3.3 0.00093202 3.3 0.0009321199999999999 0 0.0009320400000000001 0 0.00093214 3.3 0.0009320600000000001 3.3 0.00093216 0 0.0009320800000000001 0 0.00093218 3.3 0.0009321 3.3 0.0009322 0 0.00093212 0 0.00093222 3.3 0.00093214 3.3 0.00093224 0 0.00093216 0 0.00093226 3.3 0.00093218 3.3 0.00093228 0 0.0009322 0 0.0009323 3.3 0.00093222 3.3 0.0009323199999999999 0 0.0009322400000000001 0 0.00093234 3.3 0.0009322600000000001 3.3 0.00093236 0 0.0009322800000000001 0 0.00093238 3.3 0.0009323000000000001 3.3 0.0009324 0 0.00093232 0 0.00093242 3.3 0.00093234 3.3 0.00093244 0 0.00093236 0 0.00093246 3.3 0.00093238 3.3 0.00093248 0 0.0009324 0 0.0009325 3.3 0.00093242 3.3 0.0009325199999999999 0 0.00093244 0 0.0009325399999999999 3.3 0.0009324600000000001 3.3 0.00093256 0 0.0009324800000000001 0 0.00093258 3.3 0.0009325000000000001 3.3 0.0009326 0 0.00093252 0 0.00093262 3.3 0.00093254 3.3 0.00093264 0 0.00093256 0 0.00093266 3.3 0.00093258 3.3 0.00093268 0 0.0009326 0 0.0009327 3.3 0.00093262 3.3 0.00093272 0 0.00093264 0 0.0009327399999999999 3.3 0.0009326600000000001 3.3 0.00093276 0 0.0009326800000000001 0 0.00093278 3.3 0.0009327000000000001 3.3 0.0009328 0 0.0009327200000000001 0 0.00093282 3.3 0.00093274 3.3 0.00093284 0 0.00093276 0 0.00093286 3.3 0.00093278 3.3 0.00093288 0 0.0009328 0 0.0009329 3.3 0.00093282 3.3 0.00093292 0 0.00093284 0 0.0009329399999999999 3.3 0.00093286 3.3 0.0009329599999999999 0 0.0009328800000000001 0 0.00093298 3.3 0.0009329000000000001 3.3 0.000933 0 0.0009329200000000001 0 0.00093302 3.3 0.00093294 3.3 0.00093304 0 0.00093296 0 0.00093306 3.3 0.00093298 3.3 0.00093308 0 0.000933 0 0.0009331 3.3 0.00093302 3.3 0.00093312 0 0.00093304 0 0.00093314 3.3 0.00093306 3.3 0.0009331599999999999 0 0.0009330800000000001 0 0.00093318 3.3 0.0009331000000000001 3.3 0.0009332 0 0.0009331200000000001 0 0.00093322 3.3 0.0009331400000000001 3.3 0.00093324 0 0.00093316 0 0.00093326 3.3 0.00093318 3.3 0.00093328 0 0.0009332 0 0.0009333 3.3 0.00093322 3.3 0.00093332 0 0.00093324 0 0.00093334 3.3 0.00093326 3.3 0.0009333599999999999 0 0.00093328 0 0.0009333799999999999 3.3 0.0009333000000000001 3.3 0.0009334 0 0.0009333200000000001 0 0.00093342 3.3 0.0009333400000000001 3.3 0.00093344 0 0.00093336 0 0.00093346 3.3 0.00093338 3.3 0.00093348 0 0.0009334 0 0.0009335 3.3 0.00093342 3.3 0.00093352 0 0.00093344 0 0.00093354 3.3 0.00093346 3.3 0.0009335599999999999 0 0.00093348 0 0.0009335799999999999 3.3 0.0009335000000000001 3.3 0.0009336 0 0.0009335200000000001 0 0.00093362 3.3 0.0009335400000000001 3.3 0.00093364 0 0.00093356 0 0.00093366 3.3 0.00093358 3.3 0.00093368 0 0.0009336 0 0.0009337 3.3 0.00093362 3.3 0.00093372 0 0.00093364 0 0.00093374 3.3 0.00093366 3.3 0.00093376 0 0.00093368 0 0.0009337799999999999 3.3 0.0009337 3.3 0.0009337999999999999 0 0.0009337200000000001 0 0.00093382 3.3 0.0009337400000000001 3.3 0.00093384 0 0.0009337600000000001 0 0.00093386 3.3 0.00093378 3.3 0.00093388 0 0.0009338 0 0.0009339 3.3 0.00093382 3.3 0.00093392 0 0.00093384 0 0.00093394 3.3 0.00093386 3.3 0.00093396 0 0.00093388 0 0.0009339799999999999 3.3 0.0009339 3.3 0.0009339999999999999 0 0.0009339200000000001 0 0.00093402 3.3 0.0009339400000000001 3.3 0.00093404 0 0.0009339600000000001 0 0.00093406 3.3 0.00093398 3.3 0.00093408 0 0.000934 0 0.0009341 3.3 0.00093402 3.3 0.00093412 0 0.00093404 0 0.00093414 3.3 0.00093406 3.3 0.00093416 0 0.00093408 0 0.00093418 3.3 0.0009341 3.3 0.0009341999999999999 0 0.00093412 0 0.0009342199999999999 3.3 0.0009341400000000001 3.3 0.00093424 0 0.0009341600000000001 0 0.00093426 3.3 0.0009341800000000001 3.3 0.00093428 0 0.0009342 0 0.0009343 3.3 0.00093422 3.3 0.00093432 0 0.00093424 0 0.00093434 3.3 0.00093426 3.3 0.00093436 0 0.00093428 0 0.00093438 3.3 0.0009343 3.3 0.0009343999999999999 0 0.00093432 0 0.0009344199999999999 3.3 0.0009343400000000001 3.3 0.00093444 0 0.0009343600000000001 0 0.00093446 3.3 0.0009343800000000001 3.3 0.00093448 0 0.0009344 0 0.0009345 3.3 0.00093442 3.3 0.00093452 0 0.00093444 0 0.00093454 3.3 0.00093446 3.3 0.00093456 0 0.00093448 0 0.00093458 3.3 0.0009345 3.3 0.0009346 0 0.00093452 0 0.0009346199999999999 3.3 0.00093454 3.3 0.0009346399999999999 0 0.0009345600000000001 0 0.00093466 3.3 0.0009345800000000001 3.3 0.00093468 0 0.0009346000000000001 0 0.0009347 3.3 0.00093462 3.3 0.00093472 0 0.00093464 0 0.00093474 3.3 0.00093466 3.3 0.00093476 0 0.00093468 0 0.00093478 3.3 0.0009347 3.3 0.0009348 0 0.00093472 0 0.0009348199999999999 3.3 0.00093474 3.3 0.0009348399999999999 0 0.0009347600000000001 0 0.00093486 3.3 0.0009347800000000001 3.3 0.00093488 0 0.0009348000000000001 0 0.0009349 3.3 0.00093482 3.3 0.00093492 0 0.00093484 0 0.00093494 3.3 0.00093486 3.3 0.00093496 0 0.00093488 0 0.00093498 3.3 0.0009349 3.3 0.000935 0 0.00093492 0 0.00093502 3.3 0.00093494 3.3 0.0009350399999999999 0 0.00093496 0 0.0009350599999999999 3.3 0.0009349800000000001 3.3 0.00093508 0 0.0009350000000000001 0 0.0009351 3.3 0.0009350200000000001 3.3 0.00093512 0 0.00093504 0 0.00093514 3.3 0.00093506 3.3 0.00093516 0 0.00093508 0 0.00093518 3.3 0.0009351 3.3 0.0009352 0 0.00093512 0 0.00093522 3.3 0.00093514 3.3 0.0009352399999999999 0 0.00093516 0 0.0009352599999999999 3.3 0.0009351800000000001 3.3 0.00093528 0 0.0009352000000000001 0 0.0009353 3.3 0.0009352200000000001 3.3 0.00093532 0 0.00093524 0 0.00093534 3.3 0.00093526 3.3 0.00093536 0 0.00093528 0 0.00093538 3.3 0.0009353 3.3 0.0009354 0 0.00093532 0 0.00093542 3.3 0.00093534 3.3 0.00093544 0 0.00093536 0 0.0009354599999999999 3.3 0.00093538 3.3 0.0009354799999999999 0 0.0009354000000000001 0 0.0009355 3.3 0.0009354200000000001 3.3 0.00093552 0 0.0009354400000000001 0 0.00093554 3.3 0.00093546 3.3 0.00093556 0 0.00093548 0 0.00093558 3.3 0.0009355 3.3 0.0009356 0 0.00093552 0 0.00093562 3.3 0.00093554 3.3 0.00093564 0 0.00093556 0 0.0009356599999999999 3.3 0.00093558 3.3 0.0009356799999999999 0 0.0009356000000000001 0 0.0009357 3.3 0.0009356200000000001 3.3 0.00093572 0 0.0009356400000000001 0 0.00093574 3.3 0.00093566 3.3 0.00093576 0 0.00093568 0 0.00093578 3.3 0.0009357 3.3 0.0009358 0 0.00093572 0 0.00093582 3.3 0.00093574 3.3 0.00093584 0 0.00093576 0 0.00093586 3.3 0.00093578 3.3 0.0009358799999999999 0 0.0009358000000000001 0 0.0009359 3.3 0.0009358200000000001 3.3 0.00093592 0 0.0009358400000000001 0 0.00093594 3.3 0.0009358600000000001 3.3 0.00093596 0 0.00093588 0 0.00093598 3.3 0.0009359 3.3 0.000936 0 0.00093592 0 0.00093602 3.3 0.00093594 3.3 0.00093604 0 0.00093596 0 0.00093606 3.3 0.00093598 3.3 0.0009360799999999999 0 0.000936 0 0.0009360999999999999 3.3 0.0009360200000000001 3.3 0.00093612 0 0.0009360400000000001 0 0.00093614 3.3 0.0009360600000000001 3.3 0.00093616 0 0.00093608 0 0.00093618 3.3 0.0009361 3.3 0.0009362 0 0.00093612 0 0.00093622 3.3 0.00093614 3.3 0.00093624 0 0.00093616 0 0.00093626 3.3 0.00093618 3.3 0.00093628 0 0.0009362 0 0.0009362999999999999 3.3 0.0009362200000000001 3.3 0.00093632 0 0.0009362400000000001 0 0.00093634 3.3 0.0009362600000000001 3.3 0.00093636 0 0.0009362800000000001 0 0.00093638 3.3 0.0009363 3.3 0.0009364 0 0.00093632 0 0.00093642 3.3 0.00093634 3.3 0.00093644 0 0.00093636 0 0.00093646 3.3 0.00093638 3.3 0.00093648 0 0.0009364 0 0.0009364999999999999 3.3 0.00093642 3.3 0.0009365199999999999 0 0.0009364400000000001 0 0.00093654 3.3 0.0009364600000000001 3.3 0.00093656 0 0.0009364800000000001 0 0.00093658 3.3 0.0009365 3.3 0.0009366 0 0.00093652 0 0.00093662 3.3 0.00093654 3.3 0.00093664 0 0.00093656 0 0.00093666 3.3 0.00093658 3.3 0.00093668 0 0.0009366 0 0.0009367 3.3 0.00093662 3.3 0.0009367199999999999 0 0.0009366400000000001 0 0.00093674 3.3 0.0009366600000000001 3.3 0.00093676 0 0.0009366800000000001 0 0.00093678 3.3 0.0009367000000000001 3.3 0.0009368 0 0.00093672 0 0.00093682 3.3 0.00093674 3.3 0.00093684 0 0.00093676 0 0.00093686 3.3 0.00093678 3.3 0.00093688 0 0.0009368 0 0.0009369 3.3 0.00093682 3.3 0.0009369199999999999 0 0.00093684 0 0.0009369399999999999 3.3 0.0009368600000000001 3.3 0.00093696 0 0.0009368800000000001 0 0.00093698 3.3 0.0009369000000000001 3.3 0.000937 0 0.00093692 0 0.00093702 3.3 0.00093694 3.3 0.00093704 0 0.00093696 0 0.00093706 3.3 0.00093698 3.3 0.00093708 0 0.000937 0 0.0009371 3.3 0.00093702 3.3 0.0009371199999999999 0 0.00093704 0 0.0009371399999999999 3.3 0.0009370600000000001 3.3 0.00093716 0 0.0009370800000000001 0 0.00093718 3.3 0.0009371000000000001 3.3 0.0009372 0 0.00093712 0 0.00093722 3.3 0.00093714 3.3 0.00093724 0 0.00093716 0 0.00093726 3.3 0.00093718 3.3 0.00093728 0 0.0009372 0 0.0009373 3.3 0.00093722 3.3 0.00093732 0 0.00093724 0 0.0009373399999999999 3.3 0.00093726 3.3 0.0009373599999999999 0 0.0009372800000000001 0 0.00093738 3.3 0.0009373000000000001 3.3 0.0009374 0 0.0009373200000000001 0 0.00093742 3.3 0.00093734 3.3 0.00093744 0 0.00093736 0 0.00093746 3.3 0.00093738 3.3 0.00093748 0 0.0009374 0 0.0009375 3.3 0.00093742 3.3 0.00093752 0 0.00093744 0 0.0009375399999999999 3.3 0.00093746 3.3 0.0009375599999999999 0 0.0009374800000000001 0 0.00093758 3.3 0.0009375000000000001 3.3 0.0009376 0 0.0009375200000000001 0 0.00093762 3.3 0.00093754 3.3 0.00093764 0 0.00093756 0 0.00093766 3.3 0.00093758 3.3 0.00093768 0 0.0009376 0 0.0009377 3.3 0.00093762 3.3 0.00093772 0 0.00093764 0 0.00093774 3.3 0.00093766 3.3 0.0009377599999999999 0 0.00093768 0 0.0009377799999999999 3.3 0.0009377000000000001 3.3 0.0009378 0 0.0009377200000000001 0 0.00093782 3.3 0.0009377400000000001 3.3 0.00093784 0 0.00093776 0 0.00093786 3.3 0.00093778 3.3 0.00093788 0 0.0009378 0 0.0009379 3.3 0.00093782 3.3 0.00093792 0 0.00093784 0 0.00093794 3.3 0.00093786 3.3 0.0009379599999999999 0 0.00093788 0 0.0009379799999999999 3.3 0.0009379000000000001 3.3 0.000938 0 0.0009379200000000001 0 0.00093802 3.3 0.0009379400000000001 3.3 0.00093804 0 0.00093796 0 0.00093806 3.3 0.00093798 3.3 0.00093808 0 0.000938 0 0.0009381 3.3 0.00093802 3.3 0.00093812 0 0.00093804 0 0.00093814 3.3 0.00093806 3.3 0.00093816 0 0.00093808 0 0.0009381799999999999 3.3 0.0009381 3.3 0.0009381999999999999 0 0.0009381200000000001 0 0.00093822 3.3 0.0009381400000000001 3.3 0.00093824 0 0.0009381600000000001 0 0.00093826 3.3 0.00093818 3.3 0.00093828 0 0.0009382 0 0.0009383 3.3 0.00093822 3.3 0.00093832 0 0.00093824 0 0.00093834 3.3 0.00093826 3.3 0.00093836 0 0.00093828 0 0.0009383799999999999 3.3 0.0009383 3.3 0.0009383999999999999 0 0.0009383200000000001 0 0.00093842 3.3 0.0009383400000000001 3.3 0.00093844 0 0.0009383600000000001 0 0.00093846 3.3 0.00093838 3.3 0.00093848 0 0.0009384 0 0.0009385 3.3 0.00093842 3.3 0.00093852 0 0.00093844 0 0.00093854 3.3 0.00093846 3.3 0.00093856 0 0.00093848 0 0.00093858 3.3 0.0009385 3.3 0.0009385999999999999 0 0.00093852 0 0.0009386199999999999 3.3 0.0009385400000000001 3.3 0.00093864 0 0.0009385600000000001 0 0.00093866 3.3 0.0009385800000000001 3.3 0.00093868 0 0.0009386 0 0.0009387 3.3 0.00093862 3.3 0.00093872 0 0.00093864 0 0.00093874 3.3 0.00093866 3.3 0.00093876 0 0.00093868 0 0.00093878 3.3 0.0009387 3.3 0.0009387999999999999 0 0.00093872 0 0.0009388199999999999 3.3 0.0009387400000000001 3.3 0.00093884 0 0.0009387600000000001 0 0.00093886 3.3 0.0009387800000000001 3.3 0.00093888 0 0.0009388 0 0.0009389 3.3 0.00093882 3.3 0.00093892 0 0.00093884 0 0.00093894 3.3 0.00093886 3.3 0.00093896 0 0.00093888 0 0.00093898 3.3 0.0009389 3.3 0.000939 0 0.00093892 0 0.0009390199999999999 3.3 0.0009389400000000001 3.3 0.00093904 0 0.0009389600000000001 0 0.00093906 3.3 0.0009389800000000001 3.3 0.00093908 0 0.0009390000000000001 0 0.0009391 3.3 0.00093902 3.3 0.00093912 0 0.00093904 0 0.00093914 3.3 0.00093906 3.3 0.00093916 0 0.00093908 0 0.00093918 3.3 0.0009391 3.3 0.0009392 0 0.00093912 0 0.0009392199999999999 3.3 0.00093914 3.3 0.0009392399999999999 0 0.0009391600000000001 0 0.00093926 3.3 0.0009391800000000001 3.3 0.00093928 0 0.0009392000000000001 0 0.0009393 3.3 0.00093922 3.3 0.00093932 0 0.00093924 0 0.00093934 3.3 0.00093926 3.3 0.00093936 0 0.00093928 0 0.00093938 3.3 0.0009393 3.3 0.0009394 0 0.00093932 0 0.00093942 3.3 0.00093934 3.3 0.0009394399999999999 0 0.0009393600000000001 0 0.00093946 3.3 0.0009393800000000001 3.3 0.00093948 0 0.0009394000000000001 0 0.0009395 3.3 0.0009394200000000001 3.3 0.00093952 0 0.00093944 0 0.00093954 3.3 0.00093946 3.3 0.00093956 0 0.00093948 0 0.00093958 3.3 0.0009395 3.3 0.0009396 0 0.00093952 0 0.00093962 3.3 0.00093954 3.3 0.0009396399999999999 0 0.00093956 0 0.0009396599999999999 3.3 0.0009395800000000001 3.3 0.00093968 0 0.0009396000000000001 0 0.0009397 3.3 0.0009396200000000001 3.3 0.00093972 0 0.00093964 0 0.00093974 3.3 0.00093966 3.3 0.00093976 0 0.00093968 0 0.00093978 3.3 0.0009397 3.3 0.0009398 0 0.00093972 0 0.00093982 3.3 0.00093974 3.3 0.00093984 0 0.00093976 0 0.0009398599999999999 3.3 0.0009397800000000001 3.3 0.00093988 0 0.0009398000000000001 0 0.0009399 3.3 0.0009398200000000001 3.3 0.00093992 0 0.0009398400000000001 0 0.00093994 3.3 0.00093986 3.3 0.00093996 0 0.00093988 0 0.00093998 3.3 0.0009399 3.3 0.00094 0 0.00093992 0 0.00094002 3.3 0.00093994 3.3 0.00094004 0 0.00093996 0 0.0009400599999999999 3.3 0.00093998 3.3 0.0009400799999999999 0 0.0009400000000000001 0 0.0009401 3.3 0.0009400200000000001 3.3 0.00094012 0 0.0009400400000000001 0 0.00094014 3.3 0.00094006 3.3 0.00094016 0 0.00094008 0 0.00094018 3.3 0.0009401 3.3 0.0009402 0 0.00094012 0 0.00094022 3.3 0.00094014 3.3 0.00094024 0 0.00094016 0 0.0009402599999999999 3.3 0.00094018 3.3 0.0009402799999999999 0 0.0009402000000000001 0 0.0009403 3.3 0.0009402200000000001 3.3 0.00094032 0 0.0009402400000000001 0 0.00094034 3.3 0.00094026 3.3 0.00094036 0 0.00094028 0 0.00094038 3.3 0.0009403 3.3 0.0009404 0 0.00094032 0 0.00094042 3.3 0.00094034 3.3 0.00094044 0 0.00094036 0 0.00094046 3.3 0.00094038 3.3 0.0009404799999999999 0 0.0009404 0 0.0009404999999999999 3.3 0.0009404200000000001 3.3 0.00094052 0 0.0009404400000000001 0 0.00094054 3.3 0.0009404600000000001 3.3 0.00094056 0 0.00094048 0 0.00094058 3.3 0.0009405 3.3 0.0009406 0 0.00094052 0 0.00094062 3.3 0.00094054 3.3 0.00094064 0 0.00094056 0 0.00094066 3.3 0.00094058 3.3 0.0009406799999999999 0 0.0009406 0 0.0009406999999999999 3.3 0.0009406200000000001 3.3 0.00094072 0 0.0009406400000000001 0 0.00094074 3.3 0.0009406600000000001 3.3 0.00094076 0 0.00094068 0 0.00094078 3.3 0.0009407 3.3 0.0009408 0 0.00094072 0 0.00094082 3.3 0.00094074 3.3 0.00094084 0 0.00094076 0 0.00094086 3.3 0.00094078 3.3 0.00094088 0 0.0009408 0 0.0009408999999999999 3.3 0.00094082 3.3 0.0009409199999999999 0 0.0009408400000000001 0 0.00094094 3.3 0.0009408600000000001 3.3 0.00094096 0 0.0009408800000000001 0 0.00094098 3.3 0.0009409 3.3 0.000941 0 0.00094092 0 0.00094102 3.3 0.00094094 3.3 0.00094104 0 0.00094096 0 0.00094106 3.3 0.00094098 3.3 0.00094108 0 0.000941 0 0.0009410999999999999 3.3 0.00094102 3.3 0.0009411199999999999 0 0.0009410400000000001 0 0.00094114 3.3 0.0009410600000000001 3.3 0.00094116 0 0.0009410800000000001 0 0.00094118 3.3 0.0009411 3.3 0.0009412 0 0.00094112 0 0.00094122 3.3 0.00094114 3.3 0.00094124 0 0.00094116 0 0.00094126 3.3 0.00094118 3.3 0.00094128 0 0.0009412 0 0.0009413 3.3 0.00094122 3.3 0.0009413199999999999 0 0.00094124 0 0.0009413399999999999 3.3 0.0009412600000000001 3.3 0.00094136 0 0.0009412800000000001 0 0.00094138 3.3 0.0009413000000000001 3.3 0.0009414 0 0.00094132 0 0.00094142 3.3 0.00094134 3.3 0.00094144 0 0.00094136 0 0.00094146 3.3 0.00094138 3.3 0.00094148 0 0.0009414 0 0.0009415 3.3 0.00094142 3.3 0.0009415199999999999 0 0.00094144 0 0.0009415399999999999 3.3 0.0009414600000000001 3.3 0.00094156 0 0.0009414800000000001 0 0.00094158 3.3 0.0009415000000000001 3.3 0.0009416 0 0.00094152 0 0.00094162 3.3 0.00094154 3.3 0.00094164 0 0.00094156 0 0.00094166 3.3 0.00094158 3.3 0.00094168 0 0.0009416 0 0.0009417 3.3 0.00094162 3.3 0.00094172 0 0.00094164 0 0.0009417399999999999 3.3 0.00094166 3.3 0.0009417599999999999 0 0.0009416800000000001 0 0.00094178 3.3 0.0009417000000000001 3.3 0.0009418 0 0.0009417200000000001 0 0.00094182 3.3 0.00094174 3.3 0.00094184 0 0.00094176 0 0.00094186 3.3 0.00094178 3.3 0.00094188 0 0.0009418 0 0.0009419 3.3 0.00094182 3.3 0.00094192 0 0.00094184 0 0.0009419399999999999 3.3 0.00094186 3.3 0.0009419599999999999 0 0.0009418800000000001 0 0.00094198 3.3 0.0009419000000000001 3.3 0.000942 0 0.0009419200000000001 0 0.00094202 3.3 0.00094194 3.3 0.00094204 0 0.00094196 0 0.00094206 3.3 0.00094198 3.3 0.00094208 0 0.000942 0 0.0009421 3.3 0.00094202 3.3 0.00094212 0 0.00094204 0 0.00094214 3.3 0.00094206 3.3 0.0009421599999999999 0 0.00094208 0 0.0009421799999999999 3.3 0.0009421000000000001 3.3 0.0009422 0 0.0009421200000000001 0 0.00094222 3.3 0.0009421400000000001 3.3 0.00094224 0 0.00094216 0 0.00094226 3.3 0.00094218 3.3 0.00094228 0 0.0009422 0 0.0009423 3.3 0.00094222 3.3 0.00094232 0 0.00094224 0 0.00094234 3.3 0.00094226 3.3 0.0009423599999999999 0 0.00094228 0 0.0009423799999999999 3.3 0.0009423000000000001 3.3 0.0009424 0 0.0009423200000000001 0 0.00094242 3.3 0.0009423400000000001 3.3 0.00094244 0 0.00094236 0 0.00094246 3.3 0.00094238 3.3 0.00094248 0 0.0009424 0 0.0009425 3.3 0.00094242 3.3 0.00094252 0 0.00094244 0 0.00094254 3.3 0.00094246 3.3 0.00094256 0 0.00094248 0 0.0009425799999999999 3.3 0.0009425000000000001 3.3 0.0009426 0 0.0009425200000000001 0 0.00094262 3.3 0.0009425400000000001 3.3 0.00094264 0 0.0009425600000000001 0 0.00094266 3.3 0.00094258 3.3 0.00094268 0 0.0009426 0 0.0009427 3.3 0.00094262 3.3 0.00094272 0 0.00094264 0 0.00094274 3.3 0.00094266 3.3 0.00094276 0 0.00094268 0 0.0009427799999999999 3.3 0.0009427 3.3 0.0009427999999999999 0 0.0009427200000000001 0 0.00094282 3.3 0.0009427400000000001 3.3 0.00094284 0 0.0009427600000000001 0 0.00094286 3.3 0.00094278 3.3 0.00094288 0 0.0009428 0 0.0009429 3.3 0.00094282 3.3 0.00094292 0 0.00094284 0 0.00094294 3.3 0.00094286 3.3 0.00094296 0 0.00094288 0 0.00094298 3.3 0.0009429 3.3 0.0009429999999999999 0 0.0009429200000000001 0 0.00094302 3.3 0.0009429400000000001 3.3 0.00094304 0 0.0009429600000000001 0 0.00094306 3.3 0.0009429800000000001 3.3 0.00094308 0 0.000943 0 0.0009431 3.3 0.00094302 3.3 0.00094312 0 0.00094304 0 0.00094314 3.3 0.00094306 3.3 0.00094316 0 0.00094308 0 0.00094318 3.3 0.0009431 3.3 0.0009431999999999999 0 0.00094312 0 0.0009432199999999999 3.3 0.0009431400000000001 3.3 0.00094324 0 0.0009431600000000001 0 0.00094326 3.3 0.0009431800000000001 3.3 0.00094328 0 0.0009432 0 0.0009433 3.3 0.00094322 3.3 0.00094332 0 0.00094324 0 0.00094334 3.3 0.00094326 3.3 0.00094336 0 0.00094328 0 0.00094338 3.3 0.0009433 3.3 0.0009434 0 0.00094332 0 0.0009434199999999999 3.3 0.0009433400000000001 3.3 0.00094344 0 0.0009433600000000001 0 0.00094346 3.3 0.0009433800000000001 3.3 0.00094348 0 0.0009434000000000001 0 0.0009435 3.3 0.00094342 3.3 0.00094352 0 0.00094344 0 0.00094354 3.3 0.00094346 3.3 0.00094356 0 0.00094348 0 0.00094358 3.3 0.0009435 3.3 0.0009436 0 0.00094352 0 0.0009436199999999999 3.3 0.00094354 3.3 0.0009436399999999999 0 0.0009435600000000001 0 0.00094366 3.3 0.0009435800000000001 3.3 0.00094368 0 0.0009436000000000001 0 0.0009437 3.3 0.00094362 3.3 0.00094372 0 0.00094364 0 0.00094374 3.3 0.00094366 3.3 0.00094376 0 0.00094368 0 0.00094378 3.3 0.0009437 3.3 0.0009438 0 0.00094372 0 0.0009438199999999999 3.3 0.00094374 3.3 0.0009438399999999999 0 0.0009437600000000001 0 0.00094386 3.3 0.0009437800000000001 3.3 0.00094388 0 0.0009438000000000001 0 0.0009439 3.3 0.00094382 3.3 0.00094392 0 0.00094384 0 0.00094394 3.3 0.00094386 3.3 0.00094396 0 0.00094388 0 0.00094398 3.3 0.0009439 3.3 0.000944 0 0.00094392 0 0.00094402 3.3 0.00094394 3.3 0.0009440399999999999 0 0.00094396 0 0.0009440599999999999 3.3 0.0009439800000000001 3.3 0.00094408 0 0.0009440000000000001 0 0.0009441 3.3 0.0009440200000000001 3.3 0.00094412 0 0.00094404 0 0.00094414 3.3 0.00094406 3.3 0.00094416 0 0.00094408 0 0.00094418 3.3 0.0009441 3.3 0.0009442 0 0.00094412 0 0.00094422 3.3 0.00094414 3.3 0.0009442399999999999 0 0.00094416 0 0.0009442599999999999 3.3 0.0009441800000000001 3.3 0.00094428 0 0.0009442000000000001 0 0.0009443 3.3 0.0009442200000000001 3.3 0.00094432 0 0.00094424 0 0.00094434 3.3 0.00094426 3.3 0.00094436 0 0.00094428 0 0.00094438 3.3 0.0009443 3.3 0.0009444 0 0.00094432 0 0.00094442 3.3 0.00094434 3.3 0.00094444 0 0.00094436 0 0.0009444599999999999 3.3 0.00094438 3.3 0.0009444799999999999 0 0.0009444000000000001 0 0.0009445 3.3 0.0009444200000000001 3.3 0.00094452 0 0.0009444400000000001 0 0.00094454 3.3 0.00094446 3.3 0.00094456 0 0.00094448 0 0.00094458 3.3 0.0009445 3.3 0.0009446 0 0.00094452 0 0.00094462 3.3 0.00094454 3.3 0.00094464 0 0.00094456 0 0.0009446599999999999 3.3 0.00094458 3.3 0.0009446799999999999 0 0.0009446000000000001 0 0.0009447 3.3 0.0009446200000000001 3.3 0.00094472 0 0.0009446400000000001 0 0.00094474 3.3 0.00094466 3.3 0.00094476 0 0.00094468 0 0.00094478 3.3 0.0009447 3.3 0.0009448 0 0.00094472 0 0.00094482 3.3 0.00094474 3.3 0.00094484 0 0.00094476 0 0.00094486 3.3 0.00094478 3.3 0.0009448799999999999 0 0.0009448 0 0.0009448999999999999 3.3 0.0009448200000000001 3.3 0.00094492 0 0.0009448400000000001 0 0.00094494 3.3 0.0009448600000000001 3.3 0.00094496 0 0.00094488 0 0.00094498 3.3 0.0009449 3.3 0.000945 0 0.00094492 0 0.00094502 3.3 0.00094494 3.3 0.00094504 0 0.00094496 0 0.00094506 3.3 0.00094498 3.3 0.0009450799999999999 0 0.000945 0 0.0009450999999999999 3.3 0.0009450200000000001 3.3 0.00094512 0 0.0009450400000000001 0 0.00094514 3.3 0.0009450600000000001 3.3 0.00094516 0 0.00094508 0 0.00094518 3.3 0.0009451 3.3 0.0009452 0 0.00094512 0 0.00094522 3.3 0.00094514 3.3 0.00094524 0 0.00094516 0 0.00094526 3.3 0.00094518 3.3 0.00094528 0 0.0009452 0 0.0009452999999999999 3.3 0.00094522 3.3 0.0009453199999999999 0 0.0009452400000000001 0 0.00094534 3.3 0.0009452600000000001 3.3 0.00094536 0 0.0009452800000000001 0 0.00094538 3.3 0.0009453 3.3 0.0009454 0 0.00094532 0 0.00094542 3.3 0.00094534 3.3 0.00094544 0 0.00094536 0 0.00094546 3.3 0.00094538 3.3 0.00094548 0 0.0009454 0 0.0009454999999999999 3.3 0.00094542 3.3 0.0009455199999999999 0 0.0009454400000000001 0 0.00094554 3.3 0.0009454600000000001 3.3 0.00094556 0 0.0009454800000000001 0 0.00094558 3.3 0.0009455 3.3 0.0009456 0 0.00094552 0 0.00094562 3.3 0.00094554 3.3 0.00094564 0 0.00094556 0 0.00094566 3.3 0.00094558 3.3 0.00094568 0 0.0009456 0 0.0009457 3.3 0.00094562 3.3 0.0009457199999999999 0 0.00094564 0 0.0009457399999999999 3.3 0.0009456600000000001 3.3 0.00094576 0 0.0009456800000000001 0 0.00094578 3.3 0.0009457000000000001 3.3 0.0009458 0 0.00094572 0 0.00094582 3.3 0.00094574 3.3 0.00094584 0 0.00094576 0 0.00094586 3.3 0.00094578 3.3 0.00094588 0 0.0009458 0 0.0009459 3.3 0.00094582 3.3 0.0009459199999999999 0 0.00094584 0 0.0009459399999999999 3.3 0.0009458600000000001 3.3 0.00094596 0 0.0009458800000000001 0 0.00094598 3.3 0.0009459000000000001 3.3 0.000946 0 0.00094592 0 0.00094602 3.3 0.00094594 3.3 0.00094604 0 0.00094596 0 0.00094606 3.3 0.00094598 3.3 0.00094608 0 0.000946 0 0.0009461 3.3 0.00094602 3.3 0.00094612 0 0.00094604 0 0.0009461399999999999 3.3 0.0009460600000000001 3.3 0.00094616 0 0.0009460800000000001 0 0.00094618 3.3 0.0009461000000000001 3.3 0.0009462 0 0.0009461200000000001 0 0.00094622 3.3 0.00094614 3.3 0.00094624 0 0.00094616 0 0.00094626 3.3 0.00094618 3.3 0.00094628 0 0.0009462 0 0.0009463 3.3 0.00094622 3.3 0.00094632 0 0.00094624 0 0.0009463399999999999 3.3 0.00094626 3.3 0.0009463599999999999 0 0.0009462800000000001 0 0.00094638 3.3 0.0009463000000000001 3.3 0.0009464 0 0.0009463200000000001 0 0.00094642 3.3 0.00094634 3.3 0.00094644 0 0.00094636 0 0.00094646 3.3 0.00094638 3.3 0.00094648 0 0.0009464 0 0.0009465 3.3 0.00094642 3.3 0.00094652 0 0.00094644 0 0.00094654 3.3 0.00094646 3.3 0.0009465599999999999 0 0.0009464800000000001 0 0.00094658 3.3 0.0009465000000000001 3.3 0.0009466 0 0.0009465200000000001 0 0.00094662 3.3 0.0009465400000000001 3.3 0.00094664 0 0.00094656 0 0.00094666 3.3 0.00094658 3.3 0.00094668 0 0.0009466 0 0.0009467 3.3 0.00094662 3.3 0.00094672 0 0.00094664 0 0.00094674 3.3 0.00094666 3.3 0.0009467599999999999 0 0.00094668 0 0.0009467799999999999 3.3 0.0009467000000000001 3.3 0.0009468 0 0.0009467200000000001 0 0.00094682 3.3 0.0009467400000000001 3.3 0.00094684 0 0.00094676 0 0.00094686 3.3 0.00094678 3.3 0.00094688 0 0.0009468 0 0.0009469 3.3 0.00094682 3.3 0.00094692 0 0.00094684 0 0.00094694 3.3 0.00094686 3.3 0.00094696 0 0.00094688 0 0.0009469799999999999 3.3 0.0009469000000000001 3.3 0.000947 0 0.0009469200000000001 0 0.00094702 3.3 0.0009469400000000001 3.3 0.00094704 0 0.0009469600000000001 0 0.00094706 3.3 0.00094698 3.3 0.00094708 0 0.000947 0 0.0009471 3.3 0.00094702 3.3 0.00094712 0 0.00094704 0 0.00094714 3.3 0.00094706 3.3 0.00094716 0 0.00094708 0 0.0009471799999999999 3.3 0.0009471 3.3 0.0009471999999999999 0 0.0009471200000000001 0 0.00094722 3.3 0.0009471400000000001 3.3 0.00094724 0 0.0009471600000000001 0 0.00094726 3.3 0.00094718 3.3 0.00094728 0 0.0009472 0 0.0009473 3.3 0.00094722 3.3 0.00094732 0 0.00094724 0 0.00094734 3.3 0.00094726 3.3 0.00094736 0 0.00094728 0 0.0009473799999999999 3.3 0.0009473 3.3 0.0009473999999999999 0 0.0009473200000000001 0 0.00094742 3.3 0.0009473400000000001 3.3 0.00094744 0 0.0009473600000000001 0 0.00094746 3.3 0.00094738 3.3 0.00094748 0 0.0009474 0 0.0009475 3.3 0.00094742 3.3 0.00094752 0 0.00094744 0 0.00094754 3.3 0.00094746 3.3 0.00094756 0 0.00094748 0 0.00094758 3.3 0.0009475 3.3 0.0009475999999999999 0 0.00094752 0 0.0009476199999999999 3.3 0.0009475400000000001 3.3 0.00094764 0 0.0009475600000000001 0 0.00094766 3.3 0.0009475800000000001 3.3 0.00094768 0 0.0009476 0 0.0009477 3.3 0.00094762 3.3 0.00094772 0 0.00094764 0 0.00094774 3.3 0.00094766 3.3 0.00094776 0 0.00094768 0 0.00094778 3.3 0.0009477 3.3 0.0009477999999999999 0 0.00094772 0 0.0009478199999999999 3.3 0.0009477400000000001 3.3 0.00094784 0 0.0009477600000000001 0 0.00094786 3.3 0.0009477800000000001 3.3 0.00094788 0 0.0009478 0 0.0009479 3.3 0.00094782 3.3 0.00094792 0 0.00094784 0 0.00094794 3.3 0.00094786 3.3 0.00094796 0 0.00094788 0 0.00094798 3.3 0.0009479 3.3 0.000948 0 0.00094792 0 0.0009480199999999999 3.3 0.00094794 3.3 0.0009480399999999999 0 0.0009479600000000001 0 0.00094806 3.3 0.0009479800000000001 3.3 0.00094808 0 0.0009480000000000001 0 0.0009481 3.3 0.00094802 3.3 0.00094812 0 0.00094804 0 0.00094814 3.3 0.00094806 3.3 0.00094816 0 0.00094808 0 0.00094818 3.3 0.0009481 3.3 0.0009482 0 0.00094812 0 0.0009482199999999999 3.3 0.00094814 3.3 0.0009482399999999999 0 0.0009481600000000001 0 0.00094826 3.3 0.0009481800000000001 3.3 0.00094828 0 0.0009482000000000001 0 0.0009483 3.3 0.00094822 3.3 0.00094832 0 0.00094824 0 0.00094834 3.3 0.00094826 3.3 0.00094836 0 0.00094828 0 0.00094838 3.3 0.0009483 3.3 0.0009484 0 0.00094832 0 0.00094842 3.3 0.00094834 3.3 0.0009484399999999999 0 0.00094836 0 0.0009484599999999999 3.3 0.0009483800000000001 3.3 0.00094848 0 0.0009484000000000001 0 0.0009485 3.3 0.0009484200000000001 3.3 0.00094852 0 0.00094844 0 0.00094854 3.3 0.00094846 3.3 0.00094856 0 0.00094848 0 0.00094858 3.3 0.0009485 3.3 0.0009486 0 0.00094852 0 0.00094862 3.3 0.00094854 3.3 0.0009486399999999999 0 0.00094856 0 0.0009486599999999999 3.3 0.0009485800000000001 3.3 0.00094868 0 0.0009486000000000001 0 0.0009487 3.3 0.0009486200000000001 3.3 0.00094872 0 0.00094864 0 0.00094874 3.3 0.00094866 3.3 0.00094876 0 0.00094868 0 0.00094878 3.3 0.0009487 3.3 0.0009488 0 0.00094872 0 0.00094882 3.3 0.00094874 3.3 0.00094884 0 0.00094876 0 0.0009488599999999999 3.3 0.00094878 3.3 0.0009488799999999999 0 0.0009488000000000001 0 0.0009489 3.3 0.0009488200000000001 3.3 0.00094892 0 0.0009488400000000001 0 0.00094894 3.3 0.00094886 3.3 0.00094896 0 0.00094888 0 0.00094898 3.3 0.0009489 3.3 0.000949 0 0.00094892 0 0.00094902 3.3 0.00094894 3.3 0.00094904 0 0.00094896 0 0.0009490599999999999 3.3 0.00094898 3.3 0.0009490799999999999 0 0.0009490000000000001 0 0.0009491 3.3 0.0009490200000000001 3.3 0.00094912 0 0.0009490400000000001 0 0.00094914 3.3 0.00094906 3.3 0.00094916 0 0.00094908 0 0.00094918 3.3 0.0009491 3.3 0.0009492 0 0.00094912 0 0.00094922 3.3 0.00094914 3.3 0.00094924 0 0.00094916 0 0.00094926 3.3 0.00094918 3.3 0.0009492799999999999 0 0.0009492 0 0.0009492999999999999 3.3 0.0009492200000000001 3.3 0.00094932 0 0.0009492400000000001 0 0.00094934 3.3 0.0009492600000000001 3.3 0.00094936 0 0.00094928 0 0.00094938 3.3 0.0009493 3.3 0.0009494 0 0.00094932 0 0.00094942 3.3 0.00094934 3.3 0.00094944 0 0.00094936 0 0.00094946 3.3 0.00094938 3.3 0.0009494799999999999 0 0.0009494 0 0.0009494999999999999 3.3 0.0009494200000000001 3.3 0.00094952 0 0.0009494400000000001 0 0.00094954 3.3 0.0009494600000000001 3.3 0.00094956 0 0.00094948 0 0.00094958 3.3 0.0009495 3.3 0.0009496 0 0.00094952 0 0.00094962 3.3 0.00094954 3.3 0.00094964 0 0.00094956 0 0.00094966 3.3 0.00094958 3.3 0.00094968 0 0.0009496 0 0.0009496999999999999 3.3 0.0009496200000000001 3.3 0.00094972 0 0.0009496400000000001 0 0.00094974 3.3 0.0009496600000000001 3.3 0.00094976 0 0.0009496800000000001 0 0.00094978 3.3 0.0009497 3.3 0.0009498 0 0.00094972 0 0.00094982 3.3 0.00094974 3.3 0.00094984 0 0.00094976 0 0.00094986 3.3 0.00094978 3.3 0.00094988 0 0.0009498 0 0.0009498999999999999 3.3 0.00094982 3.3 0.0009499199999999999 0 0.0009498400000000001 0 0.00094994 3.3 0.0009498600000000001 3.3 0.00094996 0 0.0009498800000000001 0 0.00094998 3.3 0.0009499 3.3 0.00095 0 0.00094992 0 0.00095002 3.3 0.00094994 3.3 0.00095004 0 0.00094996 0 0.00095006 3.3 0.00094998 3.3 0.00095008 0 0.00095 0 0.0009501 3.3 0.00095002 3.3 0.0009501199999999999 0 0.0009500400000000001 0 0.00095014 3.3 0.0009500600000000001 3.3 0.00095016 0 0.0009500800000000001 0 0.00095018 3.3 0.0009501000000000001 3.3 0.0009502 0 0.00095012 0 0.00095022 3.3 0.00095014 3.3 0.00095024 0 0.00095016 0 0.00095026 3.3 0.00095018 3.3 0.00095028 0 0.0009502 0 0.0009503 3.3 0.00095022 3.3 0.0009503199999999999 0 0.00095024 0 0.0009503399999999999 3.3 0.0009502600000000001 3.3 0.00095036 0 0.0009502800000000001 0 0.00095038 3.3 0.0009503000000000001 3.3 0.0009504 0 0.00095032 0 0.00095042 3.3 0.00095034 3.3 0.00095044 0 0.00095036 0 0.00095046 3.3 0.00095038 3.3 0.00095048 0 0.0009504 0 0.0009505 3.3 0.00095042 3.3 0.0009505199999999999 0 0.00095044 0 0.0009505399999999999 3.3 0.0009504600000000001 3.3 0.00095056 0 0.0009504800000000001 0 0.00095058 3.3 0.0009505000000000001 3.3 0.0009506 0 0.00095052 0 0.00095062 3.3 0.00095054 3.3 0.00095064 0 0.00095056 0 0.00095066 3.3 0.00095058 3.3 0.00095068 0 0.0009506 0 0.0009507 3.3 0.00095062 3.3 0.00095072 0 0.00095064 0 0.0009507399999999999 3.3 0.00095066 3.3 0.0009507599999999999 0 0.0009506800000000001 0 0.00095078 3.3 0.0009507000000000001 3.3 0.0009508 0 0.0009507200000000001 0 0.00095082 3.3 0.00095074 3.3 0.00095084 0 0.00095076 0 0.00095086 3.3 0.00095078 3.3 0.00095088 0 0.0009508 0 0.0009509 3.3 0.00095082 3.3 0.00095092 0 0.00095084 0 0.0009509399999999999 3.3 0.00095086 3.3 0.0009509599999999999 0 0.0009508800000000001 0 0.00095098 3.3 0.0009509000000000001 3.3 0.000951 0 0.0009509200000000001 0 0.00095102 3.3 0.00095094 3.3 0.00095104 0 0.00095096 0 0.00095106 3.3 0.00095098 3.3 0.00095108 0 0.000951 0 0.0009511 3.3 0.00095102 3.3 0.00095112 0 0.00095104 0 0.00095114 3.3 0.00095106 3.3 0.0009511599999999999 0 0.00095108 0 0.0009511799999999999 3.3 0.0009511000000000001 3.3 0.0009512 0 0.0009511200000000001 0 0.00095122 3.3 0.0009511400000000001 3.3 0.00095124 0 0.00095116 0 0.00095126 3.3 0.00095118 3.3 0.00095128 0 0.0009512 0 0.0009513 3.3 0.00095122 3.3 0.00095132 0 0.00095124 0 0.00095134 3.3 0.00095126 3.3 0.0009513599999999999 0 0.00095128 0 0.0009513799999999999 3.3 0.0009513000000000001 3.3 0.0009514 0 0.0009513200000000001 0 0.00095142 3.3 0.0009513400000000001 3.3 0.00095144 0 0.00095136 0 0.00095146 3.3 0.00095138 3.3 0.00095148 0 0.0009514 0 0.0009515 3.3 0.00095142 3.3 0.00095152 0 0.00095144 0 0.00095154 3.3 0.00095146 3.3 0.00095156 0 0.00095148 0 0.0009515799999999999 3.3 0.0009515 3.3 0.0009515999999999999 0 0.0009515200000000001 0 0.00095162 3.3 0.0009515400000000001 3.3 0.00095164 0 0.0009515600000000001 0 0.00095166 3.3 0.00095158 3.3 0.00095168 0 0.0009516 0 0.0009517 3.3 0.00095162 3.3 0.00095172 0 0.00095164 0 0.00095174 3.3 0.00095166 3.3 0.00095176 0 0.00095168 0 0.0009517799999999999 3.3 0.0009517 3.3 0.0009517999999999999 0 0.0009517200000000001 0 0.00095182 3.3 0.0009517400000000001 3.3 0.00095184 0 0.0009517600000000001 0 0.00095186 3.3 0.00095178 3.3 0.00095188 0 0.0009518 0 0.0009519 3.3 0.00095182 3.3 0.00095192 0 0.00095184 0 0.00095194 3.3 0.00095186 3.3 0.00095196 0 0.00095188 0 0.00095198 3.3 0.0009519 3.3 0.0009519999999999999 0 0.00095192 0 0.0009520199999999999 3.3 0.0009519400000000001 3.3 0.00095204 0 0.0009519600000000001 0 0.00095206 3.3 0.0009519800000000001 3.3 0.00095208 0 0.000952 0 0.0009521 3.3 0.00095202 3.3 0.00095212 0 0.00095204 0 0.00095214 3.3 0.00095206 3.3 0.00095216 0 0.00095208 0 0.00095218 3.3 0.0009521 3.3 0.0009521999999999999 0 0.00095212 0 0.0009522199999999999 3.3 0.0009521400000000001 3.3 0.00095224 0 0.0009521600000000001 0 0.00095226 3.3 0.0009521800000000001 3.3 0.00095228 0 0.0009522 0 0.0009523 3.3 0.00095222 3.3 0.00095232 0 0.00095224 0 0.00095234 3.3 0.00095226 3.3 0.00095236 0 0.00095228 0 0.00095238 3.3 0.0009523 3.3 0.0009524 0 0.00095232 0 0.0009524199999999999 3.3 0.00095234 3.3 0.0009524399999999999 0 0.0009523600000000001 0 0.00095246 3.3 0.0009523800000000001 3.3 0.00095248 0 0.0009524000000000001 0 0.0009525 3.3 0.00095242 3.3 0.00095252 0 0.00095244 0 0.00095254 3.3 0.00095246 3.3 0.00095256 0 0.00095248 0 0.00095258 3.3 0.0009525 3.3 0.0009526 0 0.00095252 0 0.0009526199999999999 3.3 0.00095254 3.3 0.0009526399999999999 0 0.0009525600000000001 0 0.00095266 3.3 0.0009525800000000001 3.3 0.00095268 0 0.0009526000000000001 0 0.0009527 3.3 0.00095262 3.3 0.00095272 0 0.00095264 0 0.00095274 3.3 0.00095266 3.3 0.00095276 0 0.00095268 0 0.00095278 3.3 0.0009527 3.3 0.0009528 0 0.00095272 0 0.00095282 3.3 0.00095274 3.3 0.0009528399999999999 0 0.00095276 0 0.0009528599999999999 3.3 0.0009527800000000001 3.3 0.00095288 0 0.0009528000000000001 0 0.0009529 3.3 0.0009528200000000001 3.3 0.00095292 0 0.00095284 0 0.00095294 3.3 0.00095286 3.3 0.00095296 0 0.00095288 0 0.00095298 3.3 0.0009529 3.3 0.000953 0 0.00095292 0 0.00095302 3.3 0.00095294 3.3 0.0009530399999999999 0 0.00095296 0 0.0009530599999999999 3.3 0.0009529800000000001 3.3 0.00095308 0 0.0009530000000000001 0 0.0009531 3.3 0.0009530200000000001 3.3 0.00095312 0 0.00095304 0 0.00095314 3.3 0.00095306 3.3 0.00095316 0 0.00095308 0 0.00095318 3.3 0.0009531 3.3 0.0009532 0 0.00095312 0 0.00095322 3.3 0.00095314 3.3 0.00095324 0 0.00095316 0 0.0009532599999999999 3.3 0.0009531800000000001 3.3 0.00095328 0 0.0009532000000000001 0 0.0009533 3.3 0.0009532200000000001 3.3 0.00095332 0 0.0009532400000000001 0 0.00095334 3.3 0.00095326 3.3 0.00095336 0 0.00095328 0 0.00095338 3.3 0.0009533 3.3 0.0009534 0 0.00095332 0 0.00095342 3.3 0.00095334 3.3 0.00095344 0 0.00095336 0 0.0009534599999999999 3.3 0.00095338 3.3 0.0009534799999999999 0 0.0009534000000000001 0 0.0009535 3.3 0.0009534200000000001 3.3 0.00095352 0 0.0009534400000000001 0 0.00095354 3.3 0.00095346 3.3 0.00095356 0 0.00095348 0 0.00095358 3.3 0.0009535 3.3 0.0009536 0 0.00095352 0 0.00095362 3.3 0.00095354 3.3 0.00095364 0 0.00095356 0 0.00095366 3.3 0.00095358 3.3 0.0009536799999999999 0 0.0009536000000000001 0 0.0009537 3.3 0.0009536200000000001 3.3 0.00095372 0 0.0009536400000000001 0 0.00095374 3.3 0.0009536600000000001 3.3 0.00095376 0 0.00095368 0 0.00095378 3.3 0.0009537 3.3 0.0009538 0 0.00095372 0 0.00095382 3.3 0.00095374 3.3 0.00095384 0 0.00095376 0 0.00095386 3.3 0.00095378 3.3 0.0009538799999999999 0 0.0009538 0 0.0009538999999999999 3.3 0.0009538200000000001 3.3 0.00095392 0 0.0009538400000000001 0 0.00095394 3.3 0.0009538600000000001 3.3 0.00095396 0 0.00095388 0 0.00095398 3.3 0.0009539 3.3 0.000954 0 0.00095392 0 0.00095402 3.3 0.00095394 3.3 0.00095404 0 0.00095396 0 0.00095406 3.3 0.00095398 3.3 0.0009540799999999999 0 0.000954 0 0.0009540999999999999 3.3 0.0009540200000000001 3.3 0.00095412 0 0.0009540400000000001 0 0.00095414 3.3 0.0009540600000000001 3.3 0.00095416 0 0.00095408 0 0.00095418 3.3 0.0009541 3.3 0.0009542 0 0.00095412 0 0.00095422 3.3 0.00095414 3.3 0.00095424 0 0.00095416 0 0.00095426 3.3 0.00095418 3.3 0.00095428 0 0.0009542 0 0.0009542999999999999 3.3 0.00095422 3.3 0.0009543199999999999 0 0.0009542400000000001 0 0.00095434 3.3 0.0009542600000000001 3.3 0.00095436 0 0.0009542800000000001 0 0.00095438 3.3 0.0009543 3.3 0.0009544 0 0.00095432 0 0.00095442 3.3 0.00095434 3.3 0.00095444 0 0.00095436 0 0.00095446 3.3 0.00095438 3.3 0.00095448 0 0.0009544 0 0.0009544999999999999 3.3 0.00095442 3.3 0.0009545199999999999 0 0.0009544400000000001 0 0.00095454 3.3 0.0009544600000000001 3.3 0.00095456 0 0.0009544800000000001 0 0.00095458 3.3 0.0009545 3.3 0.0009546 0 0.00095452 0 0.00095462 3.3 0.00095454 3.3 0.00095464 0 0.00095456 0 0.00095466 3.3 0.00095458 3.3 0.00095468 0 0.0009546 0 0.0009547 3.3 0.00095462 3.3 0.0009547199999999999 0 0.00095464 0 0.0009547399999999999 3.3 0.0009546600000000001 3.3 0.00095476 0 0.0009546800000000001 0 0.00095478 3.3 0.0009547000000000001 3.3 0.0009548 0 0.00095472 0 0.00095482 3.3 0.00095474 3.3 0.00095484 0 0.00095476 0 0.00095486 3.3 0.00095478 3.3 0.00095488 0 0.0009548 0 0.0009549 3.3 0.00095482 3.3 0.0009549199999999999 0 0.00095484 0 0.0009549399999999999 3.3 0.0009548600000000001 3.3 0.00095496 0 0.0009548800000000001 0 0.00095498 3.3 0.0009549000000000001 3.3 0.000955 0 0.00095492 0 0.00095502 3.3 0.00095494 3.3 0.00095504 0 0.00095496 0 0.00095506 3.3 0.00095498 3.3 0.00095508 0 0.000955 0 0.0009551 3.3 0.00095502 3.3 0.00095512 0 0.00095504 0 0.0009551399999999999 3.3 0.00095506 3.3 0.0009551599999999999 0 0.0009550800000000001 0 0.00095518 3.3 0.0009551000000000001 3.3 0.0009552 0 0.0009551200000000001 0 0.00095522 3.3 0.00095514 3.3 0.00095524 0 0.00095516 0 0.00095526 3.3 0.00095518 3.3 0.00095528 0 0.0009552 0 0.0009553 3.3 0.00095522 3.3 0.00095532 0 0.00095524 0 0.0009553399999999999 3.3 0.00095526 3.3 0.0009553599999999999 0 0.0009552800000000001 0 0.00095538 3.3 0.0009553000000000001 3.3 0.0009554 0 0.0009553200000000001 0 0.00095542 3.3 0.00095534 3.3 0.00095544 0 0.00095536 0 0.00095546 3.3 0.00095538 3.3 0.00095548 0 0.0009554 0 0.0009555 3.3 0.00095542 3.3 0.00095552 0 0.00095544 0 0.00095554 3.3 0.00095546 3.3 0.0009555599999999999 0 0.00095548 0 0.0009555799999999999 3.3 0.0009555000000000001 3.3 0.0009556 0 0.0009555200000000001 0 0.00095562 3.3 0.0009555400000000001 3.3 0.00095564 0 0.00095556 0 0.00095566 3.3 0.00095558 3.3 0.00095568 0 0.0009556 0 0.0009557 3.3 0.00095562 3.3 0.00095572 0 0.00095564 0 0.00095574 3.3 0.00095566 3.3 0.0009557599999999999 0 0.00095568 0 0.0009557799999999999 3.3 0.0009557000000000001 3.3 0.0009558 0 0.0009557200000000001 0 0.00095582 3.3 0.0009557400000000001 3.3 0.00095584 0 0.00095576 0 0.00095586 3.3 0.00095578 3.3 0.00095588 0 0.0009558 0 0.0009559 3.3 0.00095582 3.3 0.00095592 0 0.00095584 0 0.00095594 3.3 0.00095586 3.3 0.00095596 0 0.00095588 0 0.0009559799999999999 3.3 0.0009559 3.3 0.0009559999999999999 0 0.0009559200000000001 0 0.00095602 3.3 0.0009559400000000001 3.3 0.00095604 0 0.0009559600000000001 0 0.00095606 3.3 0.00095598 3.3 0.00095608 0 0.000956 0 0.0009561 3.3 0.00095602 3.3 0.00095612 0 0.00095604 0 0.00095614 3.3 0.00095606 3.3 0.00095616 0 0.00095608 0 0.0009561799999999999 3.3 0.0009561 3.3 0.0009561999999999999 0 0.0009561200000000001 0 0.00095622 3.3 0.0009561400000000001 3.3 0.00095624 0 0.0009561600000000001 0 0.00095626 3.3 0.00095618 3.3 0.00095628 0 0.0009562 0 0.0009563 3.3 0.00095622 3.3 0.00095632 0 0.00095624 0 0.00095634 3.3 0.00095626 3.3 0.00095636 0 0.00095628 0 0.00095638 3.3 0.0009563 3.3 0.0009563999999999999 0 0.0009563200000000001 0 0.00095642 3.3 0.0009563400000000001 3.3 0.00095644 0 0.0009563600000000001 0 0.00095646 3.3 0.0009563800000000001 3.3 0.00095648 0 0.0009564 0 0.0009565 3.3 0.00095642 3.3 0.00095652 0 0.00095644 0 0.00095654 3.3 0.00095646 3.3 0.00095656 0 0.00095648 0 0.00095658 3.3 0.0009565 3.3 0.0009565999999999999 0 0.00095652 0 0.0009566199999999999 3.3 0.0009565400000000001 3.3 0.00095664 0 0.0009565600000000001 0 0.00095666 3.3 0.0009565800000000001 3.3 0.00095668 0 0.0009566 0 0.0009567 3.3 0.00095662 3.3 0.00095672 0 0.00095664 0 0.00095674 3.3 0.00095666 3.3 0.00095676 0 0.00095668 0 0.00095678 3.3 0.0009567 3.3 0.0009568 0 0.00095672 0 0.0009568199999999999 3.3 0.0009567400000000001 3.3 0.00095684 0 0.0009567600000000001 0 0.00095686 3.3 0.0009567800000000001 3.3 0.00095688 0 0.0009568000000000001 0 0.0009569 3.3 0.00095682 3.3 0.00095692 0 0.00095684 0 0.00095694 3.3 0.00095686 3.3 0.00095696 0 0.00095688 0 0.00095698 3.3 0.0009569 3.3 0.000957 0 0.00095692 0 0.0009570199999999999 3.3 0.00095694 3.3 0.0009570399999999999 0 0.0009569600000000001 0 0.00095706 3.3 0.0009569800000000001 3.3 0.00095708 0 0.0009570000000000001 0 0.0009571 3.3 0.00095702 3.3 0.00095712 0 0.00095704 0 0.00095714 3.3 0.00095706 3.3 0.00095716 0 0.00095708 0 0.00095718 3.3 0.0009571 3.3 0.0009572 0 0.00095712 0 0.00095722 3.3 0.00095714 3.3 0.0009572399999999999 0 0.0009571600000000001 0 0.00095726 3.3 0.0009571800000000001 3.3 0.00095728 0 0.0009572000000000001 0 0.0009573 3.3 0.0009572200000000001 3.3 0.00095732 0 0.00095724 0 0.00095734 3.3 0.00095726 3.3 0.00095736 0 0.00095728 0 0.00095738 3.3 0.0009573 3.3 0.0009574 0 0.00095732 0 0.00095742 3.3 0.00095734 3.3 0.0009574399999999999 0 0.00095736 0 0.0009574599999999999 3.3 0.0009573800000000001 3.3 0.00095748 0 0.0009574000000000001 0 0.0009575 3.3 0.0009574200000000001 3.3 0.00095752 0 0.00095744 0 0.00095754 3.3 0.00095746 3.3 0.00095756 0 0.00095748 0 0.00095758 3.3 0.0009575 3.3 0.0009576 0 0.00095752 0 0.00095762 3.3 0.00095754 3.3 0.0009576399999999999 0 0.00095756 0 0.0009576599999999999 3.3 0.0009575800000000001 3.3 0.00095768 0 0.0009576000000000001 0 0.0009577 3.3 0.0009576200000000001 3.3 0.00095772 0 0.00095764 0 0.00095774 3.3 0.00095766 3.3 0.00095776 0 0.00095768 0 0.00095778 3.3 0.0009577 3.3 0.0009578 0 0.00095772 0 0.00095782 3.3 0.00095774 3.3 0.00095784 0 0.00095776 0 0.0009578599999999999 3.3 0.00095778 3.3 0.0009578799999999999 0 0.0009578000000000001 0 0.0009579 3.3 0.0009578200000000001 3.3 0.00095792 0 0.0009578400000000001 0 0.00095794 3.3 0.00095786 3.3 0.00095796 0 0.00095788 0 0.00095798 3.3 0.0009579 3.3 0.000958 0 0.00095792 0 0.00095802 3.3 0.00095794 3.3 0.00095804 0 0.00095796 0 0.0009580599999999999 3.3 0.00095798 3.3 0.0009580799999999999 0 0.0009580000000000001 0 0.0009581 3.3 0.0009580200000000001 3.3 0.00095812 0 0.0009580400000000001 0 0.00095814 3.3 0.00095806 3.3 0.00095816 0 0.00095808 0 0.00095818 3.3 0.0009581 3.3 0.0009582 0 0.00095812 0 0.00095822 3.3 0.00095814 3.3 0.00095824 0 0.00095816 0 0.00095826 3.3 0.00095818 3.3 0.0009582799999999999 0 0.0009582 0 0.0009582999999999999 3.3 0.0009582200000000001 3.3 0.00095832 0 0.0009582400000000001 0 0.00095834 3.3 0.0009582600000000001 3.3 0.00095836 0 0.00095828 0 0.00095838 3.3 0.0009583 3.3 0.0009584 0 0.00095832 0 0.00095842 3.3 0.00095834 3.3 0.00095844 0 0.00095836 0 0.00095846 3.3 0.00095838 3.3 0.0009584799999999999 0 0.0009584 0 0.0009584999999999999 3.3 0.0009584200000000001 3.3 0.00095852 0 0.0009584400000000001 0 0.00095854 3.3 0.0009584600000000001 3.3 0.00095856 0 0.00095848 0 0.00095858 3.3 0.0009585 3.3 0.0009586 0 0.00095852 0 0.00095862 3.3 0.00095854 3.3 0.00095864 0 0.00095856 0 0.00095866 3.3 0.00095858 3.3 0.00095868 0 0.0009586 0 0.0009586999999999999 3.3 0.00095862 3.3 0.0009587199999999999 0 0.0009586400000000001 0 0.00095874 3.3 0.0009586600000000001 3.3 0.00095876 0 0.0009586800000000001 0 0.00095878 3.3 0.0009587 3.3 0.0009588 0 0.00095872 0 0.00095882 3.3 0.00095874 3.3 0.00095884 0 0.00095876 0 0.00095886 3.3 0.00095878 3.3 0.00095888 0 0.0009588 0 0.0009588999999999999 3.3 0.00095882 3.3 0.0009589199999999999 0 0.0009588400000000001 0 0.00095894 3.3 0.0009588600000000001 3.3 0.00095896 0 0.0009588800000000001 0 0.00095898 3.3 0.0009589 3.3 0.000959 0 0.00095892 0 0.00095902 3.3 0.00095894 3.3 0.00095904 0 0.00095896 0 0.00095906 3.3 0.00095898 3.3 0.00095908 0 0.000959 0 0.0009591 3.3 0.00095902 3.3 0.0009591199999999999 0 0.00095904 0 0.0009591399999999999 3.3 0.0009590600000000001 3.3 0.00095916 0 0.0009590800000000001 0 0.00095918 3.3 0.0009591000000000001 3.3 0.0009592 0 0.00095912 0 0.00095922 3.3 0.00095914 3.3 0.00095924 0 0.00095916 0 0.00095926 3.3 0.00095918 3.3 0.00095928 0 0.0009592 0 0.0009593 3.3 0.00095922 3.3 0.0009593199999999999 0 0.00095924 0 0.0009593399999999999 3.3 0.0009592600000000001 3.3 0.00095936 0 0.0009592800000000001 0 0.00095938 3.3 0.0009593000000000001 3.3 0.0009594 0 0.00095932 0 0.00095942 3.3 0.00095934 3.3 0.00095944 0 0.00095936 0 0.00095946 3.3 0.00095938 3.3 0.00095948 0 0.0009594 0 0.0009595 3.3 0.00095942 3.3 0.00095952 0 0.00095944 0 0.0009595399999999999 3.3 0.00095946 3.3 0.0009595599999999999 0 0.0009594800000000001 0 0.00095958 3.3 0.0009595000000000001 3.3 0.0009596 0 0.0009595200000000001 0 0.00095962 3.3 0.00095954 3.3 0.00095964 0 0.00095956 0 0.00095966 3.3 0.00095958 3.3 0.00095968 0 0.0009596 0 0.0009597 3.3 0.00095962 3.3 0.00095972 0 0.00095964 0 0.0009597399999999999 3.3 0.00095966 3.3 0.0009597599999999999 0 0.0009596800000000001 0 0.00095978 3.3 0.0009597000000000001 3.3 0.0009598 0 0.0009597200000000001 0 0.00095982 3.3 0.00095974 3.3 0.00095984 0 0.00095976 0 0.00095986 3.3 0.00095978 3.3 0.00095988 0 0.0009598 0 0.0009599 3.3 0.00095982 3.3 0.00095992 0 0.00095984 0 0.00095994 3.3 0.00095986 3.3 0.0009599599999999999 0 0.0009598800000000001 0 0.00095998 3.3 0.0009599000000000001 3.3 0.00096 0 0.0009599200000000001 0 0.00096002 3.3 0.0009599400000000001 3.3 0.00096004 0 0.00095996 0 0.00096006 3.3 0.00095998 3.3 0.00096008 0 0.00096 0 0.0009601 3.3 0.00096002 3.3 0.00096012 0 0.00096004 0 0.00096014 3.3 0.00096006 3.3 0.0009601599999999999 0 0.00096008 0 0.0009601799999999999 3.3 0.0009601000000000001 3.3 0.0009602 0 0.0009601200000000001 0 0.00096022 3.3 0.0009601400000000001 3.3 0.00096024 0 0.00096016 0 0.00096026 3.3 0.00096018 3.3 0.00096028 0 0.0009602 0 0.0009603 3.3 0.00096022 3.3 0.00096032 0 0.00096024 0 0.00096034 3.3 0.00096026 3.3 0.00096036 0 0.00096028 0 0.0009603799999999999 3.3 0.0009603000000000001 3.3 0.0009604 0 0.0009603200000000001 0 0.00096042 3.3 0.0009603400000000001 3.3 0.00096044 0 0.0009603600000000001 0 0.00096046 3.3 0.00096038 3.3 0.00096048 0 0.0009604 0 0.0009605 3.3 0.00096042 3.3 0.00096052 0 0.00096044 0 0.00096054 3.3 0.00096046 3.3 0.00096056 0 0.00096048 0 0.0009605799999999999 3.3 0.0009605 3.3 0.0009605999999999999 0 0.0009605200000000001 0 0.00096062 3.3 0.0009605400000000001 3.3 0.00096064 0 0.0009605600000000001 0 0.00096066 3.3 0.00096058 3.3 0.00096068 0 0.0009606 0 0.0009607 3.3 0.00096062 3.3 0.00096072 0 0.00096064 0 0.00096074 3.3 0.00096066 3.3 0.00096076 0 0.00096068 0 0.0009607799999999999 3.3 0.0009607 3.3 0.0009607999999999999 0 0.0009607200000000001 0 0.00096082 3.3 0.0009607400000000001 3.3 0.00096084 0 0.0009607600000000001 0 0.00096086 3.3 0.00096078 3.3 0.00096088 0 0.0009608 0 0.0009609 3.3 0.00096082 3.3 0.00096092 0 0.00096084 0 0.00096094 3.3 0.00096086 3.3 0.00096096 0 0.00096088 0 0.00096098 3.3 0.0009609 3.3 0.0009609999999999999 0 0.00096092 0 0.0009610199999999999 3.3 0.0009609400000000001 3.3 0.00096104 0 0.0009609600000000001 0 0.00096106 3.3 0.0009609800000000001 3.3 0.00096108 0 0.000961 0 0.0009611 3.3 0.00096102 3.3 0.00096112 0 0.00096104 0 0.00096114 3.3 0.00096106 3.3 0.00096116 0 0.00096108 0 0.00096118 3.3 0.0009611 3.3 0.0009611999999999999 0 0.00096112 0 0.0009612199999999999 3.3 0.0009611400000000001 3.3 0.00096124 0 0.0009611600000000001 0 0.00096126 3.3 0.0009611800000000001 3.3 0.00096128 0 0.0009612 0 0.0009613 3.3 0.00096122 3.3 0.00096132 0 0.00096124 0 0.00096134 3.3 0.00096126 3.3 0.00096136 0 0.00096128 0 0.00096138 3.3 0.0009613 3.3 0.0009614 0 0.00096132 0 0.0009614199999999999 3.3 0.00096134 3.3 0.0009614399999999999 0 0.0009613600000000001 0 0.00096146 3.3 0.0009613800000000001 3.3 0.00096148 0 0.0009614000000000001 0 0.0009615 3.3 0.00096142 3.3 0.00096152 0 0.00096144 0 0.00096154 3.3 0.00096146 3.3 0.00096156 0 0.00096148 0 0.00096158 3.3 0.0009615 3.3 0.0009616 0 0.00096152 0 0.0009616199999999999 3.3 0.00096154 3.3 0.0009616399999999999 0 0.0009615600000000001 0 0.00096166 3.3 0.0009615800000000001 3.3 0.00096168 0 0.0009616000000000001 0 0.0009617 3.3 0.00096162 3.3 0.00096172 0 0.00096164 0 0.00096174 3.3 0.00096166 3.3 0.00096176 0 0.00096168 0 0.00096178 3.3 0.0009617 3.3 0.0009618 0 0.00096172 0 0.00096182 3.3 0.00096174 3.3 0.0009618399999999999 0 0.00096176 0 0.0009618599999999999 3.3 0.0009617800000000001 3.3 0.00096188 0 0.0009618000000000001 0 0.0009619 3.3 0.0009618200000000001 3.3 0.00096192 0 0.00096184 0 0.00096194 3.3 0.00096186 3.3 0.00096196 0 0.00096188 0 0.00096198 3.3 0.0009619 3.3 0.000962 0 0.00096192 0 0.00096202 3.3 0.00096194 3.3 0.0009620399999999999 0 0.00096196 0 0.0009620599999999999 3.3 0.0009619800000000001 3.3 0.00096208 0 0.0009620000000000001 0 0.0009621 3.3 0.0009620200000000001 3.3 0.00096212 0 0.00096204 0 0.00096214 3.3 0.00096206 3.3 0.00096216 0 0.00096208 0 0.00096218 3.3 0.0009621 3.3 0.0009622 0 0.00096212 0 0.00096222 3.3 0.00096214 3.3 0.00096224 0 0.00096216 0 0.0009622599999999999 3.3 0.00096218 3.3 0.0009622799999999999 0 0.0009622000000000001 0 0.0009623 3.3 0.0009622200000000001 3.3 0.00096232 0 0.0009622400000000001 0 0.00096234 3.3 0.00096226 3.3 0.00096236 0 0.00096228 0 0.00096238 3.3 0.0009623 3.3 0.0009624 0 0.00096232 0 0.00096242 3.3 0.00096234 3.3 0.00096244 0 0.00096236 0 0.0009624599999999999 3.3 0.00096238 3.3 0.0009624799999999999 0 0.0009624000000000001 0 0.0009625 3.3 0.0009624200000000001 3.3 0.00096252 0 0.0009624400000000001 0 0.00096254 3.3 0.00096246 3.3 0.00096256 0 0.00096248 0 0.00096258 3.3 0.0009625 3.3 0.0009626 0 0.00096252 0 0.00096262 3.3 0.00096254 3.3 0.00096264 0 0.00096256 0 0.00096266 3.3 0.00096258 3.3 0.0009626799999999999 0 0.0009626 0 0.0009626999999999999 3.3 0.0009626200000000001 3.3 0.00096272 0 0.0009626400000000001 0 0.00096274 3.3 0.0009626600000000001 3.3 0.00096276 0 0.00096268 0 0.00096278 3.3 0.0009627 3.3 0.0009628 0 0.00096272 0 0.00096282 3.3 0.00096274 3.3 0.00096284 0 0.00096276 0 0.00096286 3.3 0.00096278 3.3 0.0009628799999999999 0 0.0009628 0 0.0009628999999999999 3.3 0.0009628200000000001 3.3 0.00096292 0 0.0009628400000000001 0 0.00096294 3.3 0.0009628600000000001 3.3 0.00096296 0 0.00096288 0 0.00096298 3.3 0.0009629 3.3 0.000963 0 0.00096292 0 0.00096302 3.3 0.00096294 3.3 0.00096304 0 0.00096296 0 0.00096306 3.3 0.00096298 3.3 0.00096308 0 0.000963 0 0.0009630999999999999 3.3 0.00096302 3.3 0.0009631199999999999 0 0.0009630400000000001 0 0.00096314 3.3 0.0009630600000000001 3.3 0.00096316 0 0.0009630800000000001 0 0.00096318 3.3 0.0009631 3.3 0.0009632 0 0.00096312 0 0.00096322 3.3 0.00096314 3.3 0.00096324 0 0.00096316 0 0.00096326 3.3 0.00096318 3.3 0.00096328 0 0.0009632 0 0.0009632999999999999 3.3 0.00096322 3.3 0.0009633199999999999 0 0.0009632400000000001 0 0.00096334 3.3 0.0009632600000000001 3.3 0.00096336 0 0.0009632800000000001 0 0.00096338 3.3 0.0009633 3.3 0.0009634 0 0.00096332 0 0.00096342 3.3 0.00096334 3.3 0.00096344 0 0.00096336 0 0.00096346 3.3 0.00096338 3.3 0.00096348 0 0.0009634 0 0.0009635 3.3 0.00096342 3.3 0.0009635199999999999 0 0.0009634400000000001 0 0.00096354 3.3 0.0009634600000000001 3.3 0.00096356 0 0.0009634800000000001 0 0.00096358 3.3 0.0009635000000000001 3.3 0.0009636 0 0.00096352 0 0.00096362 3.3 0.00096354 3.3 0.00096364 0 0.00096356 0 0.00096366 3.3 0.00096358 3.3 0.00096368 0 0.0009636 0 0.0009637 3.3 0.00096362 3.3 0.0009637199999999999 0 0.00096364 0 0.0009637399999999999 3.3 0.0009636600000000001 3.3 0.00096376 0 0.0009636800000000001 0 0.00096378 3.3 0.0009637000000000001 3.3 0.0009638 0 0.00096372 0 0.00096382 3.3 0.00096374 3.3 0.00096384 0 0.00096376 0 0.00096386 3.3 0.00096378 3.3 0.00096388 0 0.0009638 0 0.0009639 3.3 0.00096382 3.3 0.00096392 0 0.00096384 0 0.0009639399999999999 3.3 0.0009638600000000001 3.3 0.00096396 0 0.0009638800000000001 0 0.00096398 3.3 0.0009639000000000001 3.3 0.000964 0 0.0009639200000000001 0 0.00096402 3.3 0.00096394 3.3 0.00096404 0 0.00096396 0 0.00096406 3.3 0.00096398 3.3 0.00096408 0 0.000964 0 0.0009641 3.3 0.00096402 3.3 0.00096412 0 0.00096404 0 0.0009641399999999999 3.3 0.00096406 3.3 0.0009641599999999999 0 0.0009640800000000001 0 0.00096418 3.3 0.0009641000000000001 3.3 0.0009642 0 0.0009641200000000001 0 0.00096422 3.3 0.00096414 3.3 0.00096424 0 0.00096416 0 0.00096426 3.3 0.00096418 3.3 0.00096428 0 0.0009642 0 0.0009643 3.3 0.00096422 3.3 0.00096432 0 0.00096424 0 0.0009643399999999999 3.3 0.00096426 3.3 0.0009643599999999999 0 0.0009642800000000001 0 0.00096438 3.3 0.0009643000000000001 3.3 0.0009644 0 0.0009643200000000001 0 0.00096442 3.3 0.00096434 3.3 0.00096444 0 0.00096436 0 0.00096446 3.3 0.00096438 3.3 0.00096448 0 0.0009644 0 0.0009645 3.3 0.00096442 3.3 0.00096452 0 0.00096444 0 0.00096454 3.3 0.00096446 3.3 0.0009645599999999999 0 0.00096448 0 0.0009645799999999999 3.3 0.0009645000000000001 3.3 0.0009646 0 0.0009645200000000001 0 0.00096462 3.3 0.0009645400000000001 3.3 0.00096464 0 0.00096456 0 0.00096466 3.3 0.00096458 3.3 0.00096468 0 0.0009646 0 0.0009647 3.3 0.00096462 3.3 0.00096472 0 0.00096464 0 0.00096474 3.3 0.00096466 3.3 0.0009647599999999999 0 0.00096468 0 0.0009647799999999999 3.3 0.0009647000000000001 3.3 0.0009648 0 0.0009647200000000001 0 0.00096482 3.3 0.0009647400000000001 3.3 0.00096484 0 0.00096476 0 0.00096486 3.3 0.00096478 3.3 0.00096488 0 0.0009648 0 0.0009649 3.3 0.00096482 3.3 0.00096492 0 0.00096484 0 0.00096494 3.3 0.00096486 3.3 0.00096496 0 0.00096488 0 0.0009649799999999999 3.3 0.0009649 3.3 0.0009649999999999999 0 0.0009649200000000001 0 0.00096502 3.3 0.0009649400000000001 3.3 0.00096504 0 0.0009649600000000001 0 0.00096506 3.3 0.00096498 3.3 0.00096508 0 0.000965 0 0.0009651 3.3 0.00096502 3.3 0.00096512 0 0.00096504 0 0.00096514 3.3 0.00096506 3.3 0.00096516 0 0.00096508 0 0.0009651799999999999 3.3 0.0009651 3.3 0.0009651999999999999 0 0.0009651200000000001 0 0.00096522 3.3 0.0009651400000000001 3.3 0.00096524 0 0.0009651600000000001 0 0.00096526 3.3 0.00096518 3.3 0.00096528 0 0.0009652 0 0.0009653 3.3 0.00096522 3.3 0.00096532 0 0.00096524 0 0.00096534 3.3 0.00096526 3.3 0.00096536 0 0.00096528 0 0.00096538 3.3 0.0009653 3.3 0.0009653999999999999 0 0.00096532 0 0.0009654199999999999 3.3 0.0009653400000000001 3.3 0.00096544 0 0.0009653600000000001 0 0.00096546 3.3 0.0009653800000000001 3.3 0.00096548 0 0.0009654 0 0.0009655 3.3 0.00096542 3.3 0.00096552 0 0.00096544 0 0.00096554 3.3 0.00096546 3.3 0.00096556 0 0.00096548 0 0.00096558 3.3 0.0009655 3.3 0.0009655999999999999 0 0.00096552 0 0.0009656199999999999 3.3 0.0009655400000000001 3.3 0.00096564 0 0.0009655600000000001 0 0.00096566 3.3 0.0009655800000000001 3.3 0.00096568 0 0.0009656 0 0.0009657 3.3 0.00096562 3.3 0.00096572 0 0.00096564 0 0.00096574 3.3 0.00096566 3.3 0.00096576 0 0.00096568 0 0.00096578 3.3 0.0009657 3.3 0.0009658 0 0.00096572 0 0.0009658199999999999 3.3 0.00096574 3.3 0.0009658399999999999 0 0.0009657600000000001 0 0.00096586 3.3 0.0009657800000000001 3.3 0.00096588 0 0.0009658000000000001 0 0.0009659 3.3 0.00096582 3.3 0.00096592 0 0.00096584 0 0.00096594 3.3 0.00096586 3.3 0.00096596 0 0.00096588 0 0.00096598 3.3 0.0009659 3.3 0.000966 0 0.00096592 0 0.0009660199999999999 3.3 0.00096594 3.3 0.0009660399999999999 0 0.0009659600000000001 0 0.00096606 3.3 0.0009659800000000001 3.3 0.00096608 0 0.0009660000000000001 0 0.0009661 3.3 0.00096602 3.3 0.00096612 0 0.00096604 0 0.00096614 3.3 0.00096606 3.3 0.00096616 0 0.00096608 0 0.00096618 3.3 0.0009661 3.3 0.0009662 0 0.00096612 0 0.00096622 3.3 0.00096614 3.3 0.0009662399999999999 0 0.00096616 0 0.0009662599999999999 3.3 0.0009661800000000001 3.3 0.00096628 0 0.0009662000000000001 0 0.0009663 3.3 0.0009662200000000001 3.3 0.00096632 0 0.00096624 0 0.00096634 3.3 0.00096626 3.3 0.00096636 0 0.00096628 0 0.00096638 3.3 0.0009663 3.3 0.0009664 0 0.00096632 0 0.00096642 3.3 0.00096634 3.3 0.0009664399999999999 0 0.00096636 0 0.0009664599999999999 3.3 0.0009663800000000001 3.3 0.00096648 0 0.0009664000000000001 0 0.0009665 3.3 0.0009664200000000001 3.3 0.00096652 0 0.00096644 0 0.00096654 3.3 0.00096646 3.3 0.00096656 0 0.00096648 0 0.00096658 3.3 0.0009665 3.3 0.0009666 0 0.00096652 0 0.00096662 3.3 0.00096654 3.3 0.00096664 0 0.00096656 0 0.0009666599999999999 3.3 0.00096658 3.3 0.0009666799999999999 0 0.0009666000000000001 0 0.0009667 3.3 0.0009666200000000001 3.3 0.00096672 0 0.0009666400000000001 0 0.00096674 3.3 0.00096666 3.3 0.00096676 0 0.00096668 0 0.00096678 3.3 0.0009667 3.3 0.0009668 0 0.00096672 0 0.00096682 3.3 0.00096674 3.3 0.00096684 0 0.00096676 0 0.0009668599999999999 3.3 0.00096678 3.3 0.0009668799999999999 0 0.0009668000000000001 0 0.0009669 3.3 0.0009668200000000001 3.3 0.00096692 0 0.0009668400000000001 0 0.00096694 3.3 0.00096686 3.3 0.00096696 0 0.00096688 0 0.00096698 3.3 0.0009669 3.3 0.000967 0 0.00096692 0 0.00096702 3.3 0.00096694 3.3 0.00096704 0 0.00096696 0 0.00096706 3.3 0.00096698 3.3 0.0009670799999999999 0 0.0009670000000000001 0 0.0009671 3.3 0.0009670200000000001 3.3 0.00096712 0 0.0009670400000000001 0 0.00096714 3.3 0.0009670600000000001 3.3 0.00096716 0 0.00096708 0 0.00096718 3.3 0.0009671 3.3 0.0009672 0 0.00096712 0 0.00096722 3.3 0.00096714 3.3 0.00096724 0 0.00096716 0 0.00096726 3.3 0.00096718 3.3 0.0009672799999999999 0 0.0009672 0 0.0009672999999999999 3.3 0.0009672200000000001 3.3 0.00096732 0 0.0009672400000000001 0 0.00096734 3.3 0.0009672600000000001 3.3 0.00096736 0 0.00096728 0 0.00096738 3.3 0.0009673 3.3 0.0009674 0 0.00096732 0 0.00096742 3.3 0.00096734 3.3 0.00096744 0 0.00096736 0 0.00096746 3.3 0.00096738 3.3 0.00096748 0 0.0009674 0 0.0009674999999999999 3.3 0.0009674200000000001 3.3 0.00096752 0 0.0009674400000000001 0 0.00096754 3.3 0.0009674600000000001 3.3 0.00096756 0 0.0009674800000000001 0 0.00096758 3.3 0.0009675 3.3 0.0009676 0 0.00096752 0 0.00096762 3.3 0.00096754 3.3 0.00096764 0 0.00096756 0 0.00096766 3.3 0.00096758 3.3 0.00096768 0 0.0009676 0 0.0009676999999999999 3.3 0.00096762 3.3 0.0009677199999999999 0 0.0009676400000000001 0 0.00096774 3.3 0.0009676600000000001 3.3 0.00096776 0 0.0009676800000000001 0 0.00096778 3.3 0.0009677 3.3 0.0009678 0 0.00096772 0 0.00096782 3.3 0.00096774 3.3 0.00096784 0 0.00096776 0 0.00096786 3.3 0.00096778 3.3 0.00096788 0 0.0009678 0 0.0009678999999999999 3.3 0.00096782 3.3 0.0009679199999999999 0 0.0009678400000000001 0 0.00096794 3.3 0.0009678600000000001 3.3 0.00096796 0 0.0009678800000000001 0 0.00096798 3.3 0.0009679 3.3 0.000968 0 0.00096792 0 0.00096802 3.3 0.00096794 3.3 0.00096804 0 0.00096796 0 0.00096806 3.3 0.00096798 3.3 0.00096808 0 0.000968 0 0.0009681 3.3 0.00096802 3.3 0.0009681199999999999 0 0.00096804 0 0.0009681399999999999 3.3 0.0009680600000000001 3.3 0.00096816 0 0.0009680800000000001 0 0.00096818 3.3 0.0009681000000000001 3.3 0.0009682 0 0.00096812 0 0.00096822 3.3 0.00096814 3.3 0.00096824 0 0.00096816 0 0.00096826 3.3 0.00096818 3.3 0.00096828 0 0.0009682 0 0.0009683 3.3 0.00096822 3.3 0.0009683199999999999 0 0.00096824 0 0.0009683399999999999 3.3 0.0009682600000000001 3.3 0.00096836 0 0.0009682800000000001 0 0.00096838 3.3 0.0009683000000000001 3.3 0.0009684 0 0.00096832 0 0.00096842 3.3 0.00096834 3.3 0.00096844 0 0.00096836 0 0.00096846 3.3 0.00096838 3.3 0.00096848 0 0.0009684 0 0.0009685 3.3 0.00096842 3.3 0.00096852 0 0.00096844 0 0.0009685399999999999 3.3 0.00096846 3.3 0.0009685599999999999 0 0.0009684800000000001 0 0.00096858 3.3 0.0009685000000000001 3.3 0.0009686 0 0.0009685200000000001 0 0.00096862 3.3 0.00096854 3.3 0.00096864 0 0.00096856 0 0.00096866 3.3 0.00096858 3.3 0.00096868 0 0.0009686 0 0.0009687 3.3 0.00096862 3.3 0.00096872 0 0.00096864 0 0.0009687399999999999 3.3 0.00096866 3.3 0.0009687599999999999 0 0.0009686800000000001 0 0.00096878 3.3 0.0009687000000000001 3.3 0.0009688 0 0.0009687200000000001 0 0.00096882 3.3 0.00096874 3.3 0.00096884 0 0.00096876 0 0.00096886 3.3 0.00096878 3.3 0.00096888 0 0.0009688 0 0.0009689 3.3 0.00096882 3.3 0.00096892 0 0.00096884 0 0.00096894 3.3 0.00096886 3.3 0.0009689599999999999 0 0.00096888 0 0.0009689799999999999 3.3 0.0009689000000000001 3.3 0.000969 0 0.0009689200000000001 0 0.00096902 3.3 0.0009689400000000001 3.3 0.00096904 0 0.00096896 0 0.00096906 3.3 0.00096898 3.3 0.00096908 0 0.000969 0 0.0009691 3.3 0.00096902 3.3 0.00096912 0 0.00096904 0 0.00096914 3.3 0.00096906 3.3 0.0009691599999999999 0 0.00096908 0 0.0009691799999999999 3.3 0.0009691000000000001 3.3 0.0009692 0 0.0009691200000000001 0 0.00096922 3.3 0.0009691400000000001 3.3 0.00096924 0 0.00096916 0 0.00096926 3.3 0.00096918 3.3 0.00096928 0 0.0009692 0 0.0009693 3.3 0.00096922 3.3 0.00096932 0 0.00096924 0 0.00096934 3.3 0.00096926 3.3 0.00096936 0 0.00096928 0 0.0009693799999999999 3.3 0.0009693 3.3 0.0009693999999999999 0 0.0009693200000000001 0 0.00096942 3.3 0.0009693400000000001 3.3 0.00096944 0 0.0009693600000000001 0 0.00096946 3.3 0.00096938 3.3 0.00096948 0 0.0009694 0 0.0009695 3.3 0.00096942 3.3 0.00096952 0 0.00096944 0 0.00096954 3.3 0.00096946 3.3 0.00096956 0 0.00096948 0 0.0009695799999999999 3.3 0.0009695 3.3 0.0009695999999999999 0 0.0009695200000000001 0 0.00096962 3.3 0.0009695400000000001 3.3 0.00096964 0 0.0009695600000000001 0 0.00096966 3.3 0.00096958 3.3 0.00096968 0 0.0009696 0 0.0009697 3.3 0.00096962 3.3 0.00096972 0 0.00096964 0 0.00096974 3.3 0.00096966 3.3 0.00096976 0 0.00096968 0 0.00096978 3.3 0.0009697 3.3 0.0009697999999999999 0 0.00096972 0 0.0009698199999999999 3.3 0.0009697400000000001 3.3 0.00096984 0 0.0009697600000000001 0 0.00096986 3.3 0.0009697800000000001 3.3 0.00096988 0 0.0009698 0 0.0009699 3.3 0.00096982 3.3 0.00096992 0 0.00096984 0 0.00096994 3.3 0.00096986 3.3 0.00096996 0 0.00096988 0 0.00096998 3.3 0.0009699 3.3 0.0009699999999999999 0 0.00096992 0 0.0009700199999999999 3.3 0.0009699400000000001 3.3 0.00097004 0 0.0009699600000000001 0 0.00097006 3.3 0.0009699800000000001 3.3 0.00097008 0 0.00097 0 0.0009701 3.3 0.00097002 3.3 0.00097012 0 0.00097004 0 0.00097014 3.3 0.00097006 3.3 0.00097016 0 0.00097008 0 0.00097018 3.3 0.0009701 3.3 0.0009702 0 0.00097012 0 0.0009702199999999999 3.3 0.00097014 3.3 0.0009702399999999999 0 0.0009701600000000001 0 0.00097026 3.3 0.0009701800000000001 3.3 0.00097028 0 0.0009702000000000001 0 0.0009703 3.3 0.00097022 3.3 0.00097032 0 0.00097024 0 0.00097034 3.3 0.00097026 3.3 0.00097036 0 0.00097028 0 0.00097038 3.3 0.0009703 3.3 0.0009704 0 0.00097032 0 0.0009704199999999999 3.3 0.00097034 3.3 0.0009704399999999999 0 0.0009703600000000001 0 0.00097046 3.3 0.0009703800000000001 3.3 0.00097048 0 0.0009704000000000001 0 0.0009705 3.3 0.00097042 3.3 0.00097052 0 0.00097044 0 0.00097054 3.3 0.00097046 3.3 0.00097056 0 0.00097048 0 0.00097058 3.3 0.0009705 3.3 0.0009706 0 0.00097052 0 0.00097062 3.3 0.00097054 3.3 0.0009706399999999999 0 0.0009705600000000001 0 0.00097066 3.3 0.0009705800000000001 3.3 0.00097068 0 0.0009706000000000001 0 0.0009707 3.3 0.0009706200000000001 3.3 0.00097072 0 0.00097064 0 0.00097074 3.3 0.00097066 3.3 0.00097076 0 0.00097068 0 0.00097078 3.3 0.0009707 3.3 0.0009708 0 0.00097072 0 0.00097082 3.3 0.00097074 3.3 0.0009708399999999999 0 0.00097076 0 0.0009708599999999999 3.3 0.0009707800000000001 3.3 0.00097088 0 0.0009708000000000001 0 0.0009709 3.3 0.0009708200000000001 3.3 0.00097092 0 0.00097084 0 0.00097094 3.3 0.00097086 3.3 0.00097096 0 0.00097088 0 0.00097098 3.3 0.0009709 3.3 0.000971 0 0.00097092 0 0.00097102 3.3 0.00097094 3.3 0.0009710399999999999 0 0.00097096 0 0.0009710599999999999 3.3 0.0009709800000000001 3.3 0.00097108 0 0.0009710000000000001 0 0.0009711 3.3 0.0009710200000000001 3.3 0.00097112 0 0.00097104 0 0.00097114 3.3 0.00097106 3.3 0.00097116 0 0.00097108 0 0.00097118 3.3 0.0009711 3.3 0.0009712 0 0.00097112 0 0.00097122 3.3 0.00097114 3.3 0.00097124 0 0.00097116 0 0.0009712599999999999 3.3 0.00097118 3.3 0.0009712799999999999 0 0.0009712000000000001 0 0.0009713 3.3 0.0009712200000000001 3.3 0.00097132 0 0.0009712400000000001 0 0.00097134 3.3 0.00097126 3.3 0.00097136 0 0.00097128 0 0.00097138 3.3 0.0009713 3.3 0.0009714 0 0.00097132 0 0.00097142 3.3 0.00097134 3.3 0.00097144 0 0.00097136 0 0.0009714599999999999 3.3 0.00097138 3.3 0.0009714799999999999 0 0.0009714000000000001 0 0.0009715 3.3 0.0009714200000000001 3.3 0.00097152 0 0.0009714400000000001 0 0.00097154 3.3 0.00097146 3.3 0.00097156 0 0.00097148 0 0.00097158 3.3 0.0009715 3.3 0.0009716 0 0.00097152 0 0.00097162 3.3 0.00097154 3.3 0.00097164 0 0.00097156 0 0.00097166 3.3 0.00097158 3.3 0.0009716799999999999 0 0.0009716 0 0.0009716999999999999 3.3 0.0009716200000000001 3.3 0.00097172 0 0.0009716400000000001 0 0.00097174 3.3 0.0009716600000000001 3.3 0.00097176 0 0.00097168 0 0.00097178 3.3 0.0009717 3.3 0.0009718 0 0.00097172 0 0.00097182 3.3 0.00097174 3.3 0.00097184 0 0.00097176 0 0.00097186 3.3 0.00097178 3.3 0.0009718799999999999 0 0.0009718 0 0.0009718999999999999 3.3 0.0009718200000000001 3.3 0.00097192 0 0.0009718400000000001 0 0.00097194 3.3 0.0009718600000000001 3.3 0.00097196 0 0.00097188 0 0.00097198 3.3 0.0009719 3.3 0.000972 0 0.00097192 0 0.00097202 3.3 0.00097194 3.3 0.00097204 0 0.00097196 0 0.00097206 3.3 0.00097198 3.3 0.00097208 0 0.000972 0 0.0009720999999999999 3.3 0.00097202 3.3 0.0009721199999999999 0 0.0009720400000000001 0 0.00097214 3.3 0.0009720600000000001 3.3 0.00097216 0 0.0009720800000000001 0 0.00097218 3.3 0.0009721 3.3 0.0009722 0 0.00097212 0 0.00097222 3.3 0.00097214 3.3 0.00097224 0 0.00097216 0 0.00097226 3.3 0.00097218 3.3 0.00097228 0 0.0009722 0 0.0009722999999999999 3.3 0.00097222 3.3 0.0009723199999999999 0 0.0009722400000000001 0 0.00097234 3.3 0.0009722600000000001 3.3 0.00097236 0 0.0009722800000000001 0 0.00097238 3.3 0.0009723 3.3 0.0009724 0 0.00097232 0 0.00097242 3.3 0.00097234 3.3 0.00097244 0 0.00097236 0 0.00097246 3.3 0.00097238 3.3 0.00097248 0 0.0009724 0 0.0009725 3.3 0.00097242 3.3 0.0009725199999999999 0 0.00097244 0 0.0009725399999999999 3.3 0.0009724600000000001 3.3 0.00097256 0 0.0009724800000000001 0 0.00097258 3.3 0.0009725000000000001 3.3 0.0009726 0 0.00097252 0 0.00097262 3.3 0.00097254 3.3 0.00097264 0 0.00097256 0 0.00097266 3.3 0.00097258 3.3 0.00097268 0 0.0009726 0 0.0009727 3.3 0.00097262 3.3 0.0009727199999999999 0 0.00097264 0 0.0009727399999999999 3.3 0.0009726600000000001 3.3 0.00097276 0 0.0009726800000000001 0 0.00097278 3.3 0.0009727000000000001 3.3 0.0009728 0 0.00097272 0 0.00097282 3.3 0.00097274 3.3 0.00097284 0 0.00097276 0 0.00097286 3.3 0.00097278 3.3 0.00097288 0 0.0009728 0 0.0009729 3.3 0.00097282 3.3 0.00097292 0 0.00097284 0 0.0009729399999999999 3.3 0.00097286 3.3 0.0009729599999999999 0 0.0009728800000000001 0 0.00097298 3.3 0.0009729000000000001 3.3 0.000973 0 0.0009729200000000001 0 0.00097302 3.3 0.00097294 3.3 0.00097304 0 0.00097296 0 0.00097306 3.3 0.00097298 3.3 0.00097308 0 0.000973 0 0.0009731 3.3 0.00097302 3.3 0.00097312 0 0.00097304 0 0.0009731399999999999 3.3 0.00097306 3.3 0.0009731599999999999 0 0.0009730800000000001 0 0.00097318 3.3 0.0009731000000000001 3.3 0.0009732 0 0.0009731200000000001 0 0.00097322 3.3 0.00097314 3.3 0.00097324 0 0.00097316 0 0.00097326 3.3 0.00097318 3.3 0.00097328 0 0.0009732 0 0.0009733 3.3 0.00097322 3.3 0.00097332 0 0.00097324 0 0.00097334 3.3 0.00097326 3.3 0.0009733599999999999 0 0.00097328 0 0.0009733799999999999 3.3 0.0009733000000000001 3.3 0.0009734 0 0.0009733200000000001 0 0.00097342 3.3 0.0009733400000000001 3.3 0.00097344 0 0.00097336 0 0.00097346 3.3 0.00097338 3.3 0.00097348 0 0.0009734 0 0.0009735 3.3 0.00097342 3.3 0.00097352 0 0.00097344 0 0.00097354 3.3 0.00097346 3.3 0.0009735599999999999 0 0.00097348 0 0.0009735799999999999 3.3 0.0009735000000000001 3.3 0.0009736 0 0.0009735200000000001 0 0.00097362 3.3 0.0009735400000000001 3.3 0.00097364 0 0.00097356 0 0.00097366 3.3 0.00097358 3.3 0.00097368 0 0.0009736 0 0.0009737 3.3 0.00097362 3.3 0.00097372 0 0.00097364 0 0.00097374 3.3 0.00097366 3.3 0.00097376 0 0.00097368 0 0.0009737799999999999 3.3 0.0009737000000000001 3.3 0.0009738 0 0.0009737200000000001 0 0.00097382 3.3 0.0009737400000000001 3.3 0.00097384 0 0.0009737600000000001 0 0.00097386 3.3 0.00097378 3.3 0.00097388 0 0.0009738 0 0.0009739 3.3 0.00097382 3.3 0.00097392 0 0.00097384 0 0.00097394 3.3 0.00097386 3.3 0.00097396 0 0.00097388 0 0.0009739799999999999 3.3 0.0009739 3.3 0.0009739999999999999 0 0.0009739200000000001 0 0.00097402 3.3 0.0009739400000000001 3.3 0.00097404 0 0.0009739600000000001 0 0.00097406 3.3 0.00097398 3.3 0.00097408 0 0.000974 0 0.0009741 3.3 0.00097402 3.3 0.00097412 0 0.00097404 0 0.00097414 3.3 0.00097406 3.3 0.00097416 0 0.00097408 0 0.00097418 3.3 0.0009741 3.3 0.0009741999999999999 0 0.0009741200000000001 0 0.00097422 3.3 0.0009741400000000001 3.3 0.00097424 0 0.0009741600000000001 0 0.00097426 3.3 0.0009741800000000001 3.3 0.00097428 0 0.0009742 0 0.0009743 3.3 0.00097422 3.3 0.00097432 0 0.00097424 0 0.00097434 3.3 0.00097426 3.3 0.00097436 0 0.00097428 0 0.00097438 3.3 0.0009743 3.3 0.0009743999999999999 0 0.00097432 0 0.0009744199999999999 3.3 0.0009743400000000001 3.3 0.00097444 0 0.0009743600000000001 0 0.00097446 3.3 0.0009743800000000001 3.3 0.00097448 0 0.0009744 0 0.0009745 3.3 0.00097442 3.3 0.00097452 0 0.00097444 0 0.00097454 3.3 0.00097446 3.3 0.00097456 0 0.00097448 0 0.00097458 3.3 0.0009745 3.3 0.0009745999999999999 0 0.00097452 0 0.0009746199999999999 3.3 0.0009745400000000001 3.3 0.00097464 0 0.0009745600000000001 0 0.00097466 3.3 0.0009745800000000001 3.3 0.00097468 0 0.0009746 0 0.0009747 3.3 0.00097462 3.3 0.00097472 0 0.00097464 0 0.00097474 3.3 0.00097466 3.3 0.00097476 0 0.00097468 0 0.00097478 3.3 0.0009747 3.3 0.0009748 0 0.00097472 0 0.0009748199999999999 3.3 0.00097474 3.3 0.0009748399999999999 0 0.0009747600000000001 0 0.00097486 3.3 0.0009747800000000001 3.3 0.00097488 0 0.0009748000000000001 0 0.0009749 3.3 0.00097482 3.3 0.00097492 0 0.00097484 0 0.00097494 3.3 0.00097486 3.3 0.00097496 0 0.00097488 0 0.00097498 3.3 0.0009749 3.3 0.000975 0 0.00097492 0 0.0009750199999999999 3.3 0.00097494 3.3 0.0009750399999999999 0 0.0009749600000000001 0 0.00097506 3.3 0.0009749800000000001 3.3 0.00097508 0 0.0009750000000000001 0 0.0009751 3.3 0.00097502 3.3 0.00097512 0 0.00097504 0 0.00097514 3.3 0.00097506 3.3 0.00097516 0 0.00097508 0 0.00097518 3.3 0.0009751 3.3 0.0009752 0 0.00097512 0 0.00097522 3.3 0.00097514 3.3 0.0009752399999999999 0 0.00097516 0 0.0009752599999999999 3.3 0.0009751800000000001 3.3 0.00097528 0 0.0009752000000000001 0 0.0009753 3.3 0.0009752200000000001 3.3 0.00097532 0 0.00097524 0 0.00097534 3.3 0.00097526 3.3 0.00097536 0 0.00097528 0 0.00097538 3.3 0.0009753 3.3 0.0009754 0 0.00097532 0 0.00097542 3.3 0.00097534 3.3 0.0009754399999999999 0 0.00097536 0 0.0009754599999999999 3.3 0.0009753800000000001 3.3 0.00097548 0 0.0009754000000000001 0 0.0009755 3.3 0.0009754200000000001 3.3 0.00097552 0 0.00097544 0 0.00097554 3.3 0.00097546 3.3 0.00097556 0 0.00097548 0 0.00097558 3.3 0.0009755 3.3 0.0009756 0 0.00097552 0 0.00097562 3.3 0.00097554 3.3 0.00097564 0 0.00097556 0 0.0009756599999999999 3.3 0.00097558 3.3 0.0009756799999999999 0 0.0009756000000000001 0 0.0009757 3.3 0.0009756200000000001 3.3 0.00097572 0 0.0009756400000000001 0 0.00097574 3.3 0.00097566 3.3 0.00097576 0 0.00097568 0 0.00097578 3.3 0.0009757 3.3 0.0009758 0 0.00097572 0 0.00097582 3.3 0.00097574 3.3 0.00097584 0 0.00097576 0 0.0009758599999999999 3.3 0.00097578 3.3 0.0009758799999999999 0 0.0009758000000000001 0 0.0009759 3.3 0.0009758200000000001 3.3 0.00097592 0 0.0009758400000000001 0 0.00097594 3.3 0.00097586 3.3 0.00097596 0 0.00097588 0 0.00097598 3.3 0.0009759 3.3 0.000976 0 0.00097592 0 0.00097602 3.3 0.00097594 3.3 0.00097604 0 0.00097596 0 0.00097606 3.3 0.00097598 3.3 0.0009760799999999999 0 0.000976 0 0.0009760999999999999 3.3 0.0009760200000000001 3.3 0.00097612 0 0.0009760400000000001 0 0.00097614 3.3 0.0009760600000000001 3.3 0.00097616 0 0.00097608 0 0.00097618 3.3 0.0009761 3.3 0.0009762 0 0.00097612 0 0.00097622 3.3 0.00097614 3.3 0.00097624 0 0.00097616 0 0.00097626 3.3 0.00097618 3.3 0.0009762799999999999 0 0.0009762 0 0.0009762999999999999 3.3 0.0009762200000000001 3.3 0.00097632 0 0.0009762400000000001 0 0.00097634 3.3 0.0009762600000000001 3.3 0.00097636 0 0.00097628 0 0.00097638 3.3 0.0009763 3.3 0.0009764 0 0.00097632 0 0.00097642 3.3 0.00097634 3.3 0.00097644 0 0.00097636 0 0.00097646 3.3 0.00097638 3.3 0.00097648 0 0.0009764 0 0.0009764999999999999 3.3 0.00097642 3.3 0.0009765199999999999 0 0.0009764400000000001 0 0.00097654 3.3 0.0009764600000000001 3.3 0.00097656 0 0.00097648 0 0.00097658 3.3 0.0009765 3.3 0.0009766 0 0.0009765199999999999 0 0.0009766199999999999 3.3 0.00097654 3.3 0.00097664 0 0.0009765600000000001 0 0.00097666 3.3 0.00097658 3.3 0.00097668 0 0.0009766 0 0.0009767 3.3 0.0009766199999999999 3.3 0.00097672 0 0.00097664 0 0.00097674 3.3 0.0009766599999999999 3.3 0.00097676 0 0.00097668 0 0.00097678 3.3 0.0009766999999999998 3.3 0.0009767999999999999 0 0.00097672 0 0.00097682 3.3 0.00097674 3.3 0.00097684 0 0.00097676 0 0.00097686 3.3 0.00097678 3.3 0.00097688 0 0.0009767999999999999 0 0.0009769 3.3 0.00097682 3.3 0.00097692 0 0.0009768399999999999 0 0.00097694 3.3 0.00097686 3.3 0.00097696 0 0.0009768799999999998 0 0.00097698 3.3 0.0009769 3.3 0.000977 0 0.0009769199999999998 0 0.0009770199999999999 3.3 0.00097694 3.3 0.00097704 0 0.00097696 0 0.00097706 3.3 0.00097698 3.3 0.00097708 0 0.000977 0 0.0009771 3.3 0.0009770199999999999 3.3 0.00097712 0 0.00097704 0 0.00097714 3.3 0.0009770599999999999 3.3 0.00097716 0 0.00097708 0 0.00097718 3.3 0.0009770999999999998 3.3 0.0009772 0 0.00097712 0 0.00097722 3.3 0.0009771399999999998 3.3 0.0009772399999999999 0 0.00097716 0 0.00097726 3.3 0.00097718 3.3 0.00097728 0 0.0009772 0 0.0009773 3.3 0.00097722 3.3 0.00097732 0 0.0009772399999999999 0 0.00097734 3.3 0.00097726 3.3 0.00097736 0 0.0009772799999999999 0 0.00097738 3.3 0.0009773 3.3 0.0009774 0 0.0009773199999999998 0 0.00097742 3.3 0.00097734 3.3 0.00097744 0 0.0009773599999999998 0 0.0009774599999999999 3.3 0.00097738 3.3 0.00097748 0 0.0009774 0 0.0009775 3.3 0.00097742 3.3 0.00097752 0 0.00097744 0 0.00097754 3.3 0.0009774599999999999 3.3 0.00097756 0 0.00097748 0 0.00097758 3.3 0.0009774999999999999 3.3 0.0009776 0 0.00097752 0 0.00097762 3.3 0.0009775399999999998 3.3 0.0009776399999999999 0 0.00097756 0 0.00097766 3.3 0.00097758 3.3 0.00097768 0 0.0009776 0 0.0009777 3.3 0.00097762 3.3 0.00097772 0 0.0009776399999999999 0 0.00097774 3.3 0.00097766 3.3 0.00097776 0 0.0009776799999999999 0 0.00097778 3.3 0.0009777 3.3 0.0009778 0 0.0009777199999999998 0 0.00097782 3.3 0.00097774 3.3 0.00097784 0 0.0009777599999999998 0 0.0009778599999999999 3.3 0.00097778 3.3 0.00097788 0 0.0009778 0 0.0009779 3.3 0.00097782 3.3 0.00097792 0 0.00097784 0 0.00097794 3.3 0.0009778599999999999 3.3 0.00097796 0 0.00097788 0 0.00097798 3.3 0.0009778999999999999 3.3 0.000978 0 0.00097792 0 0.00097802 3.3 0.0009779399999999998 3.3 0.00097804 0 0.00097796 0 0.00097806 3.3 0.0009779799999999998 3.3 0.0009780799999999999 0 0.000978 0 0.0009781 3.3 0.00097802 3.3 0.00097812 0 0.00097804 0 0.00097814 3.3 0.00097806 3.3 0.00097816 0 0.0009780799999999999 0 0.00097818 3.3 0.0009781 3.3 0.0009782 0 0.0009781199999999999 0 0.00097822 3.3 0.00097814 3.3 0.00097824 0 0.0009781599999999998 0 0.00097826 3.3 0.00097818 3.3 0.00097828 0 0.0009781999999999998 0 0.0009782999999999999 3.3 0.00097822 3.3 0.00097832 0 0.00097824 0 0.00097834 3.3 0.00097826 3.3 0.00097836 0 0.00097828 0 0.00097838 3.3 0.0009782999999999999 3.3 0.0009784 0 0.00097832 0 0.00097842 3.3 0.0009783399999999999 3.3 0.00097844 0 0.00097836 0 0.00097846 3.3 0.0009783799999999998 3.3 0.0009784799999999999 0 0.0009784 0 0.0009785 3.3 0.00097842 3.3 0.00097852 0 0.00097844 0 0.00097854 3.3 0.00097846 3.3 0.00097856 0 0.0009784799999999999 0 0.00097858 3.3 0.0009785 3.3 0.0009786 0 0.0009785199999999999 0 0.00097862 3.3 0.00097854 3.3 0.00097864 0 0.0009785599999999998 0 0.00097866 3.3 0.00097858 3.3 0.00097868 0 0.0009785999999999998 0 0.0009786999999999999 3.3 0.00097862 3.3 0.00097872 0 0.00097864 0 0.00097874 3.3 0.00097866 3.3 0.00097876 0 0.00097868 0 0.00097878 3.3 0.0009786999999999999 3.3 0.0009788 0 0.00097872 0 0.00097882 3.3 0.0009787399999999999 3.3 0.00097884 0 0.00097876 0 0.00097886 3.3 0.0009787799999999998 3.3 0.00097888 0 0.0009788 0 0.0009789 3.3 0.0009788199999999998 3.3 0.0009789199999999999 0 0.00097884 0 0.00097894 3.3 0.00097886 3.3 0.00097896 0 0.00097888 0 0.00097898 3.3 0.0009789 3.3 0.000979 0 0.0009789199999999999 0 0.00097902 3.3 0.00097894 3.3 0.00097904 0 0.0009789599999999999 0 0.00097906 3.3 0.00097898 3.3 0.00097908 0 0.0009789999999999998 0 0.0009791 3.3 0.00097902 3.3 0.00097912 0 0.00097904 0 0.00097914 3.3 0.00097906 3.3 0.00097916 0 0.00097908 0 0.00097918 3.3 0.0009791 3.3 0.0009792 0 0.00097912 0 0.00097922 3.3 0.0009791399999999999 3.3 0.00097924 0 0.00097916 0 0.00097926 3.3 0.0009791799999999999 3.3 0.00097928 0 0.0009792 0 0.0009793 3.3 0.0009792199999999998 3.3 0.0009793199999999999 0 0.00097924 0 0.00097934 3.3 0.00097926 3.3 0.00097936 0 0.00097928 0 0.00097938 3.3 0.0009793 3.3 0.0009794 0 0.0009793199999999999 0 0.00097942 3.3 0.00097934 3.3 0.00097944 0 0.0009793599999999999 0 0.00097946 3.3 0.00097938 3.3 0.00097948 0 0.0009793999999999998 0 0.0009795 3.3 0.00097942 3.3 0.00097952 0 0.0009794399999999998 0 0.0009795399999999999 3.3 0.00097946 3.3 0.00097956 0 0.00097948 0 0.00097958 3.3 0.0009795 3.3 0.0009796 0 0.00097952 0 0.00097962 3.3 0.0009795399999999999 3.3 0.00097964 0 0.00097956 0 0.00097966 3.3 0.0009795799999999999 3.3 0.00097968 0 0.0009796 0 0.0009797 3.3 0.0009796199999999998 3.3 0.00097972 0 0.00097964 0 0.00097974 3.3 0.0009796599999999998 3.3 0.0009797599999999999 0 0.00097968 0 0.00097978 3.3 0.0009797 3.3 0.0009798 0 0.00097972 0 0.00097982 3.3 0.00097974 3.3 0.00097984 0 0.0009797599999999999 0 0.00097986 3.3 0.00097978 3.3 0.00097988 0 0.0009797999999999999 0 0.0009799 3.3 0.00097982 3.3 0.00097992 0 0.0009798399999999998 0 0.0009799399999999999 3.3 0.00097986 3.3 0.00097996 0 0.00097988 0 0.00097998 3.3 0.0009799 3.3 0.00098 0 0.00097992 0 0.00098002 3.3 0.0009799399999999999 3.3 0.00098004 0 0.00097996 0 0.00098006 3.3 0.0009799799999999999 3.3 0.00098008 0 0.00098 0 0.0009801 3.3 0.0009800199999999998 3.3 0.00098012 0 0.00098004 0 0.00098014 3.3 0.0009800599999999998 3.3 0.0009801599999999999 0 0.00098008 0 0.00098018 3.3 0.0009801 3.3 0.0009802 0 0.00098012 0 0.00098022 3.3 0.00098014 3.3 0.00098024 0 0.0009801599999999999 0 0.00098026 3.3 0.00098018 3.3 0.00098028 0 0.0009801999999999999 0 0.0009803 3.3 0.00098022 3.3 0.00098032 0 0.0009802399999999998 0 0.00098034 3.3 0.00098026 3.3 0.00098036 0 0.0009802799999999998 0 0.0009803799999999999 3.3 0.0009803 3.3 0.0009804 0 0.00098032 0 0.00098042 3.3 0.00098034 3.3 0.00098044 0 0.00098036 0 0.00098046 3.3 0.0009803799999999999 3.3 0.00098048 0 0.0009804 0 0.0009805 3.3 0.0009804199999999999 3.3 0.00098052 0 0.00098044 0 0.00098054 3.3 0.0009804599999999998 3.3 0.00098056 0 0.00098048 0 0.00098058 3.3 0.0009804999999999998 3.3 0.0009805999999999999 0 0.00098052 0 0.00098062 3.3 0.00098054 3.3 0.00098064 0 0.00098056 0 0.00098066 3.3 0.00098058 3.3 0.00098068 0 0.0009805999999999999 0 0.0009807 3.3 0.00098062 3.3 0.00098072 0 0.0009806399999999999 0 0.00098074 3.3 0.00098066 3.3 0.00098076 0 0.0009806799999999998 0 0.0009807799999999999 3.3 0.0009807 3.3 0.0009808 0 0.00098072 0 0.00098082 3.3 0.00098074 3.3 0.00098084 0 0.00098076 0 0.00098086 3.3 0.0009807799999999999 3.3 0.00098088 0 0.0009808 0 0.0009809 3.3 0.0009808199999999999 3.3 0.00098092 0 0.00098084 0 0.00098094 3.3 0.0009808599999999998 3.3 0.00098096 0 0.00098088 0 0.00098098 3.3 0.0009808999999999998 3.3 0.0009809999999999999 0 0.00098092 0 0.00098102 3.3 0.00098094 3.3 0.00098104 0 0.00098096 0 0.00098106 3.3 0.00098098 3.3 0.00098108 0 0.0009809999999999999 0 0.0009811 3.3 0.00098102 3.3 0.00098112 0 0.0009810399999999999 0 0.00098114 3.3 0.00098106 3.3 0.00098116 0 0.0009810799999999998 0 0.00098118 3.3 0.0009811 3.3 0.0009812 0 0.0009811199999999998 0 0.0009812199999999999 3.3 0.00098114 3.3 0.00098124 0 0.00098116 0 0.00098126 3.3 0.00098118 3.3 0.00098128 0 0.0009812 0 0.0009813 3.3 0.0009812199999999999 3.3 0.00098132 0 0.00098124 0 0.00098134 3.3 0.0009812599999999999 3.3 0.00098136 0 0.00098128 0 0.00098138 3.3 0.0009812999999999998 3.3 0.0009814 0 0.00098132 0 0.00098142 3.3 0.0009813399999999998 3.3 0.0009814399999999999 0 0.00098136 0 0.00098146 3.3 0.00098138 3.3 0.00098148 0 0.0009814 0 0.0009815 3.3 0.00098142 3.3 0.00098152 0 0.0009814399999999999 0 0.00098154 3.3 0.00098146 3.3 0.00098156 0 0.0009814799999999999 0 0.00098158 3.3 0.0009815 3.3 0.0009816 0 0.0009815199999999998 0 0.0009816199999999999 3.3 0.00098154 3.3 0.00098164 0 0.00098156 0 0.00098166 3.3 0.00098158 3.3 0.00098168 0 0.0009816 0 0.0009817 3.3 0.0009816199999999999 3.3 0.00098172 0 0.00098164 0 0.00098174 3.3 0.0009816599999999999 3.3 0.00098176 0 0.00098168 0 0.00098178 3.3 0.0009816999999999998 3.3 0.0009818 0 0.00098172 0 0.00098182 3.3 0.0009817399999999998 3.3 0.0009818399999999999 0 0.00098176 0 0.00098186 3.3 0.00098178 3.3 0.00098188 0 0.0009818 0 0.0009819 3.3 0.00098182 3.3 0.00098192 0 0.0009818399999999999 0 0.00098194 3.3 0.00098186 3.3 0.00098196 0 0.0009818799999999999 0 0.00098198 3.3 0.0009819 3.3 0.000982 0 0.0009819199999999998 0 0.00098202 3.3 0.00098194 3.3 0.00098204 0 0.0009819599999999998 0 0.0009820599999999999 3.3 0.00098198 3.3 0.00098208 0 0.000982 0 0.0009821 3.3 0.00098202 3.3 0.00098212 0 0.00098204 0 0.00098214 3.3 0.0009820599999999999 3.3 0.00098216 0 0.00098208 0 0.00098218 3.3 0.0009820999999999999 3.3 0.0009822 0 0.00098212 0 0.00098222 3.3 0.0009821399999999998 3.3 0.00098224 0 0.00098216 0 0.00098226 3.3 0.0009821799999999998 3.3 0.0009822799999999999 0 0.0009822 0 0.0009823 3.3 0.00098222 3.3 0.00098232 0 0.00098224 0 0.00098234 3.3 0.00098226 3.3 0.00098236 0 0.0009822799999999999 0 0.00098238 3.3 0.0009823 3.3 0.0009824 0 0.0009823199999999999 0 0.00098242 3.3 0.00098234 3.3 0.00098244 0 0.0009823599999999998 0 0.0009824599999999999 3.3 0.00098238 3.3 0.00098248 0 0.0009824 0 0.0009825 3.3 0.00098242 3.3 0.00098252 0 0.00098244 0 0.00098254 3.3 0.0009824599999999999 3.3 0.00098256 0 0.00098248 0 0.00098258 3.3 0.0009824999999999999 3.3 0.0009826 0 0.00098252 0 0.00098262 3.3 0.0009825399999999998 3.3 0.00098264 0 0.00098256 0 0.00098266 3.3 0.0009825799999999998 3.3 0.0009826799999999999 0 0.0009826 0 0.0009827 3.3 0.00098262 3.3 0.00098272 0 0.00098264 0 0.00098274 3.3 0.00098266 3.3 0.00098276 0 0.0009826799999999999 0 0.00098278 3.3 0.0009827 3.3 0.0009828 0 0.0009827199999999999 0 0.00098282 3.3 0.00098274 3.3 0.00098284 0 0.0009827599999999998 0 0.00098286 3.3 0.00098278 3.3 0.00098288 0 0.0009827999999999998 0 0.0009828999999999999 3.3 0.00098282 3.3 0.00098292 0 0.00098284 0 0.00098294 3.3 0.00098286 3.3 0.00098296 0 0.00098288 0 0.00098298 3.3 0.0009828999999999999 3.3 0.000983 0 0.00098292 0 0.00098302 3.3 0.0009829399999999999 3.3 0.00098304 0 0.00098296 0 0.00098306 3.3 0.0009829799999999998 3.3 0.0009830799999999999 0 0.000983 0 0.0009831 3.3 0.00098302 3.3 0.00098312 0 0.00098304 0 0.00098314 3.3 0.00098306 3.3 0.00098316 0 0.0009830799999999999 0 0.00098318 3.3 0.0009831 3.3 0.0009832 0 0.0009831199999999999 0 0.00098322 3.3 0.00098314 3.3 0.00098324 0 0.0009831599999999999 0 0.00098326 3.3 0.00098318 3.3 0.00098328 0 0.0009831999999999998 0 0.0009832999999999999 3.3 0.00098322 3.3 0.00098332 0 0.00098324 0 0.00098334 3.3 0.00098326 3.3 0.00098336 0 0.00098328 0 0.00098338 3.3 0.0009832999999999999 3.3 0.0009834 0 0.00098332 0 0.00098342 3.3 0.0009833399999999999 3.3 0.00098344 0 0.00098336 0 0.00098346 3.3 0.0009833799999999998 3.3 0.00098348 0 0.0009834 0 0.0009835 3.3 0.0009834199999999998 3.3 0.0009835199999999999 0 0.00098344 0 0.00098354 3.3 0.00098346 3.3 0.00098356 0 0.00098348 0 0.00098358 3.3 0.0009835 3.3 0.0009836 0 0.0009835199999999999 0 0.00098362 3.3 0.00098354 3.3 0.00098364 0 0.0009835599999999999 0 0.00098366 3.3 0.00098358 3.3 0.00098368 0 0.0009835999999999998 0 0.0009837 3.3 0.00098362 3.3 0.00098372 0 0.0009836399999999998 0 0.0009837399999999999 3.3 0.00098366 3.3 0.00098376 0 0.00098368 0 0.00098378 3.3 0.0009837 3.3 0.0009838 0 0.00098372 0 0.00098382 3.3 0.0009837399999999999 3.3 0.00098384 0 0.00098376 0 0.00098386 3.3 0.0009837799999999999 3.3 0.00098388 0 0.0009838 0 0.0009839 3.3 0.0009838199999999998 3.3 0.0009839199999999999 0 0.00098384 0 0.00098394 3.3 0.00098386 3.3 0.00098396 0 0.00098388 0 0.00098398 3.3 0.0009839 3.3 0.000984 0 0.0009839199999999999 0 0.00098402 3.3 0.00098394 3.3 0.00098404 0 0.0009839599999999999 0 0.00098406 3.3 0.00098398 3.3 0.00098408 0 0.0009839999999999998 0 0.0009841 3.3 0.00098402 3.3 0.00098412 0 0.0009840399999999998 0 0.0009841399999999999 3.3 0.00098406 3.3 0.00098416 0 0.00098408 0 0.00098418 3.3 0.0009841 3.3 0.0009842 0 0.00098412 0 0.00098422 3.3 0.0009841399999999999 3.3 0.00098424 0 0.00098416 0 0.00098426 3.3 0.0009841799999999999 3.3 0.00098428 0 0.0009842 0 0.0009843 3.3 0.0009842199999999998 3.3 0.00098432 0 0.00098424 0 0.00098434 3.3 0.0009842599999999998 3.3 0.0009843599999999999 0 0.00098428 0 0.00098438 3.3 0.0009843 3.3 0.0009844 0 0.00098432 0 0.00098442 3.3 0.00098434 3.3 0.00098444 0 0.0009843599999999999 0 0.00098446 3.3 0.00098438 3.3 0.00098448 0 0.0009843999999999999 0 0.0009845 3.3 0.00098442 3.3 0.00098452 0 0.0009844399999999998 0 0.00098454 3.3 0.00098446 3.3 0.00098456 0 0.0009844799999999998 0 0.0009845799999999999 3.3 0.0009845 3.3 0.0009846 0 0.00098452 0 0.00098462 3.3 0.00098454 3.3 0.00098464 0 0.00098456 0 0.00098466 3.3 0.0009845799999999999 3.3 0.00098468 0 0.0009846 0 0.0009847 3.3 0.0009846199999999999 3.3 0.00098472 0 0.00098464 0 0.00098474 3.3 0.0009846599999999998 3.3 0.0009847599999999999 0 0.00098468 0 0.00098478 3.3 0.0009847 3.3 0.0009848 0 0.00098472 0 0.00098482 3.3 0.00098474 3.3 0.00098484 0 0.0009847599999999999 0 0.00098486 3.3 0.00098478 3.3 0.00098488 0 0.0009847999999999999 0 0.0009849 3.3 0.00098482 3.3 0.00098492 0 0.0009848399999999998 0 0.00098494 3.3 0.00098486 3.3 0.00098496 0 0.0009848799999999998 0 0.0009849799999999999 3.3 0.0009849 3.3 0.000985 0 0.00098492 0 0.00098502 3.3 0.00098494 3.3 0.00098504 0 0.00098496 0 0.00098506 3.3 0.0009849799999999999 3.3 0.00098508 0 0.000985 0 0.0009851 3.3 0.0009850199999999999 3.3 0.00098512 0 0.00098504 0 0.00098514 3.3 0.0009850599999999998 3.3 0.00098516 0 0.00098508 0 0.00098518 3.3 0.0009850999999999998 3.3 0.0009851999999999999 0 0.00098512 0 0.00098522 3.3 0.00098514 3.3 0.00098524 0 0.00098516 0 0.00098526 3.3 0.00098518 3.3 0.00098528 0 0.0009851999999999999 0 0.0009853 3.3 0.00098522 3.3 0.00098532 0 0.0009852399999999999 0 0.00098534 3.3 0.00098526 3.3 0.00098536 0 0.0009852799999999998 0 0.00098538 3.3 0.0009853 3.3 0.0009854 0 0.0009853199999999998 0 0.0009854199999999999 3.3 0.00098534 3.3 0.00098544 0 0.00098536 0 0.00098546 3.3 0.00098538 3.3 0.00098548 0 0.0009854 0 0.0009855 3.3 0.0009854199999999999 3.3 0.00098552 0 0.00098544 0 0.00098554 3.3 0.0009854599999999999 3.3 0.00098556 0 0.00098548 0 0.00098558 3.3 0.0009854999999999998 3.3 0.0009855999999999999 0 0.00098552 0 0.00098562 3.3 0.00098554 3.3 0.00098564 0 0.00098556 0 0.00098566 3.3 0.00098558 3.3 0.00098568 0 0.0009855999999999999 0 0.0009857 3.3 0.00098562 3.3 0.00098572 0 0.0009856399999999999 0 0.00098574 3.3 0.00098566 3.3 0.00098576 0 0.0009856799999999998 0 0.00098578 3.3 0.0009857 3.3 0.0009858 0 0.0009857199999999998 0 0.0009858199999999999 3.3 0.00098574 3.3 0.00098584 0 0.00098576 0 0.00098586 3.3 0.00098578 3.3 0.00098588 0 0.0009858 0 0.0009859 3.3 0.0009858199999999999 3.3 0.00098592 0 0.00098584 0 0.00098594 3.3 0.0009858599999999999 3.3 0.00098596 0 0.00098588 0 0.00098598 3.3 0.0009858999999999998 3.3 0.000986 0 0.00098592 0 0.00098602 3.3 0.0009859399999999998 3.3 0.0009860399999999999 0 0.00098596 0 0.00098606 3.3 0.00098598 3.3 0.00098608 0 0.000986 0 0.0009861 3.3 0.00098602 3.3 0.00098612 0 0.0009860399999999999 0 0.00098614 3.3 0.00098606 3.3 0.00098616 0 0.0009860799999999999 0 0.00098618 3.3 0.0009861 3.3 0.0009862 0 0.0009861199999999998 0 0.00098622 3.3 0.00098614 3.3 0.00098624 0 0.00098616 0 0.00098626 3.3 0.00098618 3.3 0.00098628 0 0.0009862 0 0.0009863 3.3 0.00098622 3.3 0.00098632 0 0.00098624 0 0.00098634 3.3 0.0009862599999999999 3.3 0.00098636 0 0.00098628 0 0.00098638 3.3 0.0009862999999999999 3.3 0.0009864 0 0.00098632 0 0.00098642 3.3 0.0009863399999999998 3.3 0.0009864399999999999 0 0.00098636 0 0.00098646 3.3 0.00098638 3.3 0.00098648 0 0.0009864 0 0.0009865 3.3 0.00098642 3.3 0.00098652 0 0.0009864399999999999 0 0.00098654 3.3 0.00098646 3.3 0.00098656 0 0.0009864799999999999 0 0.00098658 3.3 0.0009865 3.3 0.0009866 0 0.0009865199999999998 0 0.00098662 3.3 0.00098654 3.3 0.00098664 0 0.0009865599999999998 0 0.0009866599999999999 3.3 0.00098658 3.3 0.00098668 0 0.0009866 0 0.0009867 3.3 0.00098662 3.3 0.00098672 0 0.00098664 0 0.00098674 3.3 0.0009866599999999999 3.3 0.00098676 0 0.00098668 0 0.00098678 3.3 0.0009866999999999999 3.3 0.0009868 0 0.00098672 0 0.00098682 3.3 0.0009867399999999998 3.3 0.00098684 0 0.00098676 0 0.00098686 3.3 0.0009867799999999998 3.3 0.0009868799999999999 0 0.0009868 0 0.0009869 3.3 0.00098682 3.3 0.00098692 0 0.00098684 0 0.00098694 3.3 0.00098686 3.3 0.00098696 0 0.0009868799999999999 0 0.00098698 3.3 0.0009869 3.3 0.000987 0 0.0009869199999999999 0 0.00098702 3.3 0.00098694 3.3 0.00098704 0 0.0009869599999999998 0 0.0009870599999999999 3.3 0.00098698 3.3 0.00098708 0 0.000987 0 0.0009871 3.3 0.00098702 3.3 0.00098712 0 0.00098704 0 0.00098714 3.3 0.0009870599999999999 3.3 0.00098716 0 0.00098708 0 0.00098718 3.3 0.0009870999999999999 3.3 0.0009872 0 0.00098712 0 0.00098722 3.3 0.0009871399999999998 3.3 0.00098724 0 0.00098716 0 0.00098726 3.3 0.0009871799999999998 3.3 0.0009872799999999999 0 0.0009872 0 0.0009873 3.3 0.00098722 3.3 0.00098732 0 0.00098724 0 0.00098734 3.3 0.00098726 3.3 0.00098736 0 0.0009872799999999999 0 0.00098738 3.3 0.0009873 3.3 0.0009874 0 0.0009873199999999999 0 0.00098742 3.3 0.00098734 3.3 0.00098744 0 0.0009873599999999998 0 0.00098746 3.3 0.00098738 3.3 0.00098748 0 0.0009873999999999998 0 0.0009874999999999999 3.3 0.00098742 3.3 0.00098752 0 0.00098744 0 0.00098754 3.3 0.00098746 3.3 0.00098756 0 0.00098748 0 0.00098758 3.3 0.0009874999999999999 3.3 0.0009876 0 0.00098752 0 0.00098762 3.3 0.0009875399999999999 3.3 0.00098764 0 0.00098756 0 0.00098766 3.3 0.0009875799999999998 3.3 0.00098768 0 0.0009876 0 0.0009877 3.3 0.0009876199999999998 3.3 0.0009877199999999999 0 0.00098764 0 0.00098774 3.3 0.00098766 3.3 0.00098776 0 0.00098768 0 0.00098778 3.3 0.0009877 3.3 0.0009878 0 0.0009877199999999999 0 0.00098782 3.3 0.00098774 3.3 0.00098784 0 0.0009877599999999999 0 0.00098786 3.3 0.00098778 3.3 0.00098788 0 0.0009877999999999998 0 0.0009878999999999999 3.3 0.00098782 3.3 0.00098792 0 0.00098784 0 0.00098794 3.3 0.00098786 3.3 0.00098796 0 0.00098788 0 0.00098798 3.3 0.0009878999999999999 3.3 0.000988 0 0.00098792 0 0.00098802 3.3 0.0009879399999999999 3.3 0.00098804 0 0.00098796 0 0.00098806 3.3 0.0009879799999999998 3.3 0.00098808 0 0.000988 0 0.0009881 3.3 0.0009880199999999998 3.3 0.0009881199999999999 0 0.00098804 0 0.00098814 3.3 0.00098806 3.3 0.00098816 0 0.00098808 0 0.00098818 3.3 0.0009881 3.3 0.0009882 0 0.0009881199999999999 0 0.00098822 3.3 0.00098814 3.3 0.00098824 0 0.0009881599999999999 0 0.00098826 3.3 0.00098818 3.3 0.00098828 0 0.0009881999999999998 0 0.0009883 3.3 0.00098822 3.3 0.00098832 0 0.0009882399999999998 0 0.0009883399999999999 3.3 0.00098826 3.3 0.00098836 0 0.00098828 0 0.00098838 3.3 0.0009883 3.3 0.0009884 0 0.00098832 0 0.00098842 3.3 0.0009883399999999999 3.3 0.00098844 0 0.00098836 0 0.00098846 3.3 0.0009883799999999999 3.3 0.00098848 0 0.0009884 0 0.0009885 3.3 0.0009884199999999998 3.3 0.00098852 0 0.00098844 0 0.00098854 3.3 0.0009884599999999998 3.3 0.0009885599999999999 0 0.00098848 0 0.00098858 3.3 0.0009885 3.3 0.0009886 0 0.00098852 0 0.00098862 3.3 0.00098854 3.3 0.00098864 0 0.0009885599999999999 0 0.00098866 3.3 0.00098858 3.3 0.00098868 0 0.0009885999999999999 0 0.0009887 3.3 0.00098862 3.3 0.00098872 0 0.0009886399999999998 0 0.0009887399999999999 3.3 0.00098866 3.3 0.00098876 0 0.00098868 0 0.00098878 3.3 0.0009887 3.3 0.0009888 0 0.00098872 0 0.00098882 3.3 0.0009887399999999999 3.3 0.00098884 0 0.00098876 0 0.00098886 3.3 0.0009887799999999999 3.3 0.00098888 0 0.0009888 0 0.0009889 3.3 0.0009888199999999998 3.3 0.00098892 0 0.00098884 0 0.00098894 3.3 0.0009888599999999998 3.3 0.0009889599999999999 0 0.00098888 0 0.00098898 3.3 0.0009889 3.3 0.000989 0 0.00098892 0 0.00098902 3.3 0.00098894 3.3 0.00098904 0 0.0009889599999999999 0 0.00098906 3.3 0.00098898 3.3 0.00098908 0 0.0009889999999999999 0 0.0009891 3.3 0.00098902 3.3 0.00098912 0 0.0009890399999999998 0 0.00098914 3.3 0.00098906 3.3 0.00098916 0 0.0009890799999999998 0 0.0009891799999999999 3.3 0.0009891 3.3 0.0009892 0 0.00098912 0 0.00098922 3.3 0.00098914 3.3 0.00098924 0 0.00098916 0 0.00098926 3.3 0.0009891799999999999 3.3 0.00098928 0 0.0009892 0 0.0009893 3.3 0.0009892199999999999 3.3 0.00098932 0 0.00098924 0 0.00098934 3.3 0.0009892599999999998 3.3 0.00098936 0 0.00098928 0 0.00098938 3.3 0.0009893 3.3 0.0009894 0 0.00098932 0 0.00098942 3.3 0.00098934 3.3 0.00098944 0 0.00098936 0 0.00098946 3.3 0.00098938 3.3 0.00098948 0 0.0009893999999999999 0 0.0009895 3.3 0.00098942 3.3 0.00098952 0 0.0009894399999999999 0 0.00098954 3.3 0.00098946 3.3 0.00098956 0 0.0009894799999999998 0 0.0009895799999999999 3.3 0.0009895 3.3 0.0009896 0 0.00098952 0 0.00098962 3.3 0.00098954 3.3 0.00098964 0 0.00098956 0 0.00098966 3.3 0.0009895799999999999 3.3 0.00098968 0 0.0009896 0 0.0009897 3.3 0.0009896199999999999 3.3 0.00098972 0 0.00098964 0 0.00098974 3.3 0.0009896599999999998 3.3 0.00098976 0 0.00098968 0 0.00098978 3.3 0.0009896999999999998 3.3 0.0009897999999999999 0 0.00098972 0 0.00098982 3.3 0.00098974 3.3 0.00098984 0 0.00098976 0 0.00098986 3.3 0.00098978 3.3 0.00098988 0 0.0009897999999999999 0 0.0009899 3.3 0.00098982 3.3 0.00098992 0 0.0009898399999999999 0 0.00098994 3.3 0.00098986 3.3 0.00098996 0 0.0009898799999999998 0 0.00098998 3.3 0.0009899 3.3 0.00099 0 0.0009899199999999998 0 0.0009900199999999999 3.3 0.00098994 3.3 0.00099004 0 0.00098996 0 0.00099006 3.3 0.00098998 3.3 0.00099008 0 0.00099 0 0.0009901 3.3 0.0009900199999999999 3.3 0.00099012 0 0.00099004 0 0.00099014 3.3 0.0009900599999999999 3.3 0.00099016 0 0.00099008 0 0.00099018 3.3 0.0009900999999999998 3.3 0.0009901999999999999 0 0.00099012 0 0.00099022 3.3 0.00099014 3.3 0.00099024 0 0.00099016 0 0.00099026 3.3 0.00099018 3.3 0.00099028 0 0.0009901999999999999 0 0.0009903 3.3 0.00099022 3.3 0.00099032 0 0.0009902399999999999 0 0.00099034 3.3 0.00099026 3.3 0.00099036 0 0.0009902799999999998 0 0.00099038 3.3 0.0009903 3.3 0.0009904 0 0.0009903199999999998 0 0.0009904199999999999 3.3 0.00099034 3.3 0.00099044 0 0.00099036 0 0.00099046 3.3 0.00099038 3.3 0.00099048 0 0.0009904 0 0.0009905 3.3 0.0009904199999999999 3.3 0.00099052 0 0.00099044 0 0.00099054 3.3 0.0009904599999999999 3.3 0.00099056 0 0.00099048 0 0.00099058 3.3 0.0009904999999999998 3.3 0.0009906 0 0.00099052 0 0.00099062 3.3 0.0009905399999999998 3.3 0.0009906399999999999 0 0.00099056 0 0.00099066 3.3 0.00099058 3.3 0.00099068 0 0.0009906 0 0.0009907 3.3 0.00099062 3.3 0.00099072 0 0.0009906399999999999 0 0.00099074 3.3 0.00099066 3.3 0.00099076 0 0.0009906799999999999 0 0.00099078 3.3 0.0009907 3.3 0.0009908 0 0.0009907199999999998 0 0.00099082 3.3 0.00099074 3.3 0.00099084 0 0.0009907599999999998 0 0.0009908599999999999 3.3 0.00099078 3.3 0.00099088 0 0.0009908 0 0.0009909 3.3 0.00099082 3.3 0.00099092 0 0.00099084 0 0.00099094 3.3 0.0009908599999999999 3.3 0.00099096 0 0.00099088 0 0.00099098 3.3 0.0009908999999999999 3.3 0.000991 0 0.00099092 0 0.00099102 3.3 0.0009909399999999998 3.3 0.0009910399999999999 0 0.00099096 0 0.00099106 3.3 0.00099098 3.3 0.00099108 0 0.000991 0 0.0009911 3.3 0.00099102 3.3 0.00099112 0 0.0009910399999999999 0 0.00099114 3.3 0.00099106 3.3 0.00099116 0 0.0009910799999999999 0 0.00099118 3.3 0.0009911 3.3 0.0009912 0 0.0009911199999999998 0 0.00099122 3.3 0.00099114 3.3 0.00099124 0 0.0009911599999999998 0 0.0009912599999999999 3.3 0.00099118 3.3 0.00099128 0 0.0009912 0 0.0009913 3.3 0.00099122 3.3 0.00099132 0 0.00099124 0 0.00099134 3.3 0.0009912599999999999 3.3 0.00099136 0 0.00099128 0 0.00099138 3.3 0.0009912999999999999 3.3 0.0009914 0 0.00099132 0 0.00099142 3.3 0.0009913399999999998 3.3 0.00099144 0 0.00099136 0 0.00099146 3.3 0.0009913799999999998 3.3 0.0009914799999999999 0 0.0009914 0 0.0009915 3.3 0.00099142 3.3 0.00099152 0 0.00099144 0 0.00099154 3.3 0.00099146 3.3 0.00099156 0 0.0009914799999999999 0 0.00099158 3.3 0.0009915 3.3 0.0009916 0 0.0009915199999999999 0 0.00099162 3.3 0.00099154 3.3 0.00099164 0 0.0009915599999999998 0 0.00099166 3.3 0.00099158 3.3 0.00099168 0 0.0009915999999999998 0 0.0009916999999999999 3.3 0.00099162 3.3 0.00099172 0 0.00099164 0 0.00099174 3.3 0.00099166 3.3 0.00099176 0 0.00099168 0 0.00099178 3.3 0.0009916999999999999 3.3 0.0009918 0 0.00099172 0 0.00099182 3.3 0.0009917399999999999 3.3 0.00099184 0 0.00099176 0 0.00099186 3.3 0.0009917799999999998 3.3 0.0009918799999999999 0 0.0009918 0 0.0009919 3.3 0.00099182 3.3 0.00099192 0 0.00099184 0 0.00099194 3.3 0.00099186 3.3 0.00099196 0 0.0009918799999999999 0 0.00099198 3.3 0.0009919 3.3 0.000992 0 0.0009919199999999999 0 0.00099202 3.3 0.00099194 3.3 0.00099204 0 0.0009919599999999998 0 0.00099206 3.3 0.00099198 3.3 0.00099208 0 0.0009919999999999998 0 0.0009920999999999999 3.3 0.00099202 3.3 0.00099212 0 0.00099204 0 0.00099214 3.3 0.00099206 3.3 0.00099216 0 0.00099208 0 0.00099218 3.3 0.0009920999999999999 3.3 0.0009922 0 0.00099212 0 0.00099222 3.3 0.0009921399999999999 3.3 0.00099224 0 0.00099216 0 0.00099226 3.3 0.0009921799999999998 3.3 0.00099228 0 0.0009922 0 0.0009923 3.3 0.0009922199999999998 3.3 0.0009923199999999999 0 0.00099224 0 0.00099234 3.3 0.00099226 3.3 0.00099236 0 0.00099228 0 0.00099238 3.3 0.0009923 3.3 0.0009924 0 0.0009923199999999999 0 0.00099242 3.3 0.00099234 3.3 0.00099244 0 0.0009923599999999999 0 0.00099246 3.3 0.00099238 3.3 0.00099248 0 0.0009923999999999998 0 0.0009925 3.3 0.00099242 3.3 0.00099252 0 0.0009924399999999998 0 0.0009925399999999999 3.3 0.00099246 3.3 0.00099256 0 0.00099248 0 0.00099258 3.3 0.0009925 3.3 0.0009926 0 0.00099252 0 0.00099262 3.3 0.0009925399999999999 3.3 0.00099264 0 0.00099256 0 0.00099266 3.3 0.0009925799999999999 3.3 0.00099268 0 0.0009926 0 0.0009927 3.3 0.0009926199999999998 3.3 0.0009927199999999999 0 0.00099264 0 0.00099274 3.3 0.00099266 3.3 0.00099276 0 0.00099268 0 0.00099278 3.3 0.0009927 3.3 0.0009928 0 0.0009927199999999999 0 0.00099282 3.3 0.00099274 3.3 0.00099284 0 0.0009927599999999999 0 0.00099286 3.3 0.00099278 3.3 0.00099288 0 0.0009927999999999998 0 0.0009929 3.3 0.00099282 3.3 0.00099292 0 0.0009928399999999998 0 0.0009929399999999999 3.3 0.00099286 3.3 0.00099296 0 0.00099288 0 0.00099298 3.3 0.0009929 3.3 0.000993 0 0.00099292 0 0.00099302 3.3 0.0009929399999999999 3.3 0.00099304 0 0.00099296 0 0.00099306 3.3 0.0009929799999999999 3.3 0.00099308 0 0.000993 0 0.0009931 3.3 0.0009930199999999998 3.3 0.00099312 0 0.00099304 0 0.00099314 3.3 0.0009930599999999998 3.3 0.0009931599999999999 0 0.00099308 0 0.00099318 3.3 0.0009931 3.3 0.0009932 0 0.00099312 0 0.00099322 3.3 0.00099314 3.3 0.00099324 0 0.0009931599999999999 0 0.00099326 3.3 0.00099318 3.3 0.00099328 0 0.0009931999999999999 0 0.0009933 3.3 0.00099322 3.3 0.00099332 0 0.0009932399999999998 0 0.0009933399999999999 3.3 0.00099326 3.3 0.00099336 0 0.00099328 0 0.00099338 3.3 0.0009933 3.3 0.0009934 0 0.00099332 0 0.00099342 3.3 0.0009933399999999999 3.3 0.00099344 0 0.00099336 0 0.00099346 3.3 0.0009933799999999999 3.3 0.00099348 0 0.0009934 0 0.0009935 3.3 0.0009934199999999999 3.3 0.00099352 0 0.00099344 0 0.00099354 3.3 0.0009934599999999998 3.3 0.0009935599999999999 0 0.00099348 0 0.00099358 3.3 0.0009935 3.3 0.0009936 0 0.00099352 0 0.00099362 3.3 0.00099354 3.3 0.00099364 0 0.0009935599999999999 0 0.00099366 3.3 0.00099358 3.3 0.00099368 0 0.0009935999999999999 0 0.0009937 3.3 0.00099362 3.3 0.00099372 0 0.0009936399999999998 0 0.00099374 3.3 0.00099366 3.3 0.00099376 0 0.0009936799999999998 0 0.0009937799999999999 3.3 0.0009937 3.3 0.0009938 0 0.00099372 0 0.00099382 3.3 0.00099374 3.3 0.00099384 0 0.00099376 0 0.00099386 3.3 0.0009937799999999999 3.3 0.00099388 0 0.0009938 0 0.0009939 3.3 0.0009938199999999999 3.3 0.00099392 0 0.00099384 0 0.00099394 3.3 0.0009938599999999998 3.3 0.00099396 0 0.00099388 0 0.00099398 3.3 0.0009938999999999998 3.3 0.0009939999999999999 0 0.00099392 0 0.00099402 3.3 0.00099394 3.3 0.00099404 0 0.00099396 0 0.00099406 3.3 0.00099398 3.3 0.00099408 0 0.0009939999999999999 0 0.0009941 3.3 0.00099402 3.3 0.00099412 0 0.0009940399999999999 0 0.00099414 3.3 0.00099406 3.3 0.00099416 0 0.0009940799999999998 0 0.0009941799999999999 3.3 0.0009941 3.3 0.0009942 0 0.00099412 0 0.00099422 3.3 0.00099414 3.3 0.00099424 0 0.00099416 0 0.00099426 3.3 0.0009941799999999999 3.3 0.00099428 0 0.0009942 0 0.0009943 3.3 0.0009942199999999999 3.3 0.00099432 0 0.00099424 0 0.00099434 3.3 0.0009942599999999998 3.3 0.00099436 0 0.00099428 0 0.00099438 3.3 0.0009942999999999998 3.3 0.0009943999999999999 0 0.00099432 0 0.00099442 3.3 0.00099434 3.3 0.00099444 0 0.00099436 0 0.00099446 3.3 0.00099438 3.3 0.00099448 0 0.0009943999999999999 0 0.0009945 3.3 0.00099442 3.3 0.00099452 0 0.0009944399999999999 0 0.00099454 3.3 0.00099446 3.3 0.00099456 0 0.0009944799999999998 0 0.00099458 3.3 0.0009945 3.3 0.0009946 0 0.0009945199999999998 0 0.0009946199999999999 3.3 0.00099454 3.3 0.00099464 0 0.00099456 0 0.00099466 3.3 0.00099458 3.3 0.00099468 0 0.0009946 0 0.0009947 3.3 0.0009946199999999999 3.3 0.00099472 0 0.00099464 0 0.00099474 3.3 0.0009946599999999999 3.3 0.00099476 0 0.00099468 0 0.00099478 3.3 0.0009946999999999998 3.3 0.0009948 0 0.00099472 0 0.00099482 3.3 0.0009947399999999998 3.3 0.0009948399999999999 0 0.00099476 0 0.00099486 3.3 0.00099478 3.3 0.00099488 0 0.0009948 0 0.0009949 3.3 0.00099482 3.3 0.00099492 0 0.0009948399999999999 0 0.00099494 3.3 0.00099486 3.3 0.00099496 0 0.0009948799999999999 0 0.00099498 3.3 0.0009949 3.3 0.000995 0 0.0009949199999999998 0 0.0009950199999999999 3.3 0.00099494 3.3 0.00099504 0 0.00099496 0 0.00099506 3.3 0.00099498 3.3 0.00099508 0 0.000995 0 0.0009951 3.3 0.0009950199999999999 3.3 0.00099512 0 0.00099504 0 0.00099514 3.3 0.0009950599999999999 3.3 0.00099516 0 0.00099508 0 0.00099518 3.3 0.0009950999999999998 3.3 0.0009952 0 0.00099512 0 0.00099522 3.3 0.0009951399999999998 3.3 0.0009952399999999999 0 0.00099516 0 0.00099526 3.3 0.00099518 3.3 0.00099528 0 0.0009952 0 0.0009953 3.3 0.00099522 3.3 0.00099532 0 0.0009952399999999999 0 0.00099534 3.3 0.00099526 3.3 0.00099536 0 0.0009952799999999999 0 0.00099538 3.3 0.0009953 3.3 0.0009954 0 0.0009953199999999998 0 0.00099542 3.3 0.00099534 3.3 0.00099544 0 0.0009953599999999998 0 0.0009954599999999999 3.3 0.00099538 3.3 0.00099548 0 0.0009954 0 0.0009955 3.3 0.00099542 3.3 0.00099552 0 0.00099544 0 0.00099554 3.3 0.0009954599999999999 3.3 0.00099556 0 0.00099548 0 0.00099558 3.3 0.0009954999999999999 3.3 0.0009956 0 0.00099552 0 0.00099562 3.3 0.0009955399999999998 3.3 0.00099564 0 0.00099556 0 0.00099566 3.3 0.0009955799999999998 3.3 0.0009956799999999999 0 0.0009956 0 0.0009957 3.3 0.00099562 3.3 0.00099572 0 0.00099564 0 0.00099574 3.3 0.00099566 3.3 0.00099576 0 0.0009956799999999999 0 0.00099578 3.3 0.0009957 3.3 0.0009958 0 0.0009957199999999999 0 0.00099582 3.3 0.00099574 3.3 0.00099584 0 0.0009957599999999998 0 0.0009958599999999999 3.3 0.00099578 3.3 0.00099588 0 0.0009958 0 0.0009959 3.3 0.00099582 3.3 0.00099592 0 0.00099584 0 0.00099594 3.3 0.0009958599999999999 3.3 0.00099596 0 0.00099588 0 0.00099598 3.3 0.0009958999999999999 3.3 0.000996 0 0.00099592 0 0.00099602 3.3 0.0009959399999999998 3.3 0.00099604 0 0.00099596 0 0.00099606 3.3 0.0009959799999999998 3.3 0.0009960799999999999 0 0.000996 0 0.0009961 3.3 0.00099602 3.3 0.00099612 0 0.00099604 0 0.00099614 3.3 0.00099606 3.3 0.00099616 0 0.0009960799999999999 0 0.00099618 3.3 0.0009961 3.3 0.0009962 0 0.0009961199999999999 0 0.00099622 3.3 0.00099614 3.3 0.00099624 0 0.0009961599999999998 0 0.00099626 3.3 0.00099618 3.3 0.00099628 0 0.0009961999999999998 0 0.0009962999999999999 3.3 0.00099622 3.3 0.00099632 0 0.00099624 0 0.00099634 3.3 0.00099626 3.3 0.00099636 0 0.00099628 0 0.00099638 3.3 0.0009962999999999999 3.3 0.0009964 0 0.00099632 0 0.00099642 3.3 0.0009963399999999999 3.3 0.00099644 0 0.00099636 0 0.00099646 3.3 0.0009963799999999998 3.3 0.00099648 0 0.0009964 0 0.0009965 3.3 0.00099642 3.3 0.00099652 0 0.00099644 0 0.00099654 3.3 0.00099646 3.3 0.00099656 0 0.00099648 0 0.00099658 3.3 0.0009965 3.3 0.0009966 0 0.0009965199999999999 0 0.00099662 3.3 0.00099654 3.3 0.00099664 0 0.0009965599999999999 0 0.00099666 3.3 0.00099658 3.3 0.00099668 0 0.0009965999999999998 0 0.0009966999999999999 3.3 0.00099662 3.3 0.00099672 0 0.00099664 0 0.00099674 3.3 0.00099666 3.3 0.00099676 0 0.00099668 0 0.00099678 3.3 0.0009966999999999999 3.3 0.0009968 0 0.00099672 0 0.00099682 3.3 0.0009967399999999999 3.3 0.00099684 0 0.00099676 0 0.00099686 3.3 0.0009967799999999998 3.3 0.00099688 0 0.0009968 0 0.0009969 3.3 0.0009968199999999998 3.3 0.0009969199999999999 0 0.00099684 0 0.00099694 3.3 0.00099686 3.3 0.00099696 0 0.00099688 0 0.00099698 3.3 0.0009969 3.3 0.000997 0 0.0009969199999999999 0 0.00099702 3.3 0.00099694 3.3 0.00099704 0 0.0009969599999999999 0 0.00099706 3.3 0.00099698 3.3 0.00099708 0 0.0009969999999999998 0 0.0009971 3.3 0.00099702 3.3 0.00099712 0 0.0009970399999999998 0 0.0009971399999999999 3.3 0.00099706 3.3 0.00099716 0 0.00099708 0 0.00099718 3.3 0.0009971 3.3 0.0009972 0 0.00099712 0 0.00099722 3.3 0.0009971399999999999 3.3 0.00099724 0 0.00099716 0 0.00099726 3.3 0.0009971799999999999 3.3 0.00099728 0 0.0009972 0 0.0009973 3.3 0.0009972199999999998 3.3 0.0009973199999999999 0 0.00099724 0 0.00099734 3.3 0.00099726 3.3 0.00099736 0 0.00099728 0 0.00099738 3.3 0.0009973 3.3 0.0009974 0 0.0009973199999999999 0 0.00099742 3.3 0.00099734 3.3 0.00099744 0 0.0009973599999999999 0 0.00099746 3.3 0.00099738 3.3 0.00099748 0 0.0009973999999999998 0 0.0009975 3.3 0.00099742 3.3 0.00099752 0 0.0009974399999999998 0 0.0009975399999999999 3.3 0.00099746 3.3 0.00099756 0 0.00099748 0 0.00099758 3.3 0.0009975 3.3 0.0009976 0 0.00099752 0 0.00099762 3.3 0.0009975399999999999 3.3 0.00099764 0 0.00099756 0 0.00099766 3.3 0.0009975799999999999 3.3 0.00099768 0 0.0009976 0 0.0009977 3.3 0.0009976199999999998 3.3 0.00099772 0 0.00099764 0 0.00099774 3.3 0.0009976599999999998 3.3 0.0009977599999999999 0 0.00099768 0 0.00099778 3.3 0.0009977 3.3 0.0009978 0 0.00099772 0 0.00099782 3.3 0.00099774 3.3 0.00099784 0 0.0009977599999999999 0 0.00099786 3.3 0.00099778 3.3 0.00099788 0 0.0009977999999999999 0 0.0009979 3.3 0.00099782 3.3 0.00099792 0 0.0009978399999999998 0 0.00099794 3.3 0.00099786 3.3 0.00099796 0 0.0009978799999999998 0 0.0009979799999999999 3.3 0.0009979 3.3 0.000998 0 0.00099792 0 0.00099802 3.3 0.00099794 3.3 0.00099804 0 0.00099796 0 0.00099806 3.3 0.0009979799999999999 3.3 0.00099808 0 0.000998 0 0.0009981 3.3 0.0009980199999999999 3.3 0.00099812 0 0.00099804 0 0.00099814 3.3 0.0009980599999999998 3.3 0.0009981599999999999 0 0.00099808 0 0.00099818 3.3 0.0009981 3.3 0.0009982 0 0.00099812 0 0.00099822 3.3 0.00099814 3.3 0.00099824 0 0.0009981599999999999 0 0.00099826 3.3 0.00099818 3.3 0.00099828 0 0.0009981999999999999 0 0.0009983 3.3 0.00099822 3.3 0.00099832 0 0.0009982399999999998 0 0.00099834 3.3 0.00099826 3.3 0.00099836 0 0.0009982799999999998 0 0.0009983799999999999 3.3 0.0009983 3.3 0.0009984 0 0.00099832 0 0.00099842 3.3 0.00099834 3.3 0.00099844 0 0.00099836 0 0.00099846 3.3 0.0009983799999999999 3.3 0.00099848 0 0.0009984 0 0.0009985 3.3 0.0009984199999999999 3.3 0.00099852 0 0.00099844 0 0.00099854 3.3 0.0009984599999999998 3.3 0.00099856 0 0.00099848 0 0.00099858 3.3 0.0009984999999999998 3.3 0.0009985999999999999 0 0.00099852 0 0.00099862 3.3 0.00099854 3.3 0.00099864 0 0.00099856 0 0.00099866 3.3 0.00099858 3.3 0.00099868 0 0.0009985999999999999 0 0.0009987 3.3 0.00099862 3.3 0.00099872 0 0.0009986399999999999 0 0.00099874 3.3 0.00099866 3.3 0.00099876 0 0.0009986799999999998 0 0.00099878 3.3 0.0009987 3.3 0.0009988 0 0.0009987199999999998 0 0.0009988199999999999 3.3 0.00099874 3.3 0.00099884 0 0.00099876 0 0.00099886 3.3 0.00099878 3.3 0.00099888 0 0.0009988 0 0.0009989 3.3 0.0009988199999999999 3.3 0.00099892 0 0.00099884 0 0.00099894 3.3 0.0009988599999999999 3.3 0.00099896 0 0.00099888 0 0.00099898 3.3 0.0009988999999999998 3.3 0.0009989999999999999 0 0.00099892 0 0.00099902 3.3 0.00099894 3.3 0.00099904 0 0.00099896 0 0.00099906 3.3 0.00099898 3.3 0.00099908 0 0.0009989999999999999 0 0.0009991 3.3 0.00099902 3.3 0.00099912 0 0.0009990399999999999 0 0.00099914 3.3 0.00099906 3.3 0.00099916 0 0.0009990799999999998 0 0.00099918 3.3 0.0009991 3.3 0.0009992 0 0.0009991199999999998 0 0.0009992199999999999 3.3 0.00099914 3.3 0.00099924 0 0.00099916 0 0.00099926 3.3 0.00099918 3.3 0.00099928 0 0.0009992 0 0.0009993 3.3 0.0009992199999999999 3.3 0.00099932 0 0.00099924 0 0.00099934 3.3 0.0009992599999999999 3.3 0.00099936 0 0.00099928 0 0.00099938 3.3 0.0009992999999999998 3.3 0.0009994 0 0.00099932 0 0.00099942 3.3 0.0009993399999999998 3.3 0.0009994399999999999 0 0.00099936 0 0.00099946 3.3 0.00099938 3.3 0.00099948 0 0.0009994 0 0.0009995 3.3 0.00099942 3.3 0.00099952 0 0.0009994399999999999 0 0.00099954 3.3 0.00099946 3.3 0.00099956 0 0.0009994799999999999 0 0.00099958 3.3 0.0009995 3.3 0.0009996 0 0.0009995199999999998 0 0.00099962 3.3 0.00099954 3.3 0.00099964 0 0.0009995599999999998 0 0.0009996599999999999 3.3 0.00099958 3.3 0.00099968 0 0.0009996 0 0.0009997 3.3 0.00099962 3.3 0.00099972 0 0.00099964 0 0.00099974 3.3 0.0009996599999999999 3.3 0.00099976 0 0.00099968 0 0.00099978 3.3 0.0009996999999999999 3.3 0.0009998 0 0.00099972 0 0.00099982 3.3 0.0009997399999999998 3.3 0.0009998399999999999 0 0.00099976 0 0.00099986 3.3 0.00099978 3.3 0.00099988 0 0.0009998 0 0.0009999 3.3 0.00099982 3.3 0.00099992 0 0.0009998399999999999 0 0.00099994 3.3 0.00099986 3.3 0.00099996 0 0.0009998799999999999 0 0.00099998 3.3 0.0009999 3.3 0.001 0 0.0009999199999999998 0 0.00100002 3.3 0.00099994 3.3 0.00100004 0 0.0009999599999999998 0 0.0010000599999999999 3.3 0.00099998 3.3 0.00100008 0 0.001 0 0.0010001 3.3 0.00100002 3.3 0.00100012 0 0.00100004 0 0.00100014 3.3 0.0010000599999999999 3.3 0.00100016 0 0.00100008 0 0.00100018 3.3 0.0010000999999999999 3.3 0.0010002 0 0.00100012 0 0.00100022 3.3 0.0010001399999999998 3.3 0.00100024 0 0.00100016 0 0.00100026 3.3 0.0010001799999999998 3.3 0.0010002799999999999 0 0.0010002 0 0.0010003 3.3 0.00100022 3.3 0.00100032 0 0.00100024 0 0.00100034 3.3 0.00100026 3.3 0.00100036 0 0.0010002799999999999 0 0.00100038 3.3 0.0010003 3.3 0.0010004 0 0.0010003199999999999 0 0.00100042 3.3 0.00100034 3.3 0.00100044 0 0.0010003599999999998 0 0.0010004599999999999 3.3 0.00100038 3.3 0.00100048 0 0.0010004 0 0.0010005 3.3 0.00100042 3.3 0.00100052 0 0.00100044 0 0.00100054 3.3 0.0010004599999999999 3.3 0.00100056 0 0.00100048 0 0.00100058 3.3 0.0010004999999999999 3.3 0.0010006 0 0.00100052 0 0.00100062 3.3 0.0010005399999999998 3.3 0.00100064 0 0.00100056 0 0.00100066 3.3 0.0010005799999999998 3.3 0.0010006799999999999 0 0.0010006 0 0.0010007 3.3 0.00100062 3.3 0.00100072 0 0.00100064 0 0.00100074 3.3 0.00100066 3.3 0.00100076 0 0.0010006799999999999 0 0.00100078 3.3 0.0010007 3.3 0.0010008 0 0.0010007199999999999 0 0.00100082 3.3 0.00100074 3.3 0.00100084 0 0.0010007599999999998 0 0.00100086 3.3 0.00100078 3.3 0.00100088 0 0.0010007999999999998 0 0.0010008999999999999 3.3 0.00100082 3.3 0.00100092 0 0.00100084 0 0.00100094 3.3 0.00100086 3.3 0.00100096 0 0.00100088 0 0.00100098 3.3 0.0010008999999999999 3.3 0.001001 0 0.00100092 0 0.00100102 3.3 0.0010009399999999999 3.3 0.00100104 0 0.00100096 0 0.00100106 3.3 0.0010009799999999998 3.3 0.00100108 0 0.001001 0 0.0010011 3.3 0.0010010199999999998 3.3 0.0010011199999999999 0 0.00100104 0 0.00100114 3.3 0.00100106 3.3 0.00100116 0 0.00100108 0 0.00100118 3.3 0.0010011 3.3 0.0010012 0 0.0010011199999999999 0 0.00100122 3.3 0.00100114 3.3 0.00100124 0 0.0010011599999999999 0 0.00100126 3.3 0.00100118 3.3 0.00100128 0 0.0010011999999999998 0 0.0010012999999999999 3.3 0.00100122 3.3 0.00100132 0 0.00100124 0 0.00100134 3.3 0.00100126 3.3 0.00100136 0 0.00100128 0 0.00100138 3.3 0.0010012999999999999 3.3 0.0010014 0 0.00100132 0 0.00100142 3.3 0.0010013399999999999 3.3 0.00100144 0 0.00100136 0 0.00100146 3.3 0.0010013799999999998 3.3 0.00100148 0 0.0010014 0 0.0010015 3.3 0.0010014199999999998 3.3 0.0010015199999999999 0 0.00100144 0 0.00100154 3.3 0.00100146 3.3 0.00100156 0 0.00100148 0 0.00100158 3.3 0.0010015 3.3 0.0010016 0 0.0010015199999999999 0 0.00100162 3.3 0.00100154 3.3 0.00100164 0 0.0010015599999999999 0 0.00100166 3.3 0.00100158 3.3 0.00100168 0 0.0010015999999999998 0 0.0010017 3.3 0.00100162 3.3 0.00100172 0 0.0010016399999999998 0 0.0010017399999999999 3.3 0.00100166 3.3 0.00100176 0 0.00100168 0 0.00100178 3.3 0.0010017 3.3 0.0010018 0 0.00100172 0 0.00100182 3.3 0.0010017399999999999 3.3 0.00100184 0 0.00100176 0 0.00100186 3.3 0.0010017799999999999 3.3 0.00100188 0 0.0010018 0 0.0010019 3.3 0.0010018199999999998 3.3 0.00100192 0 0.00100184 0 0.00100194 3.3 0.0010018599999999998 3.3 0.0010019599999999999 0 0.00100188 0 0.00100198 3.3 0.0010019 3.3 0.001002 0 0.00100192 0 0.00100202 3.3 0.00100194 3.3 0.00100204 0 0.0010019599999999999 0 0.00100206 3.3 0.00100198 3.3 0.00100208 0 0.0010019999999999999 0 0.0010021 3.3 0.00100202 3.3 0.00100212 0 0.0010020399999999998 0 0.0010021399999999999 3.3 0.00100206 3.3 0.00100216 0 0.00100208 0 0.00100218 3.3 0.0010021 3.3 0.0010022 0 0.00100212 0 0.00100222 3.3 0.0010021399999999999 3.3 0.00100224 0 0.00100216 0 0.00100226 3.3 0.0010021799999999999 3.3 0.00100228 0 0.0010022 0 0.0010023 3.3 0.0010022199999999998 3.3 0.00100232 0 0.00100224 0 0.00100234 3.3 0.0010022599999999998 3.3 0.0010023599999999999 0 0.00100228 0 0.00100238 3.3 0.0010023 3.3 0.0010024 0 0.00100232 0 0.00100242 3.3 0.00100234 3.3 0.00100244 0 0.0010023599999999999 0 0.00100246 3.3 0.00100238 3.3 0.00100248 0 0.0010023999999999999 0 0.0010025 3.3 0.00100242 3.3 0.00100252 0 0.0010024399999999998 0 0.00100254 3.3 0.00100246 3.3 0.00100256 0 0.0010024799999999998 0 0.0010025799999999999 3.3 0.0010025 3.3 0.0010026 0 0.00100252 0 0.00100262 3.3 0.00100254 3.3 0.00100264 0 0.00100256 0 0.00100266 3.3 0.0010025799999999999 3.3 0.00100268 0 0.0010026 0 0.0010027 3.3 0.0010026199999999999 3.3 0.00100272 0 0.00100264 0 0.00100274 3.3 0.0010026599999999998 3.3 0.00100276 0 0.00100268 0 0.00100278 3.3 0.0010026999999999998 3.3 0.0010027999999999999 0 0.00100272 0 0.00100282 3.3 0.00100274 3.3 0.00100284 0 0.00100276 0 0.00100286 3.3 0.00100278 3.3 0.00100288 0 0.0010027999999999999 0 0.0010029 3.3 0.00100282 3.3 0.00100292 0 0.0010028399999999999 0 0.00100294 3.3 0.00100286 3.3 0.00100296 0 0.0010028799999999998 0 0.0010029799999999999 3.3 0.0010029 3.3 0.001003 0 0.00100292 0 0.00100302 3.3 0.00100294 3.3 0.00100304 0 0.00100296 0 0.00100306 3.3 0.0010029799999999999 3.3 0.00100308 0 0.001003 0 0.0010031 3.3 0.0010030199999999999 3.3 0.00100312 0 0.00100304 0 0.00100314 3.3 0.0010030599999999998 3.3 0.00100316 0 0.00100308 0 0.00100318 3.3 0.0010030999999999998 3.3 0.0010031999999999999 0 0.00100312 0 0.00100322 3.3 0.00100314 3.3 0.00100324 0 0.00100316 0 0.00100326 3.3 0.00100318 3.3 0.00100328 0 0.0010031999999999999 0 0.0010033 3.3 0.00100322 3.3 0.00100332 0 0.0010032399999999999 0 0.00100334 3.3 0.00100326 3.3 0.00100336 0 0.0010032799999999998 0 0.00100338 3.3 0.0010033 3.3 0.0010034 0 0.0010033199999999998 0 0.0010034199999999999 3.3 0.00100334 3.3 0.00100344 0 0.00100336 0 0.00100346 3.3 0.00100338 3.3 0.00100348 0 0.0010034 0 0.0010035 3.3 0.0010034199999999999 3.3 0.00100352 0 0.00100344 0 0.00100354 3.3 0.0010034599999999999 3.3 0.00100356 0 0.00100348 0 0.00100358 3.3 0.0010034999999999998 3.3 0.0010035999999999999 0 0.00100352 0 0.00100362 3.3 0.00100354 3.3 0.00100364 0 0.00100356 0 0.00100366 3.3 0.00100358 3.3 0.00100368 0 0.0010035999999999999 0 0.0010037 3.3 0.00100362 3.3 0.00100372 0 0.0010036399999999999 0 0.00100374 3.3 0.00100366 3.3 0.00100376 0 0.0010036799999999999 0 0.00100378 3.3 0.0010037 3.3 0.0010038 0 0.0010037199999999998 0 0.0010038199999999999 3.3 0.00100374 3.3 0.00100384 0 0.00100376 0 0.00100386 3.3 0.00100378 3.3 0.00100388 0 0.0010038 0 0.0010039 3.3 0.0010038199999999999 3.3 0.00100392 0 0.00100384 0 0.00100394 3.3 0.0010038599999999999 3.3 0.00100396 0 0.00100388 0 0.00100398 3.3 0.0010038999999999998 3.3 0.001004 0 0.00100392 0 0.00100402 3.3 0.0010039399999999998 3.3 0.0010040399999999999 0 0.00100396 0 0.00100406 3.3 0.00100398 3.3 0.00100408 0 0.001004 0 0.0010041 3.3 0.00100402 3.3 0.00100412 0 0.0010040399999999999 0 0.00100414 3.3 0.00100406 3.3 0.00100416 0 0.0010040799999999999 0 0.00100418 3.3 0.0010041 3.3 0.0010042 0 0.0010041199999999998 0 0.00100422 3.3 0.00100414 3.3 0.00100424 0 0.0010041599999999998 0 0.0010042599999999999 3.3 0.00100418 3.3 0.00100428 0 0.0010042 0 0.0010043 3.3 0.00100422 3.3 0.00100432 0 0.00100424 0 0.00100434 3.3 0.0010042599999999999 3.3 0.00100436 0 0.00100428 0 0.00100438 3.3 0.0010042999999999999 3.3 0.0010044 0 0.00100432 0 0.00100442 3.3 0.0010043399999999998 3.3 0.0010044399999999999 0 0.00100436 0 0.00100446 3.3 0.00100438 3.3 0.00100448 0 0.0010044 0 0.0010045 3.3 0.00100442 3.3 0.00100452 0 0.0010044399999999999 0 0.00100454 3.3 0.00100446 3.3 0.00100456 0 0.0010044799999999999 0 0.00100458 3.3 0.0010045 3.3 0.0010046 0 0.0010045199999999998 0 0.00100462 3.3 0.00100454 3.3 0.00100464 0 0.0010045599999999998 0 0.0010046599999999999 3.3 0.00100458 3.3 0.00100468 0 0.0010046 0 0.0010047 3.3 0.00100462 3.3 0.00100472 0 0.00100464 0 0.00100474 3.3 0.0010046599999999999 3.3 0.00100476 0 0.00100468 0 0.00100478 3.3 0.0010046999999999999 3.3 0.0010048 0 0.00100472 0 0.00100482 3.3 0.0010047399999999998 3.3 0.00100484 0 0.00100476 0 0.00100486 3.3 0.0010047799999999998 3.3 0.0010048799999999999 0 0.0010048 0 0.0010049 3.3 0.00100482 3.3 0.00100492 0 0.00100484 0 0.00100494 3.3 0.00100486 3.3 0.00100496 0 0.0010048799999999999 0 0.00100498 3.3 0.0010049 3.3 0.001005 0 0.0010049199999999999 0 0.00100502 3.3 0.00100494 3.3 0.00100504 0 0.0010049599999999998 0 0.00100506 3.3 0.00100498 3.3 0.00100508 0 0.0010049999999999998 0 0.0010050999999999999 3.3 0.00100502 3.3 0.00100512 0 0.00100504 0 0.00100514 3.3 0.00100506 3.3 0.00100516 0 0.00100508 0 0.00100518 3.3 0.0010050999999999999 3.3 0.0010052 0 0.00100512 0 0.00100522 3.3 0.0010051399999999999 3.3 0.00100524 0 0.00100516 0 0.00100526 3.3 0.0010051799999999998 3.3 0.0010052799999999999 0 0.0010052 0 0.0010053 3.3 0.00100522 3.3 0.00100532 0 0.00100524 0 0.00100534 3.3 0.00100526 3.3 0.00100536 0 0.0010052799999999999 0 0.00100538 3.3 0.0010053 3.3 0.0010054 0 0.0010053199999999999 0 0.00100542 3.3 0.00100534 3.3 0.00100544 0 0.0010053599999999998 0 0.00100546 3.3 0.00100538 3.3 0.00100548 0 0.0010053999999999998 0 0.0010054999999999999 3.3 0.00100542 3.3 0.00100552 0 0.00100544 0 0.00100554 3.3 0.00100546 3.3 0.00100556 0 0.00100548 0 0.00100558 3.3 0.0010054999999999999 3.3 0.0010056 0 0.00100552 0 0.00100562 3.3 0.0010055399999999999 3.3 0.00100564 0 0.00100556 0 0.00100566 3.3 0.0010055799999999998 3.3 0.00100568 0 0.0010056 0 0.0010057 3.3 0.0010056199999999998 3.3 0.0010057199999999999 0 0.00100564 0 0.00100574 3.3 0.00100566 3.3 0.00100576 0 0.00100568 0 0.00100578 3.3 0.0010057 3.3 0.0010058 0 0.0010057199999999999 0 0.00100582 3.3 0.00100574 3.3 0.00100584 0 0.0010057599999999999 0 0.00100586 3.3 0.00100578 3.3 0.00100588 0 0.0010057999999999998 0 0.0010059 3.3 0.00100582 3.3 0.00100592 0 0.0010058399999999998 0 0.0010059399999999999 3.3 0.00100586 3.3 0.00100596 0 0.00100588 0 0.00100598 3.3 0.0010059 3.3 0.001006 0 0.00100592 0 0.00100602 3.3 0.0010059399999999999 3.3 0.00100604 0 0.00100596 0 0.00100606 3.3 0.0010059799999999999 3.3 0.00100608 0 0.001006 0 0.0010061 3.3 0.0010060199999999998 3.3 0.0010061199999999999 0 0.00100604 0 0.00100614 3.3 0.00100606 3.3 0.00100616 0 0.00100608 0 0.00100618 3.3 0.0010061 3.3 0.0010062 0 0.0010061199999999999 0 0.00100622 3.3 0.00100614 3.3 0.00100624 0 0.0010061599999999999 0 0.00100626 3.3 0.00100618 3.3 0.00100628 0 0.0010061999999999998 0 0.0010063 3.3 0.00100622 3.3 0.00100632 0 0.0010062399999999998 0 0.0010063399999999999 3.3 0.00100626 3.3 0.00100636 0 0.00100628 0 0.00100638 3.3 0.0010063 3.3 0.0010064 0 0.00100632 0 0.00100642 3.3 0.0010063399999999999 3.3 0.00100644 0 0.00100636 0 0.00100646 3.3 0.0010063799999999999 3.3 0.00100648 0 0.0010064 0 0.0010065 3.3 0.0010064199999999998 3.3 0.00100652 0 0.00100644 0 0.00100654 3.3 0.0010064599999999998 3.3 0.0010065599999999999 0 0.00100648 0 0.00100658 3.3 0.0010065 3.3 0.0010066 0 0.00100652 0 0.00100662 3.3 0.00100654 3.3 0.00100664 0 0.0010065599999999999 0 0.00100666 3.3 0.00100658 3.3 0.00100668 0 0.0010065999999999999 0 0.0010067 3.3 0.00100662 3.3 0.00100672 0 0.0010066399999999998 0 0.00100674 3.3 0.00100666 3.3 0.00100676 0 0.00100668 0 0.00100678 3.3 0.0010067 3.3 0.0010068 0 0.00100672 0 0.00100682 3.3 0.00100674 3.3 0.00100684 0 0.00100676 0 0.00100686 3.3 0.0010067799999999999 3.3 0.00100688 0 0.0010068 0 0.0010069 3.3 0.0010068199999999999 3.3 0.00100692 0 0.00100684 0 0.00100694 3.3 0.0010068599999999998 3.3 0.0010069599999999999 0 0.00100688 0 0.00100698 3.3 0.0010069 3.3 0.001007 0 0.00100692 0 0.00100702 3.3 0.00100694 3.3 0.00100704 0 0.0010069599999999999 0 0.00100706 3.3 0.00100698 3.3 0.00100708 0 0.0010069999999999999 0 0.0010071 3.3 0.00100702 3.3 0.00100712 0 0.0010070399999999998 0 0.00100714 3.3 0.00100706 3.3 0.00100716 0 0.0010070799999999998 0 0.0010071799999999999 3.3 0.0010071 3.3 0.0010072 0 0.00100712 0 0.00100722 3.3 0.00100714 3.3 0.00100724 0 0.00100716 0 0.00100726 3.3 0.0010071799999999999 3.3 0.00100728 0 0.0010072 0 0.0010073 3.3 0.0010072199999999999 3.3 0.00100732 0 0.00100724 0 0.00100734 3.3 0.0010072599999999998 3.3 0.00100736 0 0.00100728 0 0.00100738 3.3 0.0010072999999999998 3.3 0.0010073999999999999 0 0.00100732 0 0.00100742 3.3 0.00100734 3.3 0.00100744 0 0.00100736 0 0.00100746 3.3 0.00100738 3.3 0.00100748 0 0.0010073999999999999 0 0.0010075 3.3 0.00100742 3.3 0.00100752 0 0.0010074399999999999 0 0.00100754 3.3 0.00100746 3.3 0.00100756 0 0.0010074799999999998 0 0.0010075799999999999 3.3 0.0010075 3.3 0.0010076 0 0.00100752 0 0.00100762 3.3 0.00100754 3.3 0.00100764 0 0.00100756 0 0.00100766 3.3 0.0010075799999999999 3.3 0.00100768 0 0.0010076 0 0.0010077 3.3 0.0010076199999999999 3.3 0.00100772 0 0.00100764 0 0.00100774 3.3 0.0010076599999999998 3.3 0.00100776 0 0.00100768 0 0.00100778 3.3 0.0010076999999999998 3.3 0.0010077999999999999 0 0.00100772 0 0.00100782 3.3 0.00100774 3.3 0.00100784 0 0.00100776 0 0.00100786 3.3 0.00100778 3.3 0.00100788 0 0.0010077999999999999 0 0.0010079 3.3 0.00100782 3.3 0.00100792 0 0.0010078399999999999 0 0.00100794 3.3 0.00100786 3.3 0.00100796 0 0.0010078799999999998 0 0.00100798 3.3 0.0010079 3.3 0.001008 0 0.0010079199999999998 0 0.0010080199999999999 3.3 0.00100794 3.3 0.00100804 0 0.00100796 0 0.00100806 3.3 0.00100798 3.3 0.00100808 0 0.001008 0 0.0010081 3.3 0.0010080199999999999 3.3 0.00100812 0 0.00100804 0 0.00100814 3.3 0.0010080599999999999 3.3 0.00100816 0 0.00100808 0 0.00100818 3.3 0.0010080999999999998 3.3 0.0010082 0 0.00100812 0 0.00100822 3.3 0.0010081399999999998 3.3 0.0010082399999999999 0 0.00100816 0 0.00100826 3.3 0.00100818 3.3 0.00100828 0 0.0010082 0 0.0010083 3.3 0.00100822 3.3 0.00100832 0 0.0010082399999999999 0 0.00100834 3.3 0.00100826 3.3 0.00100836 0 0.0010082799999999999 0 0.00100838 3.3 0.0010083 3.3 0.0010084 0 0.0010083199999999998 0 0.0010084199999999999 3.3 0.00100834 3.3 0.00100844 0 0.00100836 0 0.00100846 3.3 0.00100838 3.3 0.00100848 0 0.0010084 0 0.0010085 3.3 0.0010084199999999999 3.3 0.00100852 0 0.00100844 0 0.00100854 3.3 0.0010084599999999999 3.3 0.00100856 0 0.00100848 0 0.00100858 3.3 0.0010084999999999998 3.3 0.0010086 0 0.00100852 0 0.00100862 3.3 0.0010085399999999998 3.3 0.0010086399999999999 0 0.00100856 0 0.00100866 3.3 0.00100858 3.3 0.00100868 0 0.0010086 0 0.0010087 3.3 0.00100862 3.3 0.00100872 0 0.0010086399999999999 0 0.00100874 3.3 0.00100866 3.3 0.00100876 0 0.0010086799999999999 0 0.00100878 3.3 0.0010087 3.3 0.0010088 0 0.0010087199999999998 0 0.00100882 3.3 0.00100874 3.3 0.00100884 0 0.0010087599999999998 0 0.0010088599999999999 3.3 0.00100878 3.3 0.00100888 0 0.0010088 0 0.0010089 3.3 0.00100882 3.3 0.00100892 0 0.00100884 0 0.00100894 3.3 0.0010088599999999999 3.3 0.00100896 0 0.00100888 0 0.00100898 3.3 0.0010088999999999999 3.3 0.001009 0 0.00100892 0 0.00100902 3.3 0.0010089399999999998 3.3 0.00100904 0 0.00100896 0 0.00100906 3.3 0.0010089799999999998 3.3 0.0010090799999999999 0 0.001009 0 0.0010091 3.3 0.00100902 3.3 0.00100912 0 0.00100904 0 0.00100914 3.3 0.00100906 3.3 0.00100916 0 0.0010090799999999999 0 0.00100918 3.3 0.0010091 3.3 0.0010092 0 0.0010091199999999999 0 0.00100922 3.3 0.00100914 3.3 0.00100924 0 0.0010091599999999998 0 0.0010092599999999999 3.3 0.00100918 3.3 0.00100928 0 0.0010092 0 0.0010093 3.3 0.00100922 3.3 0.00100932 0 0.00100924 0 0.00100934 3.3 0.0010092599999999999 3.3 0.00100936 0 0.00100928 0 0.00100938 3.3 0.0010092999999999999 3.3 0.0010094 0 0.00100932 0 0.00100942 3.3 0.0010093399999999998 3.3 0.00100944 0 0.00100936 0 0.00100946 3.3 0.0010093799999999998 3.3 0.0010094799999999999 0 0.0010094 0 0.0010095 3.3 0.00100942 3.3 0.00100952 0 0.00100944 0 0.00100954 3.3 0.00100946 3.3 0.00100956 0 0.0010094799999999999 0 0.00100958 3.3 0.0010095 3.3 0.0010096 0 0.0010095199999999999 0 0.00100962 3.3 0.00100954 3.3 0.00100964 0 0.0010095599999999998 0 0.00100966 3.3 0.00100958 3.3 0.00100968 0 0.0010095999999999998 0 0.0010096999999999999 3.3 0.00100962 3.3 0.00100972 0 0.00100964 0 0.00100974 3.3 0.00100966 3.3 0.00100976 0 0.00100968 0 0.00100978 3.3 0.0010096999999999999 3.3 0.0010098 0 0.00100972 0 0.00100982 3.3 0.0010097399999999999 3.3 0.00100984 0 0.00100976 0 0.00100986 3.3 0.0010097799999999998 3.3 0.00100988 0 0.0010098 0 0.0010099 3.3 0.0010098199999999998 3.3 0.0010099199999999999 0 0.00100984 0 0.00100994 3.3 0.00100986 3.3 0.00100996 0 0.00100988 0 0.00100998 3.3 0.0010099 3.3 0.00101 0 0.0010099199999999999 0 0.00101002 3.3 0.00100994 3.3 0.00101004 0 0.0010099599999999999 0 0.00101006 3.3 0.00100998 3.3 0.00101008 0 0.0010099999999999998 0 0.0010100999999999999 3.3 0.00101002 3.3 0.00101012 0 0.00101004 0 0.00101014 3.3 0.00101006 3.3 0.00101016 0 0.00101008 0 0.00101018 3.3 0.0010100999999999999 3.3 0.0010102 0 0.00101012 0 0.00101022 3.3 0.0010101399999999999 3.3 0.00101024 0 0.00101016 0 0.00101026 3.3 0.0010101799999999998 3.3 0.00101028 0 0.0010102 0 0.0010103 3.3 0.0010102199999999998 3.3 0.0010103199999999999 0 0.00101024 0 0.00101034 3.3 0.00101026 3.3 0.00101036 0 0.00101028 0 0.00101038 3.3 0.0010103 3.3 0.0010104 0 0.0010103199999999999 0 0.00101042 3.3 0.00101034 3.3 0.00101044 0 0.0010103599999999999 0 0.00101046 3.3 0.00101038 3.3 0.00101048 0 0.0010103999999999998 0 0.0010105 3.3 0.00101042 3.3 0.00101052 0 0.0010104399999999998 0 0.0010105399999999999 3.3 0.00101046 3.3 0.00101056 0 0.00101048 0 0.00101058 3.3 0.0010105 3.3 0.0010106 0 0.00101052 0 0.00101062 3.3 0.0010105399999999999 3.3 0.00101064 0 0.00101056 0 0.00101066 3.3 0.0010105799999999999 3.3 0.00101068 0 0.0010106 0 0.0010107 3.3 0.0010106199999999998 3.3 0.0010107199999999999 0 0.00101064 0 0.00101074 3.3 0.00101066 3.3 0.00101076 0 0.00101068 0 0.00101078 3.3 0.0010107 3.3 0.0010108 0 0.0010107199999999999 0 0.00101082 3.3 0.00101074 3.3 0.00101084 0 0.0010107599999999999 0 0.00101086 3.3 0.00101078 3.3 0.00101088 0 0.0010107999999999998 0 0.0010109 3.3 0.00101082 3.3 0.00101092 0 0.0010108399999999998 0 0.0010109399999999999 3.3 0.00101086 3.3 0.00101096 0 0.00101088 0 0.00101098 3.3 0.0010109 3.3 0.001011 0 0.00101092 0 0.00101102 3.3 0.0010109399999999999 3.3 0.00101104 0 0.00101096 0 0.00101106 3.3 0.0010109799999999999 3.3 0.00101108 0 0.001011 0 0.0010111 3.3 0.0010110199999999998 3.3 0.00101112 0 0.00101104 0 0.00101114 3.3 0.0010110599999999998 3.3 0.0010111599999999999 0 0.00101108 0 0.00101118 3.3 0.0010111 3.3 0.0010112 0 0.00101112 0 0.00101122 3.3 0.00101114 3.3 0.00101124 0 0.0010111599999999999 0 0.00101126 3.3 0.00101118 3.3 0.00101128 0 0.0010111999999999999 0 0.0010113 3.3 0.00101122 3.3 0.00101132 0 0.0010112399999999998 0 0.00101134 3.3 0.00101126 3.3 0.00101136 0 0.0010112799999999998 0 0.0010113799999999999 3.3 0.0010113 3.3 0.0010114 0 0.00101132 0 0.00101142 3.3 0.00101134 3.3 0.00101144 0 0.00101136 0 0.00101146 3.3 0.0010113799999999999 3.3 0.00101148 0 0.0010114 0 0.0010115 3.3 0.0010114199999999999 3.3 0.00101152 0 0.00101144 0 0.00101154 3.3 0.0010114599999999998 3.3 0.0010115599999999999 0 0.00101148 0 0.00101158 3.3 0.0010115 3.3 0.0010116 0 0.00101152 0 0.00101162 3.3 0.00101154 3.3 0.00101164 0 0.0010115599999999999 0 0.00101166 3.3 0.00101158 3.3 0.00101168 0 0.0010115999999999999 0 0.0010117 3.3 0.00101162 3.3 0.00101172 0 0.0010116399999999998 0 0.00101174 3.3 0.00101166 3.3 0.00101176 0 0.0010116799999999998 0 0.0010117799999999999 3.3 0.0010117 3.3 0.0010118 0 0.00101172 0 0.00101182 3.3 0.00101174 3.3 0.00101184 0 0.00101176 0 0.00101186 3.3 0.0010117799999999999 3.3 0.00101188 0 0.0010118 0 0.0010119 3.3 0.0010118199999999999 3.3 0.00101192 0 0.00101184 0 0.00101194 3.3 0.0010118599999999998 3.3 0.00101196 0 0.00101188 0 0.00101198 3.3 0.0010118999999999998 3.3 0.0010119999999999999 0 0.00101192 0 0.00101202 3.3 0.00101194 3.3 0.00101204 0 0.00101196 0 0.00101206 3.3 0.00101198 3.3 0.00101208 0 0.0010119999999999999 0 0.0010121 3.3 0.00101202 3.3 0.00101212 0 0.0010120399999999999 0 0.00101214 3.3 0.00101206 3.3 0.00101216 0 0.0010120799999999998 0 0.00101218 3.3 0.0010121 3.3 0.0010122 0 0.0010121199999999998 0 0.0010122199999999999 3.3 0.00101214 3.3 0.00101224 0 0.00101216 0 0.00101226 3.3 0.00101218 3.3 0.00101228 0 0.0010122 0 0.0010123 3.3 0.0010122199999999999 3.3 0.00101232 0 0.00101224 0 0.00101234 3.3 0.0010122599999999999 3.3 0.00101236 0 0.00101228 0 0.00101238 3.3 0.0010122999999999998 3.3 0.0010123999999999999 0 0.00101232 0 0.00101242 3.3 0.00101234 3.3 0.00101244 0 0.00101236 0 0.00101246 3.3 0.00101238 3.3 0.00101248 0 0.0010123999999999999 0 0.0010125 3.3 0.00101242 3.3 0.00101252 0 0.0010124399999999999 0 0.00101254 3.3 0.00101246 3.3 0.00101256 0 0.0010124799999999998 0 0.00101258 3.3 0.0010125 3.3 0.0010126 0 0.0010125199999999998 0 0.0010126199999999999 3.3 0.00101254 3.3 0.00101264 0 0.00101256 0 0.00101266 3.3 0.00101258 3.3 0.00101268 0 0.0010126 0 0.0010127 3.3 0.0010126199999999999 3.3 0.00101272 0 0.00101264 0 0.00101274 3.3 0.0010126599999999999 3.3 0.00101276 0 0.00101268 0 0.00101278 3.3 0.0010126999999999998 3.3 0.0010128 0 0.00101272 0 0.00101282 3.3 0.0010127399999999998 3.3 0.0010128399999999999 0 0.00101276 0 0.00101286 3.3 0.00101278 3.3 0.00101288 0 0.0010128 0 0.0010129 3.3 0.00101282 3.3 0.00101292 0 0.0010128399999999999 0 0.00101294 3.3 0.00101286 3.3 0.00101296 0 0.0010128799999999999 0 0.00101298 3.3 0.0010129 3.3 0.001013 0 0.0010129199999999998 0 0.00101302 3.3 0.00101294 3.3 0.00101304 0 0.0010129599999999998 0 0.0010130599999999999 3.3 0.00101298 3.3 0.00101308 0 0.001013 0 0.0010131 3.3 0.00101302 3.3 0.00101312 0 0.00101304 0 0.00101314 3.3 0.0010130599999999999 3.3 0.00101316 0 0.00101308 0 0.00101318 3.3 0.0010130999999999999 3.3 0.0010132 0 0.00101312 0 0.00101322 3.3 0.0010131399999999998 3.3 0.0010132399999999999 0 0.00101316 0 0.00101326 3.3 0.00101318 3.3 0.00101328 0 0.0010132 0 0.0010133 3.3 0.00101322 3.3 0.00101332 0 0.0010132399999999999 0 0.00101334 3.3 0.00101326 3.3 0.00101336 0 0.0010132799999999999 0 0.00101338 3.3 0.0010133 3.3 0.0010134 0 0.0010133199999999998 0 0.00101342 3.3 0.00101334 3.3 0.00101344 0 0.0010133599999999998 0 0.0010134599999999999 3.3 0.00101338 3.3 0.00101348 0 0.0010134 0 0.0010135 3.3 0.00101342 3.3 0.00101352 0 0.00101344 0 0.00101354 3.3 0.0010134599999999999 3.3 0.00101356 0 0.00101348 0 0.00101358 3.3 0.0010134999999999999 3.3 0.0010136 0 0.00101352 0 0.00101362 3.3 0.0010135399999999998 3.3 0.00101364 0 0.00101356 0 0.00101366 3.3 0.0010135799999999998 3.3 0.0010136799999999999 0 0.0010136 0 0.0010137 3.3 0.00101362 3.3 0.00101372 0 0.00101364 0 0.00101374 3.3 0.00101366 3.3 0.00101376 0 0.0010136799999999999 0 0.00101378 3.3 0.0010137 3.3 0.0010138 0 0.0010137199999999999 0 0.00101382 3.3 0.00101374 3.3 0.00101384 0 0.0010137599999999998 0 0.0010138599999999999 3.3 0.00101378 3.3 0.00101388 0 0.0010138 0 0.0010139 3.3 0.00101382 3.3 0.00101392 0 0.00101384 0 0.00101394 3.3 0.0010138599999999999 3.3 0.00101396 0 0.00101388 0 0.00101398 3.3 0.0010138999999999999 3.3 0.001014 0 0.00101392 0 0.00101402 3.3 0.0010139399999999999 3.3 0.00101404 0 0.00101396 0 0.00101406 3.3 0.0010139799999999998 3.3 0.0010140799999999999 0 0.001014 0 0.0010141 3.3 0.00101402 3.3 0.00101412 0 0.00101404 0 0.00101414 3.3 0.00101406 3.3 0.00101416 0 0.0010140799999999999 0 0.00101418 3.3 0.0010141 3.3 0.0010142 0 0.0010141199999999999 0 0.00101422 3.3 0.00101414 3.3 0.00101424 0 0.0010141599999999998 0 0.00101426 3.3 0.00101418 3.3 0.00101428 0 0.0010141999999999998 0 0.0010142999999999999 3.3 0.00101422 3.3 0.00101432 0 0.00101424 0 0.00101434 3.3 0.00101426 3.3 0.00101436 0 0.00101428 0 0.00101438 3.3 0.0010142999999999999 3.3 0.0010144 0 0.00101432 0 0.00101442 3.3 0.0010143399999999999 3.3 0.00101444 0 0.00101436 0 0.00101446 3.3 0.0010143799999999998 3.3 0.00101448 0 0.0010144 0 0.0010145 3.3 0.0010144199999999998 3.3 0.0010145199999999999 0 0.00101444 0 0.00101454 3.3 0.00101446 3.3 0.00101456 0 0.00101448 0 0.00101458 3.3 0.0010145 3.3 0.0010146 0 0.0010145199999999999 0 0.00101462 3.3 0.00101454 3.3 0.00101464 0 0.0010145599999999999 0 0.00101466 3.3 0.00101458 3.3 0.00101468 0 0.0010145999999999998 0 0.0010146999999999999 3.3 0.00101462 3.3 0.00101472 0 0.00101464 0 0.00101474 3.3 0.00101466 3.3 0.00101476 0 0.00101468 0 0.00101478 3.3 0.0010146999999999999 3.3 0.0010148 0 0.00101472 0 0.00101482 3.3 0.0010147399999999999 3.3 0.00101484 0 0.00101476 0 0.00101486 3.3 0.0010147799999999998 3.3 0.00101488 0 0.0010148 0 0.0010149 3.3 0.0010148199999999998 3.3 0.0010149199999999999 0 0.00101484 0 0.00101494 3.3 0.00101486 3.3 0.00101496 0 0.00101488 0 0.00101498 3.3 0.0010149 3.3 0.001015 0 0.0010149199999999999 0 0.00101502 3.3 0.00101494 3.3 0.00101504 0 0.0010149599999999999 0 0.00101506 3.3 0.00101498 3.3 0.00101508 0 0.0010149999999999998 0 0.0010151 3.3 0.00101502 3.3 0.00101512 0 0.0010150399999999998 0 0.0010151399999999999 3.3 0.00101506 3.3 0.00101516 0 0.00101508 0 0.00101518 3.3 0.0010151 3.3 0.0010152 0 0.00101512 0 0.00101522 3.3 0.0010151399999999999 3.3 0.00101524 0 0.00101516 0 0.00101526 3.3 0.0010151799999999999 3.3 0.00101528 0 0.0010152 0 0.0010153 3.3 0.0010152199999999998 3.3 0.00101532 0 0.00101524 0 0.00101534 3.3 0.0010152599999999998 3.3 0.0010153599999999999 0 0.00101528 0 0.00101538 3.3 0.0010153 3.3 0.0010154 0 0.00101532 0 0.00101542 3.3 0.00101534 3.3 0.00101544 0 0.0010153599999999999 0 0.00101546 3.3 0.00101538 3.3 0.00101548 0 0.0010153999999999999 0 0.0010155 3.3 0.00101542 3.3 0.00101552 0 0.0010154399999999998 0 0.0010155399999999999 3.3 0.00101546 3.3 0.00101556 0 0.00101548 0 0.00101558 3.3 0.0010155 3.3 0.0010156 0 0.00101552 0 0.00101562 3.3 0.0010155399999999999 3.3 0.00101564 0 0.00101556 0 0.00101566 3.3 0.0010155799999999999 3.3 0.00101568 0 0.0010156 0 0.0010157 3.3 0.0010156199999999998 3.3 0.00101572 0 0.00101564 0 0.00101574 3.3 0.0010156599999999998 3.3 0.0010157599999999999 0 0.00101568 0 0.00101578 3.3 0.0010157 3.3 0.0010158 0 0.00101572 0 0.00101582 3.3 0.00101574 3.3 0.00101584 0 0.0010157599999999999 0 0.00101586 3.3 0.00101578 3.3 0.00101588 0 0.0010157999999999999 0 0.0010159 3.3 0.00101582 3.3 0.00101592 0 0.0010158399999999998 0 0.00101594 3.3 0.00101586 3.3 0.00101596 0 0.0010158799999999998 0 0.0010159799999999999 3.3 0.0010159 3.3 0.001016 0 0.00101592 0 0.00101602 3.3 0.00101594 3.3 0.00101604 0 0.00101596 0 0.00101606 3.3 0.0010159799999999999 3.3 0.00101608 0 0.001016 0 0.0010161 3.3 0.0010160199999999999 3.3 0.00101612 0 0.00101604 0 0.00101614 3.3 0.0010160599999999998 3.3 0.00101616 0 0.00101608 0 0.00101618 3.3 0.0010160999999999998 3.3 0.0010161999999999999 0 0.00101612 0 0.00101622 3.3 0.00101614 3.3 0.00101624 0 0.00101616 0 0.00101626 3.3 0.00101618 3.3 0.00101628 0 0.0010161999999999999 0 0.0010163 3.3 0.00101622 3.3 0.00101632 0 0.0010162399999999999 0 0.00101634 3.3 0.00101626 3.3 0.00101636 0 0.0010162799999999998 0 0.0010163799999999999 3.3 0.0010163 3.3 0.0010164 0 0.00101632 0 0.00101642 3.3 0.00101634 3.3 0.00101644 0 0.00101636 0 0.00101646 3.3 0.0010163799999999999 3.3 0.00101648 0 0.0010164 0 0.0010165 3.3 0.0010164199999999999 3.3 0.00101652 0 0.00101644 0 0.00101654 3.3 0.0010164599999999998 3.3 0.00101656 0 0.00101648 0 0.00101658 3.3 0.0010164999999999998 3.3 0.0010165999999999999 0 0.00101652 0 0.00101662 3.3 0.00101654 3.3 0.00101664 0 0.00101656 0 0.00101666 3.3 0.00101658 3.3 0.00101668 0 0.0010165999999999999 0 0.0010167 3.3 0.00101662 3.3 0.00101672 0 0.0010166399999999999 0 0.00101674 3.3 0.00101666 3.3 0.00101676 0 0.0010166799999999998 0 0.00101678 3.3 0.0010167 3.3 0.0010168 0 0.0010167199999999998 0 0.0010168199999999999 3.3 0.00101674 3.3 0.00101684 0 0.00101676 0 0.00101686 3.3 0.00101678 3.3 0.00101688 0 0.0010168 0 0.0010169 3.3 0.0010168199999999999 3.3 0.00101692 0 0.00101684 0 0.00101694 3.3 0.0010168599999999999 3.3 0.00101696 0 0.00101688 0 0.00101698 3.3 0.0010168999999999998 3.3 0.001017 0 0.00101692 0 0.00101702 3.3 0.0010169399999999998 3.3 0.0010170399999999999 0 0.00101696 0 0.00101706 3.3 0.00101698 3.3 0.00101708 0 0.001017 0 0.0010171 3.3 0.00101702 3.3 0.00101712 0 0.0010170399999999999 0 0.00101714 3.3 0.00101706 3.3 0.00101716 0 0.0010170799999999999 0 0.00101718 3.3 0.0010171 3.3 0.0010172 0 0.0010171199999999998 0 0.0010172199999999999 3.3 0.00101714 3.3 0.00101724 0 0.00101716 0 0.00101726 3.3 0.00101718 3.3 0.00101728 0 0.0010172 0 0.0010173 3.3 0.0010172199999999999 3.3 0.00101732 0 0.00101724 0 0.00101734 3.3 0.0010172599999999999 3.3 0.00101736 0 0.00101728 0 0.00101738 3.3 0.0010172999999999998 3.3 0.0010174 0 0.00101732 0 0.00101742 3.3 0.0010173399999999998 3.3 0.0010174399999999999 0 0.00101736 0 0.00101746 3.3 0.00101738 3.3 0.00101748 0 0.0010174 0 0.0010175 3.3 0.00101742 3.3 0.00101752 0 0.0010174399999999999 0 0.00101754 3.3 0.00101746 3.3 0.00101756 0 0.0010174799999999999 0 0.00101758 3.3 0.0010175 3.3 0.0010176 0 0.0010175199999999998 0 0.00101762 3.3 0.00101754 3.3 0.00101764 0 0.0010175599999999998 0 0.0010176599999999999 3.3 0.00101758 3.3 0.00101768 0 0.0010176 0 0.0010177 3.3 0.00101762 3.3 0.00101772 0 0.00101764 0 0.00101774 3.3 0.0010176599999999999 3.3 0.00101776 0 0.00101768 0 0.00101778 3.3 0.0010176999999999999 3.3 0.0010178 0 0.00101772 0 0.00101782 3.3 0.0010177399999999998 3.3 0.0010178399999999999 0 0.00101776 0 0.00101786 3.3 0.00101778 3.3 0.00101788 0 0.0010178 0 0.0010179 3.3 0.00101782 3.3 0.00101792 0 0.0010178399999999999 0 0.00101794 3.3 0.00101786 3.3 0.00101796 0 0.0010178799999999999 0 0.00101798 3.3 0.0010179 3.3 0.001018 0 0.0010179199999999998 0 0.00101802 3.3 0.00101794 3.3 0.00101804 0 0.0010179599999999998 0 0.0010180599999999999 3.3 0.00101798 3.3 0.00101808 0 0.001018 0 0.0010181 3.3 0.00101802 3.3 0.00101812 0 0.00101804 0 0.00101814 3.3 0.0010180599999999999 3.3 0.00101816 0 0.00101808 0 0.00101818 3.3 0.0010180999999999999 3.3 0.0010182 0 0.00101812 0 0.00101822 3.3 0.0010181399999999998 3.3 0.00101824 0 0.00101816 0 0.00101826 3.3 0.0010181799999999998 3.3 0.0010182799999999999 0 0.0010182 0 0.0010183 3.3 0.00101822 3.3 0.00101832 0 0.00101824 0 0.00101834 3.3 0.00101826 3.3 0.00101836 0 0.0010182799999999999 0 0.00101838 3.3 0.0010183 3.3 0.0010184 0 0.0010183199999999999 0 0.00101842 3.3 0.00101834 3.3 0.00101844 0 0.0010183599999999998 0 0.00101846 3.3 0.00101838 3.3 0.00101848 0 0.0010183999999999998 0 0.0010184999999999999 3.3 0.00101842 3.3 0.00101852 0 0.00101844 0 0.00101854 3.3 0.00101846 3.3 0.00101856 0 0.00101848 0 0.00101858 3.3 0.0010184999999999999 3.3 0.0010186 0 0.00101852 0 0.00101862 3.3 0.0010185399999999999 3.3 0.00101864 0 0.00101856 0 0.00101866 3.3 0.0010185799999999998 3.3 0.0010186799999999999 0 0.0010186 0 0.0010187 3.3 0.00101862 3.3 0.00101872 0 0.00101864 0 0.00101874 3.3 0.00101866 3.3 0.00101876 0 0.0010186799999999999 0 0.00101878 3.3 0.0010187 3.3 0.0010188 0 0.0010187199999999999 0 0.00101882 3.3 0.00101874 3.3 0.00101884 0 0.0010187599999999998 0 0.00101886 3.3 0.00101878 3.3 0.00101888 0 0.0010187999999999998 0 0.0010188999999999999 3.3 0.00101882 3.3 0.00101892 0 0.00101884 0 0.00101894 3.3 0.00101886 3.3 0.00101896 0 0.00101888 0 0.00101898 3.3 0.0010188999999999999 3.3 0.001019 0 0.00101892 0 0.00101902 3.3 0.0010189399999999999 3.3 0.00101904 0 0.00101896 0 0.00101906 3.3 0.0010189799999999998 3.3 0.00101908 0 0.001019 0 0.0010191 3.3 0.0010190199999999998 3.3 0.0010191199999999999 0 0.00101904 0 0.00101914 3.3 0.00101906 3.3 0.00101916 0 0.00101908 0 0.00101918 3.3 0.0010191 3.3 0.0010192 0 0.0010191199999999999 0 0.00101922 3.3 0.00101914 3.3 0.00101924 0 0.0010191599999999999 0 0.00101926 3.3 0.00101918 3.3 0.00101928 0 0.0010191999999999998 0 0.0010193 3.3 0.00101922 3.3 0.00101932 0 0.0010192399999999998 0 0.0010193399999999999 3.3 0.00101926 3.3 0.00101936 0 0.00101928 0 0.00101938 3.3 0.0010193 3.3 0.0010194 0 0.00101932 0 0.00101942 3.3 0.0010193399999999999 3.3 0.00101944 0 0.00101936 0 0.00101946 3.3 0.0010193799999999999 3.3 0.00101948 0 0.0010194 0 0.0010195 3.3 0.0010194199999999998 3.3 0.0010195199999999999 0 0.00101944 0 0.00101954 3.3 0.00101946 3.3 0.00101956 0 0.00101948 0 0.00101958 3.3 0.0010195 3.3 0.0010196 0 0.0010195199999999999 0 0.00101962 3.3 0.00101954 3.3 0.00101964 0 0.0010195599999999999 0 0.00101966 3.3 0.00101958 3.3 0.00101968 0 0.0010195999999999998 0 0.0010197 3.3 0.00101962 3.3 0.00101972 0 0.0010196399999999998 0 0.0010197399999999999 3.3 0.00101966 3.3 0.00101976 0 0.00101968 0 0.00101978 3.3 0.0010197 3.3 0.0010198 0 0.00101972 0 0.00101982 3.3 0.0010197399999999999 3.3 0.00101984 0 0.00101976 0 0.00101986 3.3 0.0010197799999999999 3.3 0.00101988 0 0.0010198 0 0.0010199 3.3 0.0010198199999999998 3.3 0.00101992 0 0.00101984 0 0.00101994 3.3 0.0010198599999999998 3.3 0.0010199599999999999 0 0.00101988 0 0.00101998 3.3 0.0010199 3.3 0.00102 0 0.00101992 0 0.00102002 3.3 0.00101994 3.3 0.00102004 0 0.0010199599999999999 0 0.00102006 3.3 0.00101998 3.3 0.00102008 0 0.0010199999999999999 0 0.0010201 3.3 0.00102002 3.3 0.00102012 0 0.0010200399999999998 0 0.00102014 3.3 0.00102006 3.3 0.00102016 0 0.0010200799999999998 0 0.0010201799999999999 3.3 0.0010201 3.3 0.0010202 0 0.00102012 0 0.00102022 3.3 0.00102014 3.3 0.00102024 0 0.00102016 0 0.00102026 3.3 0.0010201799999999999 3.3 0.00102028 0 0.0010202 0 0.0010203 3.3 0.0010202199999999999 3.3 0.00102032 0 0.00102024 0 0.00102034 3.3 0.0010202599999999998 3.3 0.0010203599999999999 0 0.00102028 0 0.00102038 3.3 0.0010203 3.3 0.0010204 0 0.00102032 0 0.00102042 3.3 0.00102034 3.3 0.00102044 0 0.0010203599999999999 0 0.00102046 3.3 0.00102038 3.3 0.00102048 0 0.0010203999999999999 0 0.0010205 3.3 0.00102042 3.3 0.00102052 0 0.0010204399999999998 0 0.00102054 3.3 0.00102046 3.3 0.00102056 0 0.0010204799999999998 0 0.0010205799999999999 3.3 0.0010205 3.3 0.0010206 0 0.00102052 0 0.00102062 3.3 0.00102054 3.3 0.00102064 0 0.00102056 0 0.00102066 3.3 0.0010205799999999999 3.3 0.00102068 0 0.0010206 0 0.0010207 3.3 0.0010206199999999999 3.3 0.00102072 0 0.00102064 0 0.00102074 3.3 0.0010206599999999998 3.3 0.00102076 0 0.00102068 0 0.00102078 3.3 0.0010206999999999998 3.3 0.0010207999999999999 0 0.00102072 0 0.00102082 3.3 0.00102074 3.3 0.00102084 0 0.00102076 0 0.00102086 3.3 0.00102078 3.3 0.00102088 0 0.0010207999999999999 0 0.0010209 3.3 0.00102082 3.3 0.00102092 0 0.0010208399999999999 0 0.00102094 3.3 0.00102086 3.3 0.00102096 0 0.0010208799999999998 0 0.0010209799999999999 3.3 0.0010209 3.3 0.001021 0 0.00102092 0 0.00102102 3.3 0.00102094 3.3 0.00102104 0 0.00102096 0 0.00102106 3.3 0.0010209799999999999 3.3 0.00102108 0 0.001021 0 0.0010211 3.3 0.0010210199999999999 3.3 0.00102112 0 0.00102104 0 0.00102114 3.3 0.0010210599999999998 3.3 0.00102116 0 0.00102108 0 0.00102118 3.3 0.0010210999999999998 3.3 0.0010211999999999999 0 0.00102112 0 0.00102122 3.3 0.00102114 3.3 0.00102124 0 0.00102116 0 0.00102126 3.3 0.00102118 3.3 0.00102128 0 0.0010211999999999999 0 0.0010213 3.3 0.00102122 3.3 0.00102132 0 0.0010212399999999999 0 0.00102134 3.3 0.00102126 3.3 0.00102136 0 0.0010212799999999998 0 0.00102138 3.3 0.0010213 3.3 0.0010214 0 0.0010213199999999998 0 0.0010214199999999999 3.3 0.00102134 3.3 0.00102144 0 0.00102136 0 0.00102146 3.3 0.00102138 3.3 0.00102148 0 0.0010214 0 0.0010215 3.3 0.0010214199999999999 3.3 0.00102152 0 0.00102144 0 0.00102154 3.3 0.0010214599999999999 3.3 0.00102156 0 0.00102148 0 0.00102158 3.3 0.0010214999999999998 3.3 0.0010216 0 0.00102152 0 0.00102162 3.3 0.0010215399999999998 3.3 0.0010216399999999999 0 0.00102156 0 0.00102166 3.3 0.00102158 3.3 0.00102168 0 0.0010216 0 0.0010217 3.3 0.00102162 3.3 0.00102172 0 0.0010216399999999999 0 0.00102174 3.3 0.00102166 3.3 0.00102176 0 0.0010216799999999999 0 0.00102178 3.3 0.0010217 3.3 0.0010218 0 0.0010217199999999998 0 0.0010218199999999999 3.3 0.00102174 3.3 0.00102184 0 0.00102176 0 0.00102186 3.3 0.00102178 3.3 0.00102188 0 0.0010218 0 0.0010219 3.3 0.0010218199999999999 3.3 0.00102192 0 0.00102184 0 0.00102194 3.3 0.0010218599999999999 3.3 0.00102196 0 0.00102188 0 0.00102198 3.3 0.0010218999999999998 3.3 0.001022 0 0.00102192 0 0.00102202 3.3 0.0010219399999999998 3.3 0.0010220399999999999 0 0.00102196 0 0.00102206 3.3 0.00102198 3.3 0.00102208 0 0.001022 0 0.0010221 3.3 0.00102202 3.3 0.00102212 0 0.0010220399999999999 0 0.00102214 3.3 0.00102206 3.3 0.00102216 0 0.0010220799999999999 0 0.00102218 3.3 0.0010221 3.3 0.0010222 0 0.0010221199999999998 0 0.00102222 3.3 0.00102214 3.3 0.00102224 0 0.0010221599999999998 0 0.0010222599999999999 3.3 0.00102218 3.3 0.00102228 0 0.0010222 0 0.0010223 3.3 0.00102222 3.3 0.00102232 0 0.00102224 0 0.00102234 3.3 0.0010222599999999999 3.3 0.00102236 0 0.00102228 0 0.00102238 3.3 0.0010222999999999999 3.3 0.0010224 0 0.00102232 0 0.00102242 3.3 0.0010223399999999998 3.3 0.00102244 0 0.00102236 0 0.00102246 3.3 0.0010223799999999998 3.3 0.0010224799999999999 0 0.0010224 0 0.0010225 3.3 0.00102242 3.3 0.00102252 0 0.00102244 0 0.00102254 3.3 0.00102246 3.3 0.00102256 0 0.0010224799999999999 0 0.00102258 3.3 0.0010225 3.3 0.0010226 0 0.0010225199999999999 0 0.00102262 3.3 0.00102254 3.3 0.00102264 0 0.0010225599999999998 0 0.0010226599999999999 3.3 0.00102258 3.3 0.00102268 0 0.0010226 0 0.0010227 3.3 0.00102262 3.3 0.00102272 0 0.00102264 0 0.00102274 3.3 0.0010226599999999999 3.3 0.00102276 0 0.00102268 0 0.00102278 3.3 0.0010226999999999999 3.3 0.0010228 0 0.00102272 0 0.00102282 3.3 0.0010227399999999998 3.3 0.00102284 0 0.00102276 0 0.00102286 3.3 0.0010227799999999998 3.3 0.0010228799999999999 0 0.0010228 0 0.0010229 3.3 0.00102282 3.3 0.00102292 0 0.00102284 0 0.00102294 3.3 0.00102286 3.3 0.00102296 0 0.0010228799999999999 0 0.00102298 3.3 0.0010229 3.3 0.001023 0 0.0010229199999999999 0 0.00102302 3.3 0.00102294 3.3 0.00102304 0 0.0010229599999999998 0 0.00102306 3.3 0.00102298 3.3 0.00102308 0 0.0010229999999999998 0 0.0010230999999999999 3.3 0.00102302 3.3 0.00102312 0 0.00102304 0 0.00102314 3.3 0.00102306 3.3 0.00102316 0 0.00102308 0 0.00102318 3.3 0.0010230999999999999 3.3 0.0010232 0 0.00102312 0 0.00102322 3.3 0.0010231399999999999 3.3 0.00102324 0 0.00102316 0 0.00102326 3.3 0.0010231799999999998 3.3 0.00102328 0 0.0010232 0 0.0010233 3.3 0.0010232199999999998 3.3 0.0010233199999999999 0 0.00102324 0 0.00102334 3.3 0.00102326 3.3 0.00102336 0 0.00102328 0 0.00102338 3.3 0.0010233 3.3 0.0010234 0 0.0010233199999999999 0 0.00102342 3.3 0.00102334 3.3 0.00102344 0 0.0010233599999999999 0 0.00102346 3.3 0.00102338 3.3 0.00102348 0 0.0010233999999999998 0 0.0010234999999999999 3.3 0.00102342 3.3 0.00102352 0 0.00102344 0 0.00102354 3.3 0.00102346 3.3 0.00102356 0 0.00102348 0 0.00102358 3.3 0.0010234999999999999 3.3 0.0010236 0 0.00102352 0 0.00102362 3.3 0.0010235399999999999 3.3 0.00102364 0 0.00102356 0 0.00102366 3.3 0.0010235799999999998 3.3 0.00102368 0 0.0010236 0 0.0010237 3.3 0.0010236199999999998 3.3 0.0010237199999999999 0 0.00102364 0 0.00102374 3.3 0.00102366 3.3 0.00102376 0 0.00102368 0 0.00102378 3.3 0.0010237 3.3 0.0010238 0 0.0010237199999999999 0 0.00102382 3.3 0.00102374 3.3 0.00102384 0 0.0010237599999999999 0 0.00102386 3.3 0.00102378 3.3 0.00102388 0 0.0010237999999999998 0 0.0010239 3.3 0.00102382 3.3 0.00102392 0 0.0010238399999999998 0 0.0010239399999999999 3.3 0.00102386 3.3 0.00102396 0 0.00102388 0 0.00102398 3.3 0.0010239 3.3 0.001024 0 0.00102392 0 0.00102402 3.3 0.0010239399999999999 3.3 0.00102404 0 0.00102396 0 0.00102406 3.3 0.0010239799999999999 3.3 0.00102408 0 0.001024 0 0.0010241 3.3 0.0010240199999999998 3.3 0.0010241199999999999 0 0.00102404 0 0.00102414 3.3 0.00102406 3.3 0.00102416 0 0.00102408 0 0.00102418 3.3 0.0010241 3.3 0.0010242 0 0.0010241199999999999 0 0.00102422 3.3 0.00102414 3.3 0.00102424 0 0.0010241599999999999 0 0.00102426 3.3 0.00102418 3.3 0.00102428 0 0.0010241999999999999 0 0.0010243 3.3 0.00102422 3.3 0.00102432 0 0.0010242399999999998 0 0.0010243399999999999 3.3 0.00102426 3.3 0.00102436 0 0.00102428 0 0.00102438 3.3 0.0010243 3.3 0.0010244 0 0.00102432 0 0.00102442 3.3 0.0010243399999999999 3.3 0.00102444 0 0.00102436 0 0.00102446 3.3 0.0010243799999999999 3.3 0.00102448 0 0.0010244 0 0.0010245 3.3 0.0010244199999999998 3.3 0.00102452 0 0.00102444 0 0.00102454 3.3 0.0010244599999999998 3.3 0.0010245599999999999 0 0.00102448 0 0.00102458 3.3 0.0010245 3.3 0.0010246 0 0.00102452 0 0.00102462 3.3 0.00102454 3.3 0.00102464 0 0.0010245599999999999 0 0.00102466 3.3 0.00102458 3.3 0.00102468 0 0.0010245999999999999 0 0.0010247 3.3 0.00102462 3.3 0.00102472 0 0.0010246399999999998 0 0.00102474 3.3 0.00102466 3.3 0.00102476 0 0.0010246799999999998 0 0.0010247799999999999 3.3 0.0010247 3.3 0.0010248 0 0.00102472 0 0.00102482 3.3 0.00102474 3.3 0.00102484 0 0.00102476 0 0.00102486 3.3 0.0010247799999999999 3.3 0.00102488 0 0.0010248 0 0.0010249 3.3 0.0010248199999999999 3.3 0.00102492 0 0.00102484 0 0.00102494 3.3 0.0010248599999999998 3.3 0.0010249599999999999 0 0.00102488 0 0.00102498 3.3 0.0010249 3.3 0.001025 0 0.00102492 0 0.00102502 3.3 0.00102494 3.3 0.00102504 0 0.0010249599999999999 0 0.00102506 3.3 0.00102498 3.3 0.00102508 0 0.0010249999999999999 0 0.0010251 3.3 0.00102502 3.3 0.00102512 0 0.0010250399999999998 0 0.00102514 3.3 0.00102506 3.3 0.00102516 0 0.0010250799999999998 0 0.0010251799999999999 3.3 0.0010251 3.3 0.0010252 0 0.00102512 0 0.00102522 3.3 0.00102514 3.3 0.00102524 0 0.00102516 0 0.00102526 3.3 0.0010251799999999999 3.3 0.00102528 0 0.0010252 0 0.0010253 3.3 0.0010252199999999999 3.3 0.00102532 0 0.00102524 0 0.00102534 3.3 0.0010252599999999998 3.3 0.00102536 0 0.00102528 0 0.00102538 3.3 0.0010252999999999998 3.3 0.0010253999999999999 0 0.00102532 0 0.00102542 3.3 0.00102534 3.3 0.00102544 0 0.00102536 0 0.00102546 3.3 0.00102538 3.3 0.00102548 0 0.0010253999999999999 0 0.0010255 3.3 0.00102542 3.3 0.00102552 0 0.0010254399999999999 0 0.00102554 3.3 0.00102546 3.3 0.00102556 0 0.0010254799999999998 0 0.00102558 3.3 0.0010255 3.3 0.0010256 0 0.0010255199999999998 0 0.0010256199999999999 3.3 0.00102554 3.3 0.00102564 0 0.00102556 0 0.00102566 3.3 0.00102558 3.3 0.00102568 0 0.0010256 0 0.0010257 3.3 0.0010256199999999999 3.3 0.00102572 0 0.00102564 0 0.00102574 3.3 0.0010256599999999999 3.3 0.00102576 0 0.00102568 0 0.00102578 3.3 0.0010256999999999998 3.3 0.0010257999999999999 0 0.00102572 0 0.00102582 3.3 0.00102574 3.3 0.00102584 0 0.00102576 0 0.00102586 3.3 0.00102578 3.3 0.00102588 0 0.0010257999999999999 0 0.0010259 3.3 0.00102582 3.3 0.00102592 0 0.0010258399999999999 0 0.00102594 3.3 0.00102586 3.3 0.00102596 0 0.0010258799999999998 0 0.00102598 3.3 0.0010259 3.3 0.001026 0 0.0010259199999999998 0 0.0010260199999999999 3.3 0.00102594 3.3 0.00102604 0 0.00102596 0 0.00102606 3.3 0.00102598 3.3 0.00102608 0 0.001026 0 0.0010261 3.3 0.0010260199999999999 3.3 0.00102612 0 0.00102604 0 0.00102614 3.3 0.0010260599999999999 3.3 0.00102616 0 0.00102608 0 0.00102618 3.3 0.0010260999999999998 3.3 0.0010262 0 0.00102612 0 0.00102622 3.3 0.0010261399999999998 3.3 0.0010262399999999999 0 0.00102616 0 0.00102626 3.3 0.00102618 3.3 0.00102628 0 0.0010262 0 0.0010263 3.3 0.00102622 3.3 0.00102632 0 0.0010262399999999999 0 0.00102634 3.3 0.00102626 3.3 0.00102636 0 0.0010262799999999999 0 0.00102638 3.3 0.0010263 3.3 0.0010264 0 0.0010263199999999998 0 0.00102642 3.3 0.00102634 3.3 0.00102644 0 0.0010263599999999998 0 0.0010264599999999999 3.3 0.00102638 3.3 0.00102648 0 0.0010264 0 0.0010265 3.3 0.00102642 3.3 0.00102652 0 0.00102644 0 0.00102654 3.3 0.0010264599999999999 3.3 0.00102656 0 0.00102648 0 0.00102658 3.3 0.0010264999999999999 3.3 0.0010266 0 0.00102652 0 0.00102662 3.3 0.0010265399999999998 3.3 0.0010266399999999999 0 0.00102656 0 0.00102666 3.3 0.00102658 3.3 0.00102668 0 0.0010266 0 0.0010267 3.3 0.00102662 3.3 0.00102672 0 0.0010266399999999999 0 0.00102674 3.3 0.00102666 3.3 0.00102676 0 0.0010266799999999999 0 0.00102678 3.3 0.0010267 3.3 0.0010268 0 0.0010267199999999998 0 0.00102682 3.3 0.00102674 3.3 0.00102684 0 0.0010267599999999998 0 0.0010268599999999999 3.3 0.00102678 3.3 0.00102688 0 0.0010268 0 0.0010269 3.3 0.00102682 3.3 0.00102692 0 0.00102684 0 0.00102694 3.3 0.0010268599999999999 3.3 0.00102696 0 0.00102688 0 0.00102698 3.3 0.0010268999999999999 3.3 0.001027 0 0.00102692 0 0.00102702 3.3 0.0010269399999999998 3.3 0.00102704 0 0.00102696 0 0.00102706 3.3 0.0010269799999999998 3.3 0.0010270799999999999 0 0.001027 0 0.0010271 3.3 0.00102702 3.3 0.00102712 0 0.00102704 0 0.00102714 3.3 0.00102706 3.3 0.00102716 0 0.0010270799999999999 0 0.00102718 3.3 0.0010271 3.3 0.0010272 0 0.0010271199999999999 0 0.00102722 3.3 0.00102714 3.3 0.00102724 0 0.0010271599999999998 0 0.00102726 3.3 0.00102718 3.3 0.00102728 0 0.0010271999999999998 0 0.0010272999999999999 3.3 0.00102722 3.3 0.00102732 0 0.00102724 0 0.00102734 3.3 0.00102726 3.3 0.00102736 0 0.00102728 0 0.00102738 3.3 0.0010272999999999999 3.3 0.0010274 0 0.00102732 0 0.00102742 3.3 0.0010273399999999999 3.3 0.00102744 0 0.00102736 0 0.00102746 3.3 0.0010273799999999998 3.3 0.0010274799999999999 0 0.0010274 0 0.0010275 3.3 0.00102742 3.3 0.00102752 0 0.00102744 0 0.00102754 3.3 0.00102746 3.3 0.00102756 0 0.0010274799999999999 0 0.00102758 3.3 0.0010275 3.3 0.0010276 0 0.0010275199999999999 0 0.00102762 3.3 0.00102754 3.3 0.00102764 0 0.0010275599999999998 0 0.00102766 3.3 0.00102758 3.3 0.00102768 0 0.0010275999999999998 0 0.0010276999999999999 3.3 0.00102762 3.3 0.00102772 0 0.00102764 0 0.00102774 3.3 0.00102766 3.3 0.00102776 0 0.00102768 0 0.00102778 3.3 0.0010276999999999999 3.3 0.0010278 0 0.00102772 0 0.00102782 3.3 0.0010277399999999999 3.3 0.00102784 0 0.00102776 0 0.00102786 3.3 0.0010277799999999998 3.3 0.00102788 0 0.0010278 0 0.0010279 3.3 0.0010278199999999998 3.3 0.0010279199999999999 0 0.00102784 0 0.00102794 3.3 0.00102786 3.3 0.00102796 0 0.00102788 0 0.00102798 3.3 0.0010279 3.3 0.001028 0 0.0010279199999999999 0 0.00102802 3.3 0.00102794 3.3 0.00102804 0 0.0010279599999999999 0 0.00102806 3.3 0.00102798 3.3 0.00102808 0 0.0010279999999999998 0 0.0010280999999999999 3.3 0.00102802 3.3 0.00102812 0 0.00102804 0 0.00102814 3.3 0.00102806 3.3 0.00102816 0 0.00102808 0 0.00102818 3.3 0.0010280999999999999 3.3 0.0010282 0 0.00102812 0 0.00102822 3.3 0.0010281399999999999 3.3 0.00102824 0 0.00102816 0 0.00102826 3.3 0.0010281799999999998 3.3 0.00102828 0 0.0010282 0 0.0010283 3.3 0.0010282199999999998 3.3 0.0010283199999999999 0 0.00102824 0 0.00102834 3.3 0.00102826 3.3 0.00102836 0 0.00102828 0 0.00102838 3.3 0.0010283 3.3 0.0010284 0 0.0010283199999999999 0 0.00102842 3.3 0.00102834 3.3 0.00102844 0 0.0010283599999999999 0 0.00102846 3.3 0.00102838 3.3 0.00102848 0 0.0010283999999999998 0 0.0010285 3.3 0.00102842 3.3 0.00102852 0 0.0010284399999999998 0 0.0010285399999999999 3.3 0.00102846 3.3 0.00102856 0 0.00102848 0 0.00102858 3.3 0.0010285 3.3 0.0010286 0 0.00102852 0 0.00102862 3.3 0.0010285399999999999 3.3 0.00102864 0 0.00102856 0 0.00102866 3.3 0.0010285799999999999 3.3 0.00102868 0 0.0010286 0 0.0010287 3.3 0.0010286199999999998 3.3 0.00102872 0 0.00102864 0 0.00102874 3.3 0.0010286599999999998 3.3 0.0010287599999999999 0 0.00102868 0 0.00102878 3.3 0.0010287 3.3 0.0010288 0 0.00102872 0 0.00102882 3.3 0.00102874 3.3 0.00102884 0 0.0010287599999999999 0 0.00102886 3.3 0.00102878 3.3 0.00102888 0 0.0010287999999999999 0 0.0010289 3.3 0.00102882 3.3 0.00102892 0 0.0010288399999999998 0 0.0010289399999999999 3.3 0.00102886 3.3 0.00102896 0 0.00102888 0 0.00102898 3.3 0.0010289 3.3 0.001029 0 0.00102892 0 0.00102902 3.3 0.0010289399999999999 3.3 0.00102904 0 0.00102896 0 0.00102906 3.3 0.0010289799999999999 3.3 0.00102908 0 0.001029 0 0.0010291 3.3 0.0010290199999999998 3.3 0.00102912 0 0.00102904 0 0.00102914 3.3 0.0010290599999999998 3.3 0.0010291599999999999 0 0.00102908 0 0.00102918 3.3 0.0010291 3.3 0.0010292 0 0.00102912 0 0.00102922 3.3 0.00102914 3.3 0.00102924 0 0.0010291599999999999 0 0.00102926 3.3 0.00102918 3.3 0.00102928 0 0.0010291999999999999 0 0.0010293 3.3 0.00102922 3.3 0.00102932 0 0.0010292399999999998 0 0.00102934 3.3 0.00102926 3.3 0.00102936 0 0.0010292799999999998 0 0.0010293799999999999 3.3 0.0010293 3.3 0.0010294 0 0.00102932 0 0.00102942 3.3 0.00102934 3.3 0.00102944 0 0.00102936 0 0.00102946 3.3 0.0010293799999999999 3.3 0.00102948 0 0.0010294 0 0.0010295 3.3 0.0010294199999999999 3.3 0.00102952 0 0.00102944 0 0.00102954 3.3 0.0010294599999999998 3.3 0.00102956 0 0.00102948 0 0.00102958 3.3 0.0010294999999999998 3.3 0.0010295999999999999 0 0.00102952 0 0.00102962 3.3 0.00102954 3.3 0.00102964 0 0.00102956 0 0.00102966 3.3 0.00102958 3.3 0.00102968 0 0.0010295999999999999 0 0.0010297 3.3 0.00102962 3.3 0.00102972 0 0.0010296399999999999 0 0.00102974 3.3 0.00102966 3.3 0.00102976 0 0.0010296799999999998 0 0.0010297799999999999 3.3 0.0010297 3.3 0.0010298 0 0.00102972 0 0.00102982 3.3 0.00102974 3.3 0.00102984 0 0.00102976 0 0.00102986 3.3 0.0010297799999999999 3.3 0.00102988 0 0.0010298 0 0.0010299 3.3 0.0010298199999999999 3.3 0.00102992 0 0.00102984 0 0.00102994 3.3 0.0010298599999999998 3.3 0.00102996 0 0.00102988 0 0.00102998 3.3 0.0010298999999999998 3.3 0.0010299999999999999 0 0.00102992 0 0.00103002 3.3 0.00102994 3.3 0.00103004 0 0.00102996 0 0.00103006 3.3 0.00102998 3.3 0.00103008 0 0.0010299999999999999 0 0.0010301 3.3 0.00103002 3.3 0.00103012 0 0.0010300399999999999 0 0.00103014 3.3 0.00103006 3.3 0.00103016 0 0.0010300799999999998 0 0.00103018 3.3 0.0010301 3.3 0.0010302 0 0.0010301199999999998 0 0.0010302199999999999 3.3 0.00103014 3.3 0.00103024 0 0.00103016 0 0.00103026 3.3 0.00103018 3.3 0.00103028 0 0.0010302 0 0.0010303 3.3 0.0010302199999999999 3.3 0.00103032 0 0.00103024 0 0.00103034 3.3 0.0010302599999999999 3.3 0.00103036 0 0.00103028 0 0.00103038 3.3 0.0010302999999999998 3.3 0.0010304 0 0.00103032 0 0.00103042 3.3 0.0010303399999999998 3.3 0.0010304399999999999 0 0.00103036 0 0.00103046 3.3 0.00103038 3.3 0.00103048 0 0.0010304 0 0.0010305 3.3 0.00103042 3.3 0.00103052 0 0.0010304399999999999 0 0.00103054 3.3 0.00103046 3.3 0.00103056 0 0.0010304799999999999 0 0.00103058 3.3 0.0010305 3.3 0.0010306 0 0.0010305199999999998 0 0.0010306199999999999 3.3 0.00103054 3.3 0.00103064 0 0.00103056 0 0.00103066 3.3 0.00103058 3.3 0.00103068 0 0.0010306 0 0.0010307 3.3 0.0010306199999999999 3.3 0.00103072 0 0.00103064 0 0.00103074 3.3 0.0010306599999999999 3.3 0.00103076 0 0.00103068 0 0.00103078 3.3 0.0010306999999999998 3.3 0.0010308 0 0.00103072 0 0.00103082 3.3 0.0010307399999999998 3.3 0.0010308399999999999 0 0.00103076 0 0.00103086 3.3 0.00103078 3.3 0.00103088 0 0.0010308 0 0.0010309 3.3 0.00103082 3.3 0.00103092 0 0.0010308399999999999 0 0.00103094 3.3 0.00103086 3.3 0.00103096 0 0.0010308799999999999 0 0.00103098 3.3 0.0010309 3.3 0.001031 0 0.0010309199999999998 0 0.00103102 3.3 0.00103094 3.3 0.00103104 0 0.0010309599999999998 0 0.0010310599999999999 3.3 0.00103098 3.3 0.00103108 0 0.001031 0 0.0010311 3.3 0.00103102 3.3 0.00103112 0 0.00103104 0 0.00103114 3.3 0.0010310599999999999 3.3 0.00103116 0 0.00103108 0 0.00103118 3.3 0.0010310999999999999 3.3 0.0010312 0 0.00103112 0 0.00103122 3.3 0.0010311399999999998 3.3 0.0010312399999999999 0 0.00103116 0 0.00103126 3.3 0.00103118 3.3 0.00103128 0 0.0010312 0 0.0010313 3.3 0.00103122 3.3 0.00103132 0 0.0010312399999999999 0 0.00103134 3.3 0.00103126 3.3 0.00103136 0 0.0010312799999999999 0 0.00103138 3.3 0.0010313 3.3 0.0010314 0 0.0010313199999999998 0 0.00103142 3.3 0.00103134 3.3 0.00103144 0 0.0010313599999999998 0 0.0010314599999999999 3.3 0.00103138 3.3 0.00103148 0 0.0010314 0 0.0010315 3.3 0.00103142 3.3 0.00103152 0 0.00103144 0 0.00103154 3.3 0.0010314599999999999 3.3 0.00103156 0 0.00103148 0 0.00103158 3.3 0.0010314999999999999 3.3 0.0010316 0 0.00103152 0 0.00103162 3.3 0.0010315399999999998 3.3 0.00103164 0 0.00103156 0 0.00103166 3.3 0.0010315799999999998 3.3 0.0010316799999999999 0 0.0010316 0 0.0010317 3.3 0.00103162 3.3 0.00103172 0 0.00103164 0 0.00103174 3.3 0.00103166 3.3 0.00103176 0 0.0010316799999999999 0 0.00103178 3.3 0.0010317 3.3 0.0010318 0 0.0010317199999999999 0 0.00103182 3.3 0.00103174 3.3 0.00103184 0 0.0010317599999999998 0 0.00103186 3.3 0.00103178 3.3 0.00103188 0 0.0010317999999999998 0 0.0010318999999999999 3.3 0.00103182 3.3 0.00103192 0 0.00103184 0 0.00103194 3.3 0.00103186 3.3 0.00103196 0 0.00103188 0 0.00103198 3.3 0.0010318999999999999 3.3 0.001032 0 0.00103192 0 0.00103202 3.3 0.0010319399999999999 3.3 0.00103204 0 0.00103196 0 0.00103206 3.3 0.0010319799999999998 3.3 0.0010320799999999999 0 0.001032 0 0.0010321 3.3 0.00103202 3.3 0.00103212 0 0.00103204 0 0.00103214 3.3 0.00103206 3.3 0.00103216 0 0.0010320799999999999 0 0.00103218 3.3 0.0010321 3.3 0.0010322 0 0.0010321199999999999 0 0.00103222 3.3 0.00103214 3.3 0.00103224 0 0.0010321599999999998 0 0.00103226 3.3 0.00103218 3.3 0.00103228 0 0.0010321999999999998 0 0.0010322999999999999 3.3 0.00103222 3.3 0.00103232 0 0.00103224 0 0.00103234 3.3 0.00103226 3.3 0.00103236 0 0.00103228 0 0.00103238 3.3 0.0010322999999999999 3.3 0.0010324 0 0.00103232 0 0.00103242 3.3 0.0010323399999999999 3.3 0.00103244 0 0.00103236 0 0.00103246 3.3 0.0010323799999999998 3.3 0.00103248 0 0.0010324 0 0.0010325 3.3 0.0010324199999999998 3.3 0.0010325199999999999 0 0.00103244 0 0.00103254 3.3 0.00103246 3.3 0.00103256 0 0.00103248 0 0.00103258 3.3 0.0010325 3.3 0.0010326 0 0.0010325199999999999 0 0.00103262 3.3 0.00103254 3.3 0.00103264 0 0.0010325599999999999 0 0.00103266 3.3 0.00103258 3.3 0.00103268 0 0.0010325999999999998 0 0.0010327 3.3 0.00103262 3.3 0.00103272 0 0.0010326399999999998 0 0.0010327399999999999 3.3 0.00103266 3.3 0.00103276 0 0.00103268 0 0.00103278 3.3 0.0010327 3.3 0.0010328 0 0.00103272 0 0.00103282 3.3 0.0010327399999999999 3.3 0.00103284 0 0.00103276 0 0.00103286 3.3 0.0010327799999999999 3.3 0.00103288 0 0.0010328 0 0.0010329 3.3 0.0010328199999999998 3.3 0.0010329199999999999 0 0.00103284 0 0.00103294 3.3 0.00103286 3.3 0.00103296 0 0.00103288 0 0.00103298 3.3 0.0010329 3.3 0.001033 0 0.0010329199999999999 0 0.00103302 3.3 0.00103294 3.3 0.00103304 0 0.0010329599999999999 0 0.00103306 3.3 0.00103298 3.3 0.00103308 0 0.0010329999999999998 0 0.0010331 3.3 0.00103302 3.3 0.00103312 0 0.0010330399999999998 0 0.0010331399999999999 3.3 0.00103306 3.3 0.00103316 0 0.00103308 0 0.00103318 3.3 0.0010331 3.3 0.0010332 0 0.00103312 0 0.00103322 3.3 0.0010331399999999999 3.3 0.00103324 0 0.00103316 0 0.00103326 3.3 0.0010331799999999999 3.3 0.00103328 0 0.0010332 0 0.0010333 3.3 0.0010332199999999998 3.3 0.00103332 0 0.00103324 0 0.00103334 3.3 0.0010332599999999998 3.3 0.0010333599999999999 0 0.00103328 0 0.00103338 3.3 0.0010333 3.3 0.0010334 0 0.00103332 0 0.00103342 3.3 0.00103334 3.3 0.00103344 0 0.0010333599999999999 0 0.00103346 3.3 0.00103338 3.3 0.00103348 0 0.0010333999999999999 0 0.0010335 3.3 0.00103342 3.3 0.00103352 0 0.0010334399999999998 0 0.00103354 3.3 0.00103346 3.3 0.00103356 0 0.0010334799999999998 0 0.0010335799999999999 3.3 0.0010335 3.3 0.0010336 0 0.00103352 0 0.00103362 3.3 0.00103354 3.3 0.00103364 0 0.00103356 0 0.00103366 3.3 0.0010335799999999999 3.3 0.00103368 0 0.0010336 0 0.0010337 3.3 0.0010336199999999999 3.3 0.00103372 0 0.00103364 0 0.00103374 3.3 0.0010336599999999998 3.3 0.0010337599999999999 0 0.00103368 0 0.00103378 3.3 0.0010337 3.3 0.0010338 0 0.00103372 0 0.00103382 3.3 0.00103374 3.3 0.00103384 0 0.0010337599999999999 0 0.00103386 3.3 0.00103378 3.3 0.00103388 0 0.0010337999999999999 0 0.0010339 3.3 0.00103382 3.3 0.00103392 0 0.0010338399999999998 0 0.00103394 3.3 0.00103386 3.3 0.00103396 0 0.0010338799999999998 0 0.0010339799999999999 3.3 0.0010339 3.3 0.001034 0 0.00103392 0 0.00103402 3.3 0.00103394 3.3 0.00103404 0 0.00103396 0 0.00103406 3.3 0.0010339799999999999 3.3 0.00103408 0 0.001034 0 0.0010341 3.3 0.0010340199999999999 3.3 0.00103412 0 0.00103404 0 0.00103414 3.3 0.0010340599999999998 3.3 0.00103416 0 0.00103408 0 0.00103418 3.3 0.0010340999999999998 3.3 0.0010341999999999999 0 0.00103412 0 0.00103422 3.3 0.00103414 3.3 0.00103424 0 0.00103416 0 0.00103426 3.3 0.00103418 3.3 0.00103428 0 0.0010341999999999999 0 0.0010343 3.3 0.00103422 3.3 0.00103432 0 0.0010342399999999999 0 0.00103434 3.3 0.00103426 3.3 0.00103436 0 0.0010342799999999998 0 0.0010343799999999999 3.3 0.0010343 3.3 0.0010344 0 0.0010343199999999998 0 0.0010344199999999999 3.3 0.00103434 3.3 0.00103444 0 0.00103436 0 0.00103446 3.3 0.0010343799999999999 3.3 0.00103448 0 0.0010344 0 0.0010345 3.3 0.0010344199999999999 3.3 0.00103452 0 0.00103444 0 0.00103454 3.3 0.0010344599999999999 3.3 0.00103456 0 0.00103448 0 0.00103458 3.3 0.0010344999999999998 3.3 0.0010345999999999999 0 0.00103452 0 0.00103462 3.3 0.00103454 3.3 0.00103464 0 0.00103456 0 0.00103466 3.3 0.00103458 3.3 0.00103468 0 0.0010345999999999999 0 0.0010347 3.3 0.00103462 3.3 0.00103472 0 0.0010346399999999999 0 0.00103474 3.3 0.00103466 3.3 0.00103476 0 0.0010346799999999998 0 0.00103478 3.3 0.0010347 3.3 0.0010348 0 0.0010347199999999998 0 0.0010348199999999999 3.3 0.00103474 3.3 0.00103484 0 0.00103476 0 0.00103486 3.3 0.00103478 3.3 0.00103488 0 0.0010348 0 0.0010349 3.3 0.0010348199999999999 3.3 0.00103492 0 0.00103484 0 0.00103494 3.3 0.0010348599999999999 3.3 0.00103496 0 0.00103488 0 0.00103498 3.3 0.0010348999999999998 3.3 0.001035 0 0.00103492 0 0.00103502 3.3 0.0010349399999999998 3.3 0.0010350399999999999 0 0.00103496 0 0.00103506 3.3 0.00103498 3.3 0.00103508 0 0.001035 0 0.0010351 3.3 0.00103502 3.3 0.00103512 0 0.0010350399999999999 0 0.00103514 3.3 0.00103506 3.3 0.00103516 0 0.0010350799999999999 0 0.00103518 3.3 0.0010351 3.3 0.0010352 0 0.0010351199999999998 0 0.0010352199999999999 3.3 0.00103514 3.3 0.00103524 0 0.00103516 0 0.00103526 3.3 0.00103518 3.3 0.00103528 0 0.0010352 0 0.0010353 3.3 0.0010352199999999999 3.3 0.00103532 0 0.00103524 0 0.00103534 3.3 0.0010352599999999999 3.3 0.00103536 0 0.00103528 0 0.00103538 3.3 0.0010352999999999998 3.3 0.0010354 0 0.00103532 0 0.00103542 3.3 0.0010353399999999998 3.3 0.0010354399999999999 0 0.00103536 0 0.00103546 3.3 0.00103538 3.3 0.00103548 0 0.0010354 0 0.0010355 3.3 0.00103542 3.3 0.00103552 0 0.0010354399999999999 0 0.00103554 3.3 0.00103546 3.3 0.00103556 0 0.0010354799999999999 0 0.00103558 3.3 0.0010355 3.3 0.0010356 0 0.0010355199999999998 0 0.00103562 3.3 0.00103554 3.3 0.00103564 0 0.0010355599999999998 0 0.0010356599999999999 3.3 0.00103558 3.3 0.00103568 0 0.0010356 0 0.0010357 3.3 0.00103562 3.3 0.00103572 0 0.00103564 0 0.00103574 3.3 0.0010356599999999999 3.3 0.00103576 0 0.00103568 0 0.00103578 3.3 0.0010356999999999999 3.3 0.0010358 0 0.00103572 0 0.00103582 3.3 0.0010357399999999998 3.3 0.00103584 0 0.00103576 0 0.00103586 3.3 0.0010357799999999998 3.3 0.0010358799999999999 0 0.0010358 0 0.0010359 3.3 0.00103582 3.3 0.00103592 0 0.00103584 0 0.00103594 3.3 0.00103586 3.3 0.00103596 0 0.0010358799999999999 0 0.00103598 3.3 0.0010359 3.3 0.001036 0 0.0010359199999999999 0 0.00103602 3.3 0.00103594 3.3 0.00103604 0 0.0010359599999999998 0 0.0010360599999999999 3.3 0.00103598 3.3 0.00103608 0 0.001036 0 0.0010361 3.3 0.00103602 3.3 0.00103612 0 0.00103604 0 0.00103614 3.3 0.0010360599999999999 3.3 0.00103616 0 0.00103608 0 0.00103618 3.3 0.0010360999999999999 3.3 0.0010362 0 0.00103612 0 0.00103622 3.3 0.0010361399999999998 3.3 0.00103624 0 0.00103616 0 0.00103626 3.3 0.0010361799999999998 3.3 0.0010362799999999999 0 0.0010362 0 0.0010363 3.3 0.00103622 3.3 0.00103632 0 0.00103624 0 0.00103634 3.3 0.00103626 3.3 0.00103636 0 0.0010362799999999999 0 0.00103638 3.3 0.0010363 3.3 0.0010364 0 0.0010363199999999999 0 0.00103642 3.3 0.00103634 3.3 0.00103644 0 0.0010363599999999998 0 0.00103646 3.3 0.00103638 3.3 0.00103648 0 0.0010363999999999998 0 0.0010364999999999999 3.3 0.00103642 3.3 0.00103652 0 0.00103644 0 0.00103654 3.3 0.00103646 3.3 0.00103656 0 0.00103648 0 0.00103658 3.3 0.0010364999999999999 3.3 0.0010366 0 0.00103652 0 0.00103662 3.3 0.0010365399999999999 3.3 0.00103664 0 0.00103656 0 0.00103666 3.3 0.0010365799999999998 3.3 0.00103668 0 0.0010366 0 0.0010367 3.3 0.0010366199999999998 3.3 0.0010367199999999999 0 0.00103664 0 0.00103674 3.3 0.00103666 3.3 0.00103676 0 0.00103668 0 0.00103678 3.3 0.0010367 3.3 0.0010368 0 0.0010367199999999999 0 0.00103682 3.3 0.00103674 3.3 0.00103684 0 0.0010367599999999999 0 0.00103686 3.3 0.00103678 3.3 0.00103688 0 0.0010367999999999998 0 0.0010368999999999999 3.3 0.00103682 3.3 0.00103692 0 0.00103684 0 0.00103694 3.3 0.00103686 3.3 0.00103696 0 0.00103688 0 0.00103698 3.3 0.0010368999999999999 3.3 0.001037 0 0.00103692 0 0.00103702 3.3 0.0010369399999999999 3.3 0.00103704 0 0.00103696 0 0.00103706 3.3 0.0010369799999999998 3.3 0.00103708 0 0.001037 0 0.0010371 3.3 0.0010370199999999998 3.3 0.0010371199999999999 0 0.00103704 0 0.00103714 3.3 0.00103706 3.3 0.00103716 0 0.00103708 0 0.00103718 3.3 0.0010371 3.3 0.0010372 0 0.0010371199999999999 0 0.00103722 3.3 0.00103714 3.3 0.00103724 0 0.0010371599999999999 0 0.00103726 3.3 0.00103718 3.3 0.00103728 0 0.0010371999999999998 0 0.0010373 3.3 0.00103722 3.3 0.00103732 0 0.0010372399999999998 0 0.0010373399999999999 3.3 0.00103726 3.3 0.00103736 0 0.00103728 0 0.00103738 3.3 0.0010373 3.3 0.0010374 0 0.00103732 0 0.00103742 3.3 0.0010373399999999999 3.3 0.00103744 0 0.00103736 0 0.00103746 3.3 0.0010373799999999999 3.3 0.00103748 0 0.0010374 0 0.0010375 3.3 0.0010374199999999998 3.3 0.00103752 0 0.00103744 0 0.00103754 3.3 0.0010374599999999998 3.3 0.0010375599999999999 0 0.00103748 0 0.00103758 3.3 0.0010375 3.3 0.0010376 0 0.00103752 0 0.00103762 3.3 0.00103754 3.3 0.00103764 0 0.0010375599999999999 0 0.00103766 3.3 0.00103758 3.3 0.00103768 0 0.0010375999999999999 0 0.0010377 3.3 0.00103762 3.3 0.00103772 0 0.0010376399999999998 0 0.0010377399999999999 3.3 0.00103766 3.3 0.00103776 0 0.00103768 0 0.00103778 3.3 0.0010377 3.3 0.0010378 0 0.00103772 0 0.00103782 3.3 0.0010377399999999999 3.3 0.00103784 0 0.00103776 0 0.00103786 3.3 0.0010377799999999999 3.3 0.00103788 0 0.0010378 0 0.0010379 3.3 0.0010378199999999998 3.3 0.00103792 0 0.00103784 0 0.00103794 3.3 0.0010378599999999998 3.3 0.0010379599999999999 0 0.00103788 0 0.00103798 3.3 0.0010379 3.3 0.001038 0 0.00103792 0 0.00103802 3.3 0.00103794 3.3 0.00103804 0 0.0010379599999999999 0 0.00103806 3.3 0.00103798 3.3 0.00103808 0 0.0010379999999999999 0 0.0010381 3.3 0.00103802 3.3 0.00103812 0 0.0010380399999999998 0 0.00103814 3.3 0.00103806 3.3 0.00103816 0 0.0010380799999999998 0 0.0010381799999999999 3.3 0.0010381 3.3 0.0010382 0 0.00103812 0 0.00103822 3.3 0.00103814 3.3 0.00103824 0 0.00103816 0 0.00103826 3.3 0.0010381799999999999 3.3 0.00103828 0 0.0010382 0 0.0010383 3.3 0.0010382199999999999 3.3 0.00103832 0 0.00103824 0 0.00103834 3.3 0.0010382599999999998 3.3 0.0010383599999999999 0 0.00103828 0 0.00103838 3.3 0.0010383 3.3 0.0010384 0 0.00103832 0 0.00103842 3.3 0.00103834 3.3 0.00103844 0 0.0010383599999999999 0 0.00103846 3.3 0.00103838 3.3 0.00103848 0 0.0010383999999999999 0 0.0010385 3.3 0.00103842 3.3 0.00103852 0 0.0010384399999999998 0 0.00103854 3.3 0.00103846 3.3 0.00103856 0 0.0010384799999999998 0 0.0010385799999999999 3.3 0.0010385 3.3 0.0010386 0 0.00103852 0 0.00103862 3.3 0.00103854 3.3 0.00103864 0 0.00103856 0 0.00103866 3.3 0.0010385799999999999 3.3 0.00103868 0 0.0010386 0 0.0010387 3.3 0.0010386199999999999 3.3 0.00103872 0 0.00103864 0 0.00103874 3.3 0.0010386599999999998 3.3 0.00103876 0 0.00103868 0 0.00103878 3.3 0.0010386999999999998 3.3 0.0010387999999999999 0 0.00103872 0 0.00103882 3.3 0.00103874 3.3 0.00103884 0 0.00103876 0 0.00103886 3.3 0.00103878 3.3 0.00103888 0 0.0010387999999999999 0 0.0010389 3.3 0.00103882 3.3 0.00103892 0 0.0010388399999999999 0 0.00103894 3.3 0.00103886 3.3 0.00103896 0 0.0010388799999999998 0 0.00103898 3.3 0.0010389 3.3 0.001039 0 0.0010389199999999998 0 0.0010390199999999999 3.3 0.00103894 3.3 0.00103904 0 0.00103896 0 0.00103906 3.3 0.00103898 3.3 0.00103908 0 0.001039 0 0.0010391 3.3 0.0010390199999999999 3.3 0.00103912 0 0.00103904 0 0.00103914 3.3 0.0010390599999999999 3.3 0.00103916 0 0.00103908 0 0.00103918 3.3 0.0010390999999999998 3.3 0.0010391999999999999 0 0.00103912 0 0.00103922 3.3 0.00103914 3.3 0.00103924 0 0.00103916 0 0.00103926 3.3 0.00103918 3.3 0.00103928 0 0.0010391999999999999 0 0.0010393 3.3 0.00103922 3.3 0.00103932 0 0.0010392399999999999 0 0.00103934 3.3 0.00103926 3.3 0.00103936 0 0.0010392799999999998 0 0.00103938 3.3 0.0010393 3.3 0.0010394 0 0.0010393199999999998 0 0.0010394199999999999 3.3 0.00103934 3.3 0.00103944 0 0.00103936 0 0.00103946 3.3 0.00103938 3.3 0.00103948 0 0.0010394 0 0.0010395 3.3 0.0010394199999999999 3.3 0.00103952 0 0.00103944 0 0.00103954 3.3 0.0010394599999999999 3.3 0.00103956 0 0.00103948 0 0.00103958 3.3 0.0010394999999999998 3.3 0.0010396 0 0.00103952 0 0.00103962 3.3 0.0010395399999999998 3.3 0.0010396399999999999 0 0.00103956 0 0.00103966 3.3 0.00103958 3.3 0.00103968 0 0.0010396 0 0.0010397 3.3 0.00103962 3.3 0.00103972 0 0.0010396399999999999 0 0.00103974 3.3 0.00103966 3.3 0.00103976 0 0.0010396799999999999 0 0.00103978 3.3 0.0010397 3.3 0.0010398 0 0.0010397199999999998 0 0.00103982 3.3 0.00103974 3.3 0.00103984 0 0.0010397599999999998 0 0.0010398599999999999 3.3 0.00103978 3.3 0.00103988 0 0.0010398 0 0.0010399 3.3 0.00103982 3.3 0.00103992 0 0.00103984 0 0.00103994 3.3 0.0010398599999999999 3.3 0.00103996 0 0.00103988 0 0.00103998 3.3 0.0010398999999999999 3.3 0.00104 0 0.00103992 0 0.00104002 3.3 0.0010399399999999998 3.3 0.0010400399999999999 0 0.00103996 0 0.00104006 3.3 0.00103998 3.3 0.00104008 0 0.00104 0 0.0010401 3.3 0.00104002 3.3 0.00104012 0 0.0010400399999999999 0 0.00104014 3.3 0.00104006 3.3 0.00104016 0 0.0010400799999999999 0 0.00104018 3.3 0.0010401 3.3 0.0010402 0 0.0010401199999999998 0 0.00104022 3.3 0.00104014 3.3 0.00104024 0 0.0010401599999999998 0 0.0010402599999999999 3.3 0.00104018 3.3 0.00104028 0 0.0010402 0 0.0010403 3.3 0.00104022 3.3 0.00104032 0 0.00104024 0 0.00104034 3.3 0.0010402599999999999 3.3 0.00104036 0 0.00104028 0 0.00104038 3.3 0.0010402999999999999 3.3 0.0010404 0 0.00104032 0 0.00104042 3.3 0.0010403399999999998 3.3 0.00104044 0 0.00104036 0 0.00104046 3.3 0.0010403799999999998 3.3 0.0010404799999999999 0 0.0010404 0 0.0010405 3.3 0.00104042 3.3 0.00104052 0 0.00104044 0 0.00104054 3.3 0.00104046 3.3 0.00104056 0 0.0010404799999999999 0 0.00104058 3.3 0.0010405 3.3 0.0010406 0 0.0010405199999999999 0 0.00104062 3.3 0.00104054 3.3 0.00104064 0 0.0010405599999999998 0 0.00104066 3.3 0.00104058 3.3 0.00104068 0 0.0010405999999999998 0 0.0010406999999999999 3.3 0.00104062 3.3 0.00104072 0 0.00104064 0 0.00104074 3.3 0.00104066 3.3 0.00104076 0 0.00104068 0 0.00104078 3.3 0.0010406999999999999 3.3 0.0010408 0 0.00104072 0 0.00104082 3.3 0.0010407399999999999 3.3 0.00104084 0 0.00104076 0 0.00104086 3.3 0.0010407799999999998 3.3 0.0010408799999999999 0 0.0010408 0 0.0010409 3.3 0.00104082 3.3 0.00104092 0 0.00104084 0 0.00104094 3.3 0.00104086 3.3 0.00104096 0 0.0010408799999999999 0 0.00104098 3.3 0.0010409 3.3 0.001041 0 0.0010409199999999999 0 0.00104102 3.3 0.00104094 3.3 0.00104104 0 0.0010409599999999998 0 0.00104106 3.3 0.00104098 3.3 0.00104108 0 0.0010409999999999998 0 0.0010410999999999999 3.3 0.00104102 3.3 0.00104112 0 0.00104104 0 0.00104114 3.3 0.00104106 3.3 0.00104116 0 0.00104108 0 0.00104118 3.3 0.0010410999999999999 3.3 0.0010412 0 0.00104112 0 0.00104122 3.3 0.0010411399999999999 3.3 0.00104124 0 0.00104116 0 0.00104126 3.3 0.0010411799999999998 3.3 0.00104128 0 0.0010412 0 0.0010413 3.3 0.0010412199999999998 3.3 0.0010413199999999999 0 0.00104124 0 0.00104134 3.3 0.00104126 3.3 0.00104136 0 0.00104128 0 0.00104138 3.3 0.0010413 3.3 0.0010414 0 0.0010413199999999999 0 0.00104142 3.3 0.00104134 3.3 0.00104144 0 0.0010413599999999999 0 0.00104146 3.3 0.00104138 3.3 0.00104148 0 0.0010413999999999998 0 0.0010414999999999999 3.3 0.00104142 3.3 0.00104152 0 0.00104144 0 0.00104154 3.3 0.00104146 3.3 0.00104156 0 0.00104148 0 0.00104158 3.3 0.0010414999999999999 3.3 0.0010416 0 0.00104152 0 0.00104162 3.3 0.0010415399999999999 3.3 0.00104164 0 0.00104156 0 0.00104166 3.3 0.0010415799999999998 3.3 0.00104168 0 0.0010416 0 0.0010417 3.3 0.0010416199999999998 3.3 0.0010417199999999999 0 0.00104164 0 0.00104174 3.3 0.00104166 3.3 0.00104176 0 0.00104168 0 0.00104178 3.3 0.0010417 3.3 0.0010418 0 0.0010417199999999999 0 0.00104182 3.3 0.00104174 3.3 0.00104184 0 0.0010417599999999999 0 0.00104186 3.3 0.00104178 3.3 0.00104188 0 0.0010417999999999998 0 0.0010419 3.3 0.00104182 3.3 0.00104192 0 0.0010418399999999998 0 0.0010419399999999999 3.3 0.00104186 3.3 0.00104196 0 0.00104188 0 0.00104198 3.3 0.0010419 3.3 0.001042 0 0.00104192 0 0.00104202 3.3 0.0010419399999999999 3.3 0.00104204 0 0.00104196 0 0.00104206 3.3 0.0010419799999999999 3.3 0.00104208 0 0.001042 0 0.0010421 3.3 0.0010420199999999998 3.3 0.00104212 0 0.00104204 0 0.00104214 3.3 0.0010420599999999998 3.3 0.0010421599999999999 0 0.00104208 0 0.00104218 3.3 0.0010421 3.3 0.0010422 0 0.00104212 0 0.00104222 3.3 0.00104214 3.3 0.00104224 0 0.0010421599999999999 0 0.00104226 3.3 0.00104218 3.3 0.00104228 0 0.0010421999999999999 0 0.0010423 3.3 0.00104222 3.3 0.00104232 0 0.0010422399999999998 0 0.0010423399999999999 3.3 0.00104226 3.3 0.00104236 0 0.00104228 0 0.00104238 3.3 0.0010423 3.3 0.0010424 0 0.00104232 0 0.00104242 3.3 0.0010423399999999999 3.3 0.00104244 0 0.00104236 0 0.00104246 3.3 0.0010423799999999999 3.3 0.00104248 0 0.0010424 0 0.0010425 3.3 0.0010424199999999998 3.3 0.00104252 0 0.00104244 0 0.00104254 3.3 0.0010424599999999998 3.3 0.0010425599999999999 0 0.00104248 0 0.00104258 3.3 0.0010425 3.3 0.0010426 0 0.00104252 0 0.00104262 3.3 0.00104254 3.3 0.00104264 0 0.0010425599999999999 0 0.00104266 3.3 0.00104258 3.3 0.00104268 0 0.0010425999999999999 0 0.0010427 3.3 0.00104262 3.3 0.00104272 0 0.0010426399999999998 0 0.00104274 3.3 0.00104266 3.3 0.00104276 0 0.0010426799999999998 0 0.0010427799999999999 3.3 0.0010427 3.3 0.0010428 0 0.00104272 0 0.00104282 3.3 0.00104274 3.3 0.00104284 0 0.00104276 0 0.00104286 3.3 0.0010427799999999999 3.3 0.00104288 0 0.0010428 0 0.0010429 3.3 0.0010428199999999999 3.3 0.00104292 0 0.00104284 0 0.00104294 3.3 0.0010428599999999998 3.3 0.00104296 0 0.00104288 0 0.00104298 3.3 0.0010428999999999998 3.3 0.0010429999999999999 0 0.00104292 0 0.00104302 3.3 0.00104294 3.3 0.00104304 0 0.00104296 0 0.00104306 3.3 0.00104298 3.3 0.00104308 0 0.0010429999999999999 0 0.0010431 3.3 0.00104302 3.3 0.00104312 0 0.0010430399999999999 0 0.00104314 3.3 0.00104306 3.3 0.00104316 0 0.0010430799999999998 0 0.0010431799999999999 3.3 0.0010431 3.3 0.0010432 0 0.00104312 0 0.00104322 3.3 0.00104314 3.3 0.00104324 0 0.00104316 0 0.00104326 3.3 0.0010431799999999999 3.3 0.00104328 0 0.0010432 0 0.0010433 3.3 0.0010432199999999999 3.3 0.00104332 0 0.00104324 0 0.00104334 3.3 0.0010432599999999998 3.3 0.00104336 0 0.00104328 0 0.00104338 3.3 0.0010432999999999998 3.3 0.0010433999999999999 0 0.00104332 0 0.00104342 3.3 0.00104334 3.3 0.00104344 0 0.00104336 0 0.00104346 3.3 0.00104338 3.3 0.00104348 0 0.0010433999999999999 0 0.0010435 3.3 0.00104342 3.3 0.00104352 0 0.0010434399999999999 0 0.00104354 3.3 0.00104346 3.3 0.00104356 0 0.0010434799999999998 0 0.00104358 3.3 0.0010435 3.3 0.0010436 0 0.0010435199999999998 0 0.0010436199999999999 3.3 0.00104354 3.3 0.00104364 0 0.00104356 0 0.00104366 3.3 0.00104358 3.3 0.00104368 0 0.0010436 0 0.0010437 3.3 0.0010436199999999999 3.3 0.00104372 0 0.00104364 0 0.00104374 3.3 0.0010436599999999999 3.3 0.00104376 0 0.00104368 0 0.00104378 3.3 0.0010436999999999998 3.3 0.0010438 0 0.00104372 0 0.00104382 3.3 0.0010437399999999998 3.3 0.0010438399999999999 0 0.00104376 0 0.00104386 3.3 0.00104378 3.3 0.00104388 0 0.0010438 0 0.0010439 3.3 0.00104382 3.3 0.00104392 0 0.0010438399999999999 0 0.00104394 3.3 0.00104386 3.3 0.00104396 0 0.0010438799999999999 0 0.00104398 3.3 0.0010439 3.3 0.001044 0 0.0010439199999999998 0 0.0010440199999999999 3.3 0.00104394 3.3 0.00104404 0 0.00104396 0 0.00104406 3.3 0.00104398 3.3 0.00104408 0 0.001044 0 0.0010441 3.3 0.0010440199999999999 3.3 0.00104412 0 0.00104404 0 0.00104414 3.3 0.0010440599999999999 3.3 0.00104416 0 0.00104408 0 0.00104418 3.3 0.0010440999999999998 3.3 0.0010442 0 0.00104412 0 0.00104422 3.3 0.0010441399999999998 3.3 0.0010442399999999999 0 0.00104416 0 0.00104426 3.3 0.00104418 3.3 0.00104428 0 0.0010442 0 0.0010443 3.3 0.00104422 3.3 0.00104432 0 0.0010442399999999999 0 0.00104434 3.3 0.00104426 3.3 0.00104436 0 0.0010442799999999999 0 0.00104438 3.3 0.0010443 3.3 0.0010444 0 0.0010443199999999998 0 0.00104442 3.3 0.00104434 3.3 0.00104444 0 0.0010443599999999998 0 0.0010444599999999999 3.3 0.00104438 3.3 0.00104448 0 0.0010444 0 0.0010445 3.3 0.00104442 3.3 0.00104452 0 0.00104444 0 0.00104454 3.3 0.0010444599999999999 3.3 0.00104456 0 0.00104448 0 0.00104458 3.3 0.0010444999999999999 3.3 0.0010446 0 0.00104452 0 0.00104462 3.3 0.0010445399999999998 3.3 0.0010446399999999999 0 0.00104456 0 0.00104466 3.3 0.0010445799999999998 3.3 0.0010446799999999999 0 0.0010446 0 0.0010447 3.3 0.00104462 3.3 0.00104472 0 0.0010446399999999999 0 0.00104474 3.3 0.00104466 3.3 0.00104476 0 0.0010446799999999999 0 0.00104478 3.3 0.0010447 3.3 0.0010448 0 0.0010447199999999999 0 0.00104482 3.3 0.00104474 3.3 0.00104484 0 0.0010447599999999998 0 0.0010448599999999999 3.3 0.00104478 3.3 0.00104488 0 0.0010448 0 0.0010449 3.3 0.00104482 3.3 0.00104492 0 0.00104484 0 0.00104494 3.3 0.0010448599999999999 3.3 0.00104496 0 0.00104488 0 0.00104498 3.3 0.0010448999999999999 3.3 0.001045 0 0.00104492 0 0.00104502 3.3 0.0010449399999999998 3.3 0.00104504 0 0.00104496 0 0.00104506 3.3 0.0010449799999999998 3.3 0.0010450799999999999 0 0.001045 0 0.0010451 3.3 0.00104502 3.3 0.00104512 0 0.00104504 0 0.00104514 3.3 0.00104506 3.3 0.00104516 0 0.0010450799999999999 0 0.00104518 3.3 0.0010451 3.3 0.0010452 0 0.0010451199999999999 0 0.00104522 3.3 0.00104514 3.3 0.00104524 0 0.0010451599999999998 0 0.00104526 3.3 0.00104518 3.3 0.00104528 0 0.0010451999999999998 0 0.0010452999999999999 3.3 0.00104522 3.3 0.00104532 0 0.00104524 0 0.00104534 3.3 0.00104526 3.3 0.00104536 0 0.00104528 0 0.00104538 3.3 0.0010452999999999999 3.3 0.0010454 0 0.00104532 0 0.00104542 3.3 0.0010453399999999999 3.3 0.00104544 0 0.00104536 0 0.00104546 3.3 0.0010453799999999998 3.3 0.0010454799999999999 0 0.0010454 0 0.0010455 3.3 0.00104542 3.3 0.00104552 0 0.00104544 0 0.00104554 3.3 0.00104546 3.3 0.00104556 0 0.0010454799999999999 0 0.00104558 3.3 0.0010455 3.3 0.0010456 0 0.0010455199999999999 0 0.00104562 3.3 0.00104554 3.3 0.00104564 0 0.0010455599999999998 0 0.00104566 3.3 0.00104558 3.3 0.00104568 0 0.0010455999999999998 0 0.0010456999999999999 3.3 0.00104562 3.3 0.00104572 0 0.00104564 0 0.00104574 3.3 0.00104566 3.3 0.00104576 0 0.00104568 0 0.00104578 3.3 0.0010456999999999999 3.3 0.0010458 0 0.00104572 0 0.00104582 3.3 0.0010457399999999999 3.3 0.00104584 0 0.00104576 0 0.00104586 3.3 0.0010457799999999998 3.3 0.00104588 0 0.0010458 0 0.0010459 3.3 0.0010458199999999998 3.3 0.0010459199999999999 0 0.00104584 0 0.00104594 3.3 0.00104586 3.3 0.00104596 0 0.00104588 0 0.00104598 3.3 0.0010459 3.3 0.001046 0 0.0010459199999999999 0 0.00104602 3.3 0.00104594 3.3 0.00104604 0 0.0010459599999999999 0 0.00104606 3.3 0.00104598 3.3 0.00104608 0 0.0010459999999999998 0 0.0010461 3.3 0.00104602 3.3 0.00104612 0 0.0010460399999999998 0 0.0010461399999999999 3.3 0.00104606 3.3 0.00104616 0 0.00104608 0 0.00104618 3.3 0.0010461 3.3 0.0010462 0 0.00104612 0 0.00104622 3.3 0.0010461399999999999 3.3 0.00104624 0 0.00104616 0 0.00104626 3.3 0.0010461799999999999 3.3 0.00104628 0 0.0010462 0 0.0010463 3.3 0.0010462199999999998 3.3 0.0010463199999999999 0 0.00104624 0 0.00104634 3.3 0.00104626 3.3 0.00104636 0 0.00104628 0 0.00104638 3.3 0.0010463 3.3 0.0010464 0 0.0010463199999999999 0 0.00104642 3.3 0.00104634 3.3 0.00104644 0 0.0010463599999999999 0 0.00104646 3.3 0.00104638 3.3 0.00104648 0 0.0010463999999999998 0 0.0010465 3.3 0.00104642 3.3 0.00104652 0 0.0010464399999999998 0 0.0010465399999999999 3.3 0.00104646 3.3 0.00104656 0 0.00104648 0 0.00104658 3.3 0.0010465 3.3 0.0010466 0 0.00104652 0 0.00104662 3.3 0.0010465399999999999 3.3 0.00104664 0 0.00104656 0 0.00104666 3.3 0.0010465799999999999 3.3 0.00104668 0 0.0010466 0 0.0010467 3.3 0.0010466199999999998 3.3 0.00104672 0 0.00104664 0 0.00104674 3.3 0.0010466599999999998 3.3 0.0010467599999999999 0 0.00104668 0 0.00104678 3.3 0.0010467 3.3 0.0010468 0 0.00104672 0 0.00104682 3.3 0.00104674 3.3 0.00104684 0 0.0010467599999999999 0 0.00104686 3.3 0.00104678 3.3 0.00104688 0 0.0010467999999999999 0 0.0010469 3.3 0.00104682 3.3 0.00104692 0 0.0010468399999999998 0 0.00104694 3.3 0.00104686 3.3 0.00104696 0 0.0010468799999999998 0 0.0010469799999999999 3.3 0.0010469 3.3 0.001047 0 0.00104692 0 0.00104702 3.3 0.00104694 3.3 0.00104704 0 0.00104696 0 0.00104706 3.3 0.0010469799999999999 3.3 0.00104708 0 0.001047 0 0.0010471 3.3 0.0010470199999999999 3.3 0.00104712 0 0.00104704 0 0.00104714 3.3 0.0010470599999999998 3.3 0.0010471599999999999 0 0.00104708 0 0.00104718 3.3 0.0010471 3.3 0.0010472 0 0.00104712 0 0.00104722 3.3 0.00104714 3.3 0.00104724 0 0.0010471599999999999 0 0.00104726 3.3 0.00104718 3.3 0.00104728 0 0.0010471999999999999 0 0.0010473 3.3 0.00104722 3.3 0.00104732 0 0.0010472399999999998 0 0.00104734 3.3 0.00104726 3.3 0.00104736 0 0.0010472799999999998 0 0.0010473799999999999 3.3 0.0010473 3.3 0.0010474 0 0.00104732 0 0.00104742 3.3 0.00104734 3.3 0.00104744 0 0.00104736 0 0.00104746 3.3 0.0010473799999999999 3.3 0.00104748 0 0.0010474 0 0.0010475 3.3 0.0010474199999999999 3.3 0.00104752 0 0.00104744 0 0.00104754 3.3 0.0010474599999999998 3.3 0.00104756 0 0.00104748 0 0.00104758 3.3 0.0010474999999999998 3.3 0.0010475999999999999 0 0.00104752 0 0.00104762 3.3 0.00104754 3.3 0.00104764 0 0.00104756 0 0.00104766 3.3 0.00104758 3.3 0.00104768 0 0.0010475999999999999 0 0.0010477 3.3 0.00104762 3.3 0.00104772 0 0.0010476399999999999 0 0.00104774 3.3 0.00104766 3.3 0.00104776 0 0.0010476799999999998 0 0.00104778 3.3 0.0010477 3.3 0.0010478 0 0.0010477199999999998 0 0.0010478199999999999 3.3 0.00104774 3.3 0.00104784 0 0.00104776 0 0.00104786 3.3 0.00104778 3.3 0.00104788 0 0.0010478 0 0.0010479 3.3 0.0010478199999999999 3.3 0.00104792 0 0.00104784 0 0.00104794 3.3 0.0010478599999999999 3.3 0.00104796 0 0.00104788 0 0.00104798 3.3 0.0010478999999999998 3.3 0.0010479999999999999 0 0.00104792 0 0.00104802 3.3 0.00104794 3.3 0.00104804 0 0.00104796 0 0.00104806 3.3 0.00104798 3.3 0.00104808 0 0.0010479999999999999 0 0.0010481 3.3 0.00104802 3.3 0.00104812 0 0.0010480399999999999 0 0.00104814 3.3 0.00104806 3.3 0.00104816 0 0.0010480799999999998 0 0.00104818 3.3 0.0010481 3.3 0.0010482 0 0.0010481199999999998 0 0.0010482199999999999 3.3 0.00104814 3.3 0.00104824 0 0.00104816 0 0.00104826 3.3 0.00104818 3.3 0.00104828 0 0.0010482 0 0.0010483 3.3 0.0010482199999999999 3.3 0.00104832 0 0.00104824 0 0.00104834 3.3 0.0010482599999999999 3.3 0.00104836 0 0.00104828 0 0.00104838 3.3 0.0010482999999999998 3.3 0.0010484 0 0.00104832 0 0.00104842 3.3 0.0010483399999999998 3.3 0.0010484399999999999 0 0.00104836 0 0.00104846 3.3 0.00104838 3.3 0.00104848 0 0.0010484 0 0.0010485 3.3 0.00104842 3.3 0.00104852 0 0.0010484399999999999 0 0.00104854 3.3 0.00104846 3.3 0.00104856 0 0.0010484799999999999 0 0.00104858 3.3 0.0010485 3.3 0.0010486 0 0.0010485199999999998 0 0.0010486199999999999 3.3 0.00104854 3.3 0.00104864 0 0.00104856 0 0.00104866 3.3 0.00104858 3.3 0.00104868 0 0.0010486 0 0.0010487 3.3 0.0010486199999999999 3.3 0.00104872 0 0.00104864 0 0.00104874 3.3 0.0010486599999999999 3.3 0.00104876 0 0.00104868 0 0.00104878 3.3 0.0010486999999999998 3.3 0.0010488 0 0.00104872 0 0.00104882 3.3 0.0010487399999999998 3.3 0.0010488399999999999 0 0.00104876 0 0.00104886 3.3 0.00104878 3.3 0.00104888 0 0.0010488 0 0.0010489 3.3 0.00104882 3.3 0.00104892 0 0.0010488399999999999 0 0.00104894 3.3 0.00104886 3.3 0.00104896 0 0.0010488799999999999 0 0.00104898 3.3 0.0010489 3.3 0.001049 0 0.0010489199999999998 0 0.00104902 3.3 0.00104894 3.3 0.00104904 0 0.0010489599999999998 0 0.0010490599999999999 3.3 0.00104898 3.3 0.00104908 0 0.001049 0 0.0010491 3.3 0.00104902 3.3 0.00104912 0 0.00104904 0 0.00104914 3.3 0.0010490599999999999 3.3 0.00104916 0 0.00104908 0 0.00104918 3.3 0.0010490999999999999 3.3 0.0010492 0 0.00104912 0 0.00104922 3.3 0.0010491399999999998 3.3 0.00104924 0 0.00104916 0 0.00104926 3.3 0.0010491799999999998 3.3 0.0010492799999999999 0 0.0010492 0 0.0010493 3.3 0.00104922 3.3 0.00104932 0 0.00104924 0 0.00104934 3.3 0.00104926 3.3 0.00104936 0 0.0010492799999999999 0 0.00104938 3.3 0.0010493 3.3 0.0010494 0 0.0010493199999999999 0 0.00104942 3.3 0.00104934 3.3 0.00104944 0 0.0010493599999999998 0 0.0010494599999999999 3.3 0.00104938 3.3 0.00104948 0 0.0010494 0 0.0010495 3.3 0.00104942 3.3 0.00104952 0 0.00104944 0 0.00104954 3.3 0.0010494599999999999 3.3 0.00104956 0 0.00104948 0 0.00104958 3.3 0.0010494999999999999 3.3 0.0010496 0 0.00104952 0 0.00104962 3.3 0.0010495399999999998 3.3 0.00104964 0 0.00104956 0 0.00104966 3.3 0.0010495799999999998 3.3 0.0010496799999999999 0 0.0010496 0 0.0010497 3.3 0.00104962 3.3 0.00104972 0 0.00104964 0 0.00104974 3.3 0.00104966 3.3 0.00104976 0 0.0010496799999999999 0 0.00104978 3.3 0.0010497 3.3 0.0010498 0 0.0010497199999999999 0 0.00104982 3.3 0.00104974 3.3 0.00104984 0 0.0010497599999999998 0 0.00104986 3.3 0.00104978 3.3 0.00104988 0 0.0010497999999999998 0 0.0010498999999999999 3.3 0.00104982 3.3 0.00104992 0 0.00104984 0 0.00104994 3.3 0.00104986 3.3 0.00104996 0 0.00104988 0 0.00104998 3.3 0.0010498999999999999 3.3 0.00105 0 0.00104992 0 0.00105002 3.3 0.0010499399999999999 3.3 0.00105004 0 0.00104996 0 0.00105006 3.3 0.0010499799999999998 3.3 0.00105008 0 0.00105 0 0.0010501 3.3 0.0010500199999999998 3.3 0.0010501199999999999 0 0.00105004 0 0.00105014 3.3 0.00105006 3.3 0.00105016 0 0.00105008 0 0.00105018 3.3 0.0010501 3.3 0.0010502 0 0.0010501199999999999 0 0.00105022 3.3 0.00105014 3.3 0.00105024 0 0.0010501599999999999 0 0.00105026 3.3 0.00105018 3.3 0.00105028 0 0.0010501999999999998 0 0.0010502999999999999 3.3 0.00105022 3.3 0.00105032 0 0.00105024 0 0.00105034 3.3 0.00105026 3.3 0.00105036 0 0.00105028 0 0.00105038 3.3 0.0010502999999999999 3.3 0.0010504 0 0.00105032 0 0.00105042 3.3 0.0010503399999999999 3.3 0.00105044 0 0.00105036 0 0.00105046 3.3 0.0010503799999999998 3.3 0.00105048 0 0.0010504 0 0.0010505 3.3 0.0010504199999999998 3.3 0.0010505199999999999 0 0.00105044 0 0.00105054 3.3 0.00105046 3.3 0.00105056 0 0.00105048 0 0.00105058 3.3 0.0010505 3.3 0.0010506 0 0.0010505199999999999 0 0.00105062 3.3 0.00105054 3.3 0.00105064 0 0.0010505599999999999 0 0.00105066 3.3 0.00105058 3.3 0.00105068 0 0.0010505999999999998 0 0.0010507 3.3 0.00105062 3.3 0.00105072 0 0.0010506399999999998 0 0.0010507399999999999 3.3 0.00105066 3.3 0.00105076 0 0.00105068 0 0.00105078 3.3 0.0010507 3.3 0.0010508 0 0.00105072 0 0.00105082 3.3 0.0010507399999999999 3.3 0.00105084 0 0.00105076 0 0.00105086 3.3 0.0010507799999999999 3.3 0.00105088 0 0.0010508 0 0.0010509 3.3 0.0010508199999999998 3.3 0.00105092 0 0.00105084 0 0.00105094 3.3 0.0010508599999999998 3.3 0.0010509599999999999 0 0.00105088 0 0.00105098 3.3 0.0010509 3.3 0.001051 0 0.00105092 0 0.00105102 3.3 0.00105094 3.3 0.00105104 0 0.0010509599999999999 0 0.00105106 3.3 0.00105098 3.3 0.00105108 0 0.0010509999999999999 0 0.0010511 3.3 0.00105102 3.3 0.00105112 0 0.0010510399999999998 0 0.0010511399999999999 3.3 0.00105106 3.3 0.00105116 0 0.00105108 0 0.00105118 3.3 0.0010511 3.3 0.0010512 0 0.00105112 0 0.00105122 3.3 0.0010511399999999999 3.3 0.00105124 0 0.00105116 0 0.00105126 3.3 0.0010511799999999999 3.3 0.00105128 0 0.0010512 0 0.0010513 3.3 0.0010512199999999998 3.3 0.00105132 0 0.00105124 0 0.00105134 3.3 0.0010512599999999998 3.3 0.0010513599999999999 0 0.00105128 0 0.00105138 3.3 0.0010513 3.3 0.0010514 0 0.00105132 0 0.00105142 3.3 0.00105134 3.3 0.00105144 0 0.0010513599999999999 0 0.00105146 3.3 0.00105138 3.3 0.00105148 0 0.0010513999999999999 0 0.0010515 3.3 0.00105142 3.3 0.00105152 0 0.0010514399999999998 0 0.00105154 3.3 0.00105146 3.3 0.00105156 0 0.0010514799999999998 0 0.0010515799999999999 3.3 0.0010515 3.3 0.0010516 0 0.00105152 0 0.00105162 3.3 0.00105154 3.3 0.00105164 0 0.00105156 0 0.00105166 3.3 0.0010515799999999999 3.3 0.00105168 0 0.0010516 0 0.0010517 3.3 0.0010516199999999999 3.3 0.00105172 0 0.00105164 0 0.00105174 3.3 0.0010516599999999998 3.3 0.0010517599999999999 0 0.00105168 0 0.00105178 3.3 0.0010516999999999998 3.3 0.0010517999999999999 0 0.00105172 0 0.00105182 3.3 0.00105174 3.3 0.00105184 0 0.0010517599999999999 0 0.00105186 3.3 0.00105178 3.3 0.00105188 0 0.0010517999999999999 0 0.0010519 3.3 0.00105182 3.3 0.00105192 0 0.0010518399999999998 0 0.00105194 3.3 0.00105186 3.3 0.00105196 0 0.0010518799999999998 0 0.0010519799999999999 3.3 0.0010519 3.3 0.001052 0 0.00105192 0 0.00105202 3.3 0.00105194 3.3 0.00105204 0 0.00105196 0 0.00105206 3.3 0.0010519799999999999 3.3 0.00105208 0 0.001052 0 0.0010521 3.3 0.0010520199999999999 3.3 0.00105212 0 0.00105204 0 0.00105214 3.3 0.0010520599999999998 3.3 0.00105216 0 0.00105208 0 0.00105218 3.3 0.0010520999999999998 3.3 0.0010521999999999999 0 0.00105212 0 0.00105222 3.3 0.00105214 3.3 0.00105224 0 0.00105216 0 0.00105226 3.3 0.00105218 3.3 0.00105228 0 0.0010521999999999999 0 0.0010523 3.3 0.00105222 3.3 0.00105232 0 0.0010522399999999999 0 0.00105234 3.3 0.00105226 3.3 0.00105236 0 0.0010522799999999998 0 0.00105238 3.3 0.0010523 3.3 0.0010524 0 0.0010523199999999998 0 0.0010524199999999999 3.3 0.00105234 3.3 0.00105244 0 0.00105236 0 0.00105246 3.3 0.00105238 3.3 0.00105248 0 0.0010524 0 0.0010525 3.3 0.0010524199999999999 3.3 0.00105252 0 0.00105244 0 0.00105254 3.3 0.0010524599999999999 3.3 0.00105256 0 0.00105248 0 0.00105258 3.3 0.0010524999999999998 3.3 0.0010525999999999999 0 0.00105252 0 0.00105262 3.3 0.00105254 3.3 0.00105264 0 0.00105256 0 0.00105266 3.3 0.00105258 3.3 0.00105268 0 0.0010525999999999999 0 0.0010527 3.3 0.00105262 3.3 0.00105272 0 0.0010526399999999999 0 0.00105274 3.3 0.00105266 3.3 0.00105276 0 0.0010526799999999998 0 0.00105278 3.3 0.0010527 3.3 0.0010528 0 0.0010527199999999998 0 0.0010528199999999999 3.3 0.00105274 3.3 0.00105284 0 0.00105276 0 0.00105286 3.3 0.00105278 3.3 0.00105288 0 0.0010528 0 0.0010529 3.3 0.0010528199999999999 3.3 0.00105292 0 0.00105284 0 0.00105294 3.3 0.0010528599999999999 3.3 0.00105296 0 0.00105288 0 0.00105298 3.3 0.0010528999999999998 3.3 0.001053 0 0.00105292 0 0.00105302 3.3 0.0010529399999999998 3.3 0.0010530399999999999 0 0.00105296 0 0.00105306 3.3 0.00105298 3.3 0.00105308 0 0.001053 0 0.0010531 3.3 0.00105302 3.3 0.00105312 0 0.0010530399999999999 0 0.00105314 3.3 0.00105306 3.3 0.00105316 0 0.0010530799999999999 0 0.00105318 3.3 0.0010531 3.3 0.0010532 0 0.0010531199999999998 0 0.00105322 3.3 0.00105314 3.3 0.00105324 0 0.0010531599999999998 0 0.0010532599999999999 3.3 0.00105318 3.3 0.00105328 0 0.0010532 0 0.0010533 3.3 0.00105322 3.3 0.00105332 0 0.00105324 0 0.00105334 3.3 0.0010532599999999999 3.3 0.00105336 0 0.00105328 0 0.00105338 3.3 0.0010532999999999999 3.3 0.0010534 0 0.00105332 0 0.00105342 3.3 0.0010533399999999998 3.3 0.0010534399999999999 0 0.00105336 0 0.00105346 3.3 0.00105338 3.3 0.00105348 0 0.0010534 0 0.0010535 3.3 0.00105342 3.3 0.00105352 0 0.0010534399999999999 0 0.00105354 3.3 0.00105346 3.3 0.00105356 0 0.0010534799999999999 0 0.00105358 3.3 0.0010535 3.3 0.0010536 0 0.0010535199999999998 0 0.00105362 3.3 0.00105354 3.3 0.00105364 0 0.0010535599999999998 0 0.0010536599999999999 3.3 0.00105358 3.3 0.00105368 0 0.0010536 0 0.0010537 3.3 0.00105362 3.3 0.00105372 0 0.00105364 0 0.00105374 3.3 0.0010536599999999999 3.3 0.00105376 0 0.00105368 0 0.00105378 3.3 0.0010536999999999999 3.3 0.0010538 0 0.00105372 0 0.00105382 3.3 0.0010537399999999998 3.3 0.00105384 0 0.00105376 0 0.00105386 3.3 0.0010537799999999998 3.3 0.0010538799999999999 0 0.0010538 0 0.0010539 3.3 0.00105382 3.3 0.00105392 0 0.00105384 0 0.00105394 3.3 0.00105386 3.3 0.00105396 0 0.0010538799999999999 0 0.00105398 3.3 0.0010539 3.3 0.001054 0 0.0010539199999999999 0 0.00105402 3.3 0.00105394 3.3 0.00105404 0 0.0010539599999999998 0 0.00105406 3.3 0.00105398 3.3 0.00105408 0 0.0010539999999999998 0 0.0010540999999999999 3.3 0.00105402 3.3 0.00105412 0 0.00105404 0 0.00105414 3.3 0.00105406 3.3 0.00105416 0 0.00105408 0 0.00105418 3.3 0.0010540999999999999 3.3 0.0010542 0 0.00105412 0 0.00105422 3.3 0.0010541399999999999 3.3 0.00105424 0 0.00105416 0 0.00105426 3.3 0.0010541799999999998 3.3 0.0010542799999999999 0 0.0010542 0 0.0010543 3.3 0.00105422 3.3 0.00105432 0 0.00105424 0 0.00105434 3.3 0.00105426 3.3 0.00105436 0 0.0010542799999999999 0 0.00105438 3.3 0.0010543 3.3 0.0010544 0 0.0010543199999999999 0 0.00105442 3.3 0.00105434 3.3 0.00105444 0 0.0010543599999999998 0 0.00105446 3.3 0.00105438 3.3 0.00105448 0 0.0010543999999999998 0 0.0010544999999999999 3.3 0.00105442 3.3 0.00105452 0 0.00105444 0 0.00105454 3.3 0.00105446 3.3 0.00105456 0 0.00105448 0 0.00105458 3.3 0.0010544999999999999 3.3 0.0010546 0 0.00105452 0 0.00105462 3.3 0.0010545399999999999 3.3 0.00105464 0 0.00105456 0 0.00105466 3.3 0.0010545799999999998 3.3 0.00105468 0 0.0010546 0 0.0010547 3.3 0.0010546199999999998 3.3 0.0010547199999999999 0 0.00105464 0 0.00105474 3.3 0.00105466 3.3 0.00105476 0 0.00105468 0 0.00105478 3.3 0.0010547 3.3 0.0010548 0 0.0010547199999999999 0 0.00105482 3.3 0.00105474 3.3 0.00105484 0 0.0010547599999999999 0 0.00105486 3.3 0.00105478 3.3 0.00105488 0 0.0010547999999999998 0 0.0010549 3.3 0.00105482 3.3 0.00105492 0 0.0010548399999999998 0 0.0010549399999999999 3.3 0.00105486 3.3 0.00105496 0 0.00105488 0 0.00105498 3.3 0.0010549 3.3 0.001055 0 0.00105492 0 0.00105502 3.3 0.0010549399999999999 3.3 0.00105504 0 0.00105496 0 0.00105506 3.3 0.0010549799999999999 3.3 0.00105508 0 0.001055 0 0.0010551 3.3 0.0010550199999999998 3.3 0.0010551199999999999 0 0.00105504 0 0.00105514 3.3 0.00105506 3.3 0.00105516 0 0.00105508 0 0.00105518 3.3 0.0010551 3.3 0.0010552 0 0.0010551199999999999 0 0.00105522 3.3 0.00105514 3.3 0.00105524 0 0.0010551599999999999 0 0.00105526 3.3 0.00105518 3.3 0.00105528 0 0.0010551999999999998 0 0.0010553 3.3 0.00105522 3.3 0.00105532 0 0.0010552399999999998 0 0.0010553399999999999 3.3 0.00105526 3.3 0.00105536 0 0.00105528 0 0.00105538 3.3 0.0010553 3.3 0.0010554 0 0.00105532 0 0.00105542 3.3 0.0010553399999999999 3.3 0.00105544 0 0.00105536 0 0.00105546 3.3 0.0010553799999999999 3.3 0.00105548 0 0.0010554 0 0.0010555 3.3 0.0010554199999999998 3.3 0.00105552 0 0.00105544 0 0.00105554 3.3 0.0010554599999999998 3.3 0.0010555599999999999 0 0.00105548 0 0.00105558 3.3 0.0010555 3.3 0.0010556 0 0.00105552 0 0.00105562 3.3 0.00105554 3.3 0.00105564 0 0.0010555599999999999 0 0.00105566 3.3 0.00105558 3.3 0.00105568 0 0.0010555999999999999 0 0.0010557 3.3 0.00105562 3.3 0.00105572 0 0.0010556399999999998 0 0.0010557399999999999 3.3 0.00105566 3.3 0.00105576 0 0.00105568 0 0.00105578 3.3 0.0010557 3.3 0.0010558 0 0.00105572 0 0.00105582 3.3 0.0010557399999999999 3.3 0.00105584 0 0.00105576 0 0.00105586 3.3 0.0010557799999999999 3.3 0.00105588 0 0.0010558 0 0.0010559 3.3 0.0010558199999999998 3.3 0.00105592 0 0.00105584 0 0.00105594 3.3 0.0010558599999999998 3.3 0.0010559599999999999 0 0.00105588 0 0.00105598 3.3 0.0010559 3.3 0.001056 0 0.00105592 0 0.00105602 3.3 0.00105594 3.3 0.00105604 0 0.0010559599999999999 0 0.00105606 3.3 0.00105598 3.3 0.00105608 0 0.0010559999999999999 0 0.0010561 3.3 0.00105602 3.3 0.00105612 0 0.0010560399999999998 0 0.00105614 3.3 0.00105606 3.3 0.00105616 0 0.0010560799999999998 0 0.0010561799999999999 3.3 0.0010561 3.3 0.0010562 0 0.00105612 0 0.00105622 3.3 0.00105614 3.3 0.00105624 0 0.00105616 0 0.00105626 3.3 0.0010561799999999999 3.3 0.00105628 0 0.0010562 0 0.0010563 3.3 0.0010562199999999999 3.3 0.00105632 0 0.00105624 0 0.00105634 3.3 0.0010562599999999998 3.3 0.00105636 0 0.00105628 0 0.00105638 3.3 0.0010562999999999998 3.3 0.0010563999999999999 0 0.00105632 0 0.00105642 3.3 0.00105634 3.3 0.00105644 0 0.00105636 0 0.00105646 3.3 0.00105638 3.3 0.00105648 0 0.0010563999999999999 0 0.0010565 3.3 0.00105642 3.3 0.00105652 0 0.0010564399999999999 0 0.00105654 3.3 0.00105646 3.3 0.00105656 0 0.0010564799999999998 0 0.0010565799999999999 3.3 0.0010565 3.3 0.0010566 0 0.00105652 0 0.00105662 3.3 0.00105654 3.3 0.00105664 0 0.00105656 0 0.00105666 3.3 0.0010565799999999999 3.3 0.00105668 0 0.0010566 0 0.0010567 3.3 0.0010566199999999999 3.3 0.00105672 0 0.00105664 0 0.00105674 3.3 0.0010566599999999998 3.3 0.00105676 0 0.00105668 0 0.00105678 3.3 0.0010566999999999998 3.3 0.0010567999999999999 0 0.00105672 0 0.00105682 3.3 0.00105674 3.3 0.00105684 0 0.00105676 0 0.00105686 3.3 0.00105678 3.3 0.00105688 0 0.0010567999999999999 0 0.0010569 3.3 0.00105682 3.3 0.00105692 0 0.0010568399999999999 0 0.00105694 3.3 0.00105686 3.3 0.00105696 0 0.0010568799999999998 0 0.00105698 3.3 0.0010569 3.3 0.001057 0 0.0010569199999999998 0 0.0010570199999999999 3.3 0.00105694 3.3 0.00105704 0 0.00105696 0 0.00105706 3.3 0.00105698 3.3 0.00105708 0 0.001057 0 0.0010571 3.3 0.0010570199999999999 3.3 0.00105712 0 0.00105704 0 0.00105714 3.3 0.0010570599999999999 3.3 0.00105716 0 0.00105708 0 0.00105718 3.3 0.0010570999999999998 3.3 0.0010572 0 0.00105712 0 0.00105722 3.3 0.0010571399999999998 3.3 0.0010572399999999999 0 0.00105716 0 0.00105726 3.3 0.00105718 3.3 0.00105728 0 0.0010572 0 0.0010573 3.3 0.00105722 3.3 0.00105732 0 0.0010572399999999999 0 0.00105734 3.3 0.00105726 3.3 0.00105736 0 0.0010572799999999999 0 0.00105738 3.3 0.0010573 3.3 0.0010574 0 0.0010573199999999998 0 0.0010574199999999999 3.3 0.00105734 3.3 0.00105744 0 0.00105736 0 0.00105746 3.3 0.00105738 3.3 0.00105748 0 0.0010574 0 0.0010575 3.3 0.0010574199999999999 3.3 0.00105752 0 0.00105744 0 0.00105754 3.3 0.0010574599999999999 3.3 0.00105756 0 0.00105748 0 0.00105758 3.3 0.0010574999999999998 3.3 0.0010576 0 0.00105752 0 0.00105762 3.3 0.0010575399999999998 3.3 0.0010576399999999999 0 0.00105756 0 0.00105766 3.3 0.00105758 3.3 0.00105768 0 0.0010576 0 0.0010577 3.3 0.00105762 3.3 0.00105772 0 0.0010576399999999999 0 0.00105774 3.3 0.00105766 3.3 0.00105776 0 0.0010576799999999999 0 0.00105778 3.3 0.0010577 3.3 0.0010578 0 0.0010577199999999998 0 0.00105782 3.3 0.00105774 3.3 0.00105784 0 0.0010577599999999998 0 0.0010578599999999999 3.3 0.00105778 3.3 0.00105788 0 0.0010578 0 0.0010579 3.3 0.00105782 3.3 0.00105792 0 0.00105784 0 0.00105794 3.3 0.0010578599999999999 3.3 0.00105796 0 0.00105788 0 0.00105798 3.3 0.0010578999999999999 3.3 0.001058 0 0.00105792 0 0.00105802 3.3 0.0010579399999999998 3.3 0.00105804 0 0.00105796 0 0.00105806 3.3 0.0010579799999999998 3.3 0.0010580799999999999 0 0.001058 0 0.0010581 3.3 0.00105802 3.3 0.00105812 0 0.00105804 0 0.00105814 3.3 0.00105806 3.3 0.00105816 0 0.0010580799999999999 0 0.00105818 3.3 0.0010581 3.3 0.0010582 0 0.0010581199999999999 0 0.00105822 3.3 0.00105814 3.3 0.00105824 0 0.0010581599999999998 0 0.0010582599999999999 3.3 0.00105818 3.3 0.00105828 0 0.0010582 0 0.0010583 3.3 0.00105822 3.3 0.00105832 0 0.00105824 0 0.00105834 3.3 0.0010582599999999999 3.3 0.00105836 0 0.00105828 0 0.00105838 3.3 0.0010582999999999999 3.3 0.0010584 0 0.00105832 0 0.00105842 3.3 0.0010583399999999998 3.3 0.00105844 0 0.00105836 0 0.00105846 3.3 0.0010583799999999998 3.3 0.0010584799999999999 0 0.0010584 0 0.0010585 3.3 0.00105842 3.3 0.00105852 0 0.00105844 0 0.00105854 3.3 0.00105846 3.3 0.00105856 0 0.0010584799999999999 0 0.00105858 3.3 0.0010585 3.3 0.0010586 0 0.0010585199999999999 0 0.00105862 3.3 0.00105854 3.3 0.00105864 0 0.0010585599999999998 0 0.00105866 3.3 0.00105858 3.3 0.00105868 0 0.0010585999999999998 0 0.0010586999999999999 3.3 0.00105862 3.3 0.00105872 0 0.00105864 0 0.00105874 3.3 0.00105866 3.3 0.00105876 0 0.00105868 0 0.00105878 3.3 0.0010586999999999999 3.3 0.0010588 0 0.00105872 0 0.00105882 3.3 0.0010587399999999999 3.3 0.00105884 0 0.00105876 0 0.00105886 3.3 0.0010587799999999998 3.3 0.0010588799999999999 0 0.0010588 0 0.0010589 3.3 0.00105882 3.3 0.00105892 0 0.00105884 0 0.00105894 3.3 0.00105886 3.3 0.00105896 0 0.0010588799999999999 0 0.00105898 3.3 0.0010589 3.3 0.001059 0 0.0010589199999999999 0 0.00105902 3.3 0.00105894 3.3 0.00105904 0 0.0010589599999999998 0 0.00105906 3.3 0.00105898 3.3 0.00105908 0 0.0010589999999999998 0 0.0010590999999999999 3.3 0.00105902 3.3 0.00105912 0 0.00105904 0 0.00105914 3.3 0.00105906 3.3 0.00105916 0 0.00105908 0 0.00105918 3.3 0.0010590999999999999 3.3 0.0010592 0 0.00105912 0 0.00105922 3.3 0.0010591399999999999 3.3 0.00105924 0 0.00105916 0 0.00105926 3.3 0.0010591799999999998 3.3 0.00105928 0 0.0010592 0 0.0010593 3.3 0.0010592199999999998 3.3 0.0010593199999999999 0 0.00105924 0 0.00105934 3.3 0.00105926 3.3 0.00105936 0 0.00105928 0 0.00105938 3.3 0.0010593 3.3 0.0010594 0 0.0010593199999999999 0 0.00105942 3.3 0.00105934 3.3 0.00105944 0 0.0010593599999999999 0 0.00105946 3.3 0.00105938 3.3 0.00105948 0 0.0010593999999999998 0 0.0010595 3.3 0.00105942 3.3 0.00105952 0 0.0010594399999999998 0 0.0010595399999999999 3.3 0.00105946 3.3 0.00105956 0 0.00105948 0 0.00105958 3.3 0.0010595 3.3 0.0010596 0 0.00105952 0 0.00105962 3.3 0.0010595399999999999 3.3 0.00105964 0 0.00105956 0 0.00105966 3.3 0.0010595799999999999 3.3 0.00105968 0 0.0010596 0 0.0010597 3.3 0.0010596199999999998 3.3 0.0010597199999999999 0 0.00105964 0 0.00105974 3.3 0.00105966 3.3 0.00105976 0 0.00105968 0 0.00105978 3.3 0.0010597 3.3 0.0010598 0 0.0010597199999999999 0 0.00105982 3.3 0.00105974 3.3 0.00105984 0 0.0010597599999999999 0 0.00105986 3.3 0.00105978 3.3 0.00105988 0 0.0010597999999999998 0 0.0010599 3.3 0.00105982 3.3 0.00105992 0 0.0010598399999999998 0 0.0010599399999999999 3.3 0.00105986 3.3 0.00105996 0 0.00105988 0 0.00105998 3.3 0.0010599 3.3 0.00106 0 0.00105992 0 0.00106002 3.3 0.0010599399999999999 3.3 0.00106004 0 0.00105996 0 0.00106006 3.3 0.0010599799999999999 3.3 0.00106008 0 0.00106 0 0.0010601 3.3 0.0010600199999999998 3.3 0.00106012 0 0.00106004 0 0.00106014 3.3 0.0010600599999999998 3.3 0.0010601599999999999 0 0.00106008 0 0.00106018 3.3 0.0010601 3.3 0.0010602 0 0.00106012 0 0.00106022 3.3 0.00106014 3.3 0.00106024 0 0.0010601599999999999 0 0.00106026 3.3 0.00106018 3.3 0.00106028 0 0.0010601999999999999 0 0.0010603 3.3 0.00106022 3.3 0.00106032 0 0.0010602399999999998 0 0.00106034 3.3 0.00106026 3.3 0.00106036 0 0.0010602799999999998 0 0.0010603799999999999 3.3 0.0010603 3.3 0.0010604 0 0.00106032 0 0.00106042 3.3 0.00106034 3.3 0.00106044 0 0.00106036 0 0.00106046 3.3 0.0010603799999999999 3.3 0.00106048 0 0.0010604 0 0.0010605 3.3 0.0010604199999999999 3.3 0.00106052 0 0.00106044 0 0.00106054 3.3 0.0010604599999999998 3.3 0.0010605599999999999 0 0.00106048 0 0.00106058 3.3 0.0010605 3.3 0.0010606 0 0.00106052 0 0.00106062 3.3 0.00106054 3.3 0.00106064 0 0.0010605599999999999 0 0.00106066 3.3 0.00106058 3.3 0.00106068 0 0.0010605999999999999 0 0.0010607 3.3 0.00106062 3.3 0.00106072 0 0.0010606399999999998 0 0.00106074 3.3 0.00106066 3.3 0.00106076 0 0.0010606799999999998 0 0.0010607799999999999 3.3 0.0010607 3.3 0.0010608 0 0.00106072 0 0.00106082 3.3 0.00106074 3.3 0.00106084 0 0.00106076 0 0.00106086 3.3 0.0010607799999999999 3.3 0.00106088 0 0.0010608 0 0.0010609 3.3 0.0010608199999999999 3.3 0.00106092 0 0.00106084 0 0.00106094 3.3 0.0010608599999999998 3.3 0.00106096 0 0.00106088 0 0.00106098 3.3 0.0010608999999999998 3.3 0.0010609999999999999 0 0.00106092 0 0.00106102 3.3 0.00106094 3.3 0.00106104 0 0.00106096 0 0.00106106 3.3 0.00106098 3.3 0.00106108 0 0.0010609999999999999 0 0.0010611 3.3 0.00106102 3.3 0.00106112 0 0.0010610399999999999 0 0.00106114 3.3 0.00106106 3.3 0.00106116 0 0.0010610799999999998 0 0.00106118 3.3 0.0010611 3.3 0.0010612 0 0.0010611199999999998 0 0.0010612199999999999 3.3 0.00106114 3.3 0.00106124 0 0.00106116 0 0.00106126 3.3 0.00106118 3.3 0.00106128 0 0.0010612 0 0.0010613 3.3 0.0010612199999999999 3.3 0.00106132 0 0.00106124 0 0.00106134 3.3 0.0010612599999999999 3.3 0.00106136 0 0.00106128 0 0.00106138 3.3 0.0010612999999999998 3.3 0.0010613999999999999 0 0.00106132 0 0.00106142 3.3 0.00106134 3.3 0.00106144 0 0.00106136 0 0.00106146 3.3 0.00106138 3.3 0.00106148 0 0.0010613999999999999 0 0.0010615 3.3 0.00106142 3.3 0.00106152 0 0.0010614399999999999 0 0.00106154 3.3 0.00106146 3.3 0.00106156 0 0.0010614799999999998 0 0.00106158 3.3 0.0010615 3.3 0.0010616 0 0.0010615199999999998 0 0.0010616199999999999 3.3 0.00106154 3.3 0.00106164 0 0.00106156 0 0.00106166 3.3 0.00106158 3.3 0.00106168 0 0.0010616 0 0.0010617 3.3 0.0010616199999999999 3.3 0.00106172 0 0.00106164 0 0.00106174 3.3 0.0010616599999999999 3.3 0.00106176 0 0.00106168 0 0.00106178 3.3 0.0010616999999999998 3.3 0.0010618 0 0.00106172 0 0.00106182 3.3 0.0010617399999999998 3.3 0.0010618399999999999 0 0.00106176 0 0.00106186 3.3 0.00106178 3.3 0.00106188 0 0.0010618 0 0.0010619 3.3 0.00106182 3.3 0.00106192 0 0.0010618399999999999 0 0.00106194 3.3 0.00106186 3.3 0.00106196 0 0.0010618799999999999 0 0.00106198 3.3 0.0010619 3.3 0.001062 0 0.0010619199999999998 0 0.0010620199999999999 3.3 0.00106194 3.3 0.00106204 0 0.0010619599999999998 0 0.0010620599999999999 3.3 0.00106198 3.3 0.00106208 0 0.001062 0 0.0010621 3.3 0.0010620199999999999 3.3 0.00106212 0 0.00106204 0 0.00106214 3.3 0.0010620599999999999 3.3 0.00106216 0 0.00106208 0 0.00106218 3.3 0.0010620999999999998 3.3 0.0010622 0 0.00106212 0 0.00106222 3.3 0.0010621399999999998 3.3 0.0010622399999999999 0 0.00106216 0 0.00106226 3.3 0.00106218 3.3 0.00106228 0 0.0010622 0 0.0010623 3.3 0.00106222 3.3 0.00106232 0 0.0010622399999999999 0 0.00106234 3.3 0.00106226 3.3 0.00106236 0 0.0010622799999999999 0 0.00106238 3.3 0.0010623 3.3 0.0010624 0 0.0010623199999999998 0 0.00106242 3.3 0.00106234 3.3 0.00106244 0 0.0010623599999999998 0 0.0010624599999999999 3.3 0.00106238 3.3 0.00106248 0 0.0010624 0 0.0010625 3.3 0.00106242 3.3 0.00106252 0 0.00106244 0 0.00106254 3.3 0.0010624599999999999 3.3 0.00106256 0 0.00106248 0 0.00106258 3.3 0.0010624999999999999 3.3 0.0010626 0 0.00106252 0 0.00106262 3.3 0.0010625399999999998 3.3 0.00106264 0 0.00106256 0 0.00106266 3.3 0.0010625799999999998 3.3 0.0010626799999999999 0 0.0010626 0 0.0010627 3.3 0.00106262 3.3 0.00106272 0 0.00106264 0 0.00106274 3.3 0.00106266 3.3 0.00106276 0 0.0010626799999999999 0 0.00106278 3.3 0.0010627 3.3 0.0010628 0 0.0010627199999999999 0 0.00106282 3.3 0.00106274 3.3 0.00106284 0 0.0010627599999999998 0 0.0010628599999999999 3.3 0.00106278 3.3 0.00106288 0 0.0010628 0 0.0010629 3.3 0.00106282 3.3 0.00106292 0 0.00106284 0 0.00106294 3.3 0.0010628599999999999 3.3 0.00106296 0 0.00106288 0 0.00106298 3.3 0.0010628999999999999 3.3 0.001063 0 0.00106292 0 0.00106302 3.3 0.0010629399999999998 3.3 0.00106304 0 0.00106296 0 0.00106306 3.3 0.0010629799999999998 3.3 0.0010630799999999999 0 0.001063 0 0.0010631 3.3 0.00106302 3.3 0.00106312 0 0.00106304 0 0.00106314 3.3 0.00106306 3.3 0.00106316 0 0.0010630799999999999 0 0.00106318 3.3 0.0010631 3.3 0.0010632 0 0.0010631199999999999 0 0.00106322 3.3 0.00106314 3.3 0.00106324 0 0.0010631599999999998 0 0.00106326 3.3 0.00106318 3.3 0.00106328 0 0.0010631999999999998 0 0.0010632999999999999 3.3 0.00106322 3.3 0.00106332 0 0.00106324 0 0.00106334 3.3 0.00106326 3.3 0.00106336 0 0.00106328 0 0.00106338 3.3 0.0010632999999999999 3.3 0.0010634 0 0.00106332 0 0.00106342 3.3 0.0010633399999999999 3.3 0.00106344 0 0.00106336 0 0.00106346 3.3 0.0010633799999999998 3.3 0.00106348 0 0.0010634 0 0.0010635 3.3 0.0010634199999999998 3.3 0.0010635199999999999 0 0.00106344 0 0.00106354 3.3 0.00106346 3.3 0.00106356 0 0.00106348 0 0.00106358 3.3 0.0010635 3.3 0.0010636 0 0.0010635199999999999 0 0.00106362 3.3 0.00106354 3.3 0.00106364 0 0.0010635599999999999 0 0.00106366 3.3 0.00106358 3.3 0.00106368 0 0.0010635999999999998 0 0.0010636999999999999 3.3 0.00106362 3.3 0.00106372 0 0.00106364 0 0.00106374 3.3 0.00106366 3.3 0.00106376 0 0.00106368 0 0.00106378 3.3 0.0010636999999999999 3.3 0.0010638 0 0.00106372 0 0.00106382 3.3 0.0010637399999999999 3.3 0.00106384 0 0.00106376 0 0.00106386 3.3 0.0010637799999999998 3.3 0.00106388 0 0.0010638 0 0.0010639 3.3 0.0010638199999999998 3.3 0.0010639199999999999 0 0.00106384 0 0.00106394 3.3 0.00106386 3.3 0.00106396 0 0.00106388 0 0.00106398 3.3 0.0010639 3.3 0.001064 0 0.0010639199999999999 0 0.00106402 3.3 0.00106394 3.3 0.00106404 0 0.0010639599999999999 0 0.00106406 3.3 0.00106398 3.3 0.00106408 0 0.0010639999999999998 0 0.0010641 3.3 0.00106402 3.3 0.00106412 0 0.0010640399999999998 0 0.0010641399999999999 3.3 0.00106406 3.3 0.00106416 0 0.00106408 0 0.00106418 3.3 0.0010641 3.3 0.0010642 0 0.00106412 0 0.00106422 3.3 0.0010641399999999999 3.3 0.00106424 0 0.00106416 0 0.00106426 3.3 0.0010641799999999999 3.3 0.00106428 0 0.0010642 0 0.0010643 3.3 0.0010642199999999998 3.3 0.00106432 0 0.00106424 0 0.00106434 3.3 0.0010642599999999998 3.3 0.0010643599999999999 0 0.00106428 0 0.00106438 3.3 0.0010643 3.3 0.0010644 0 0.00106432 0 0.00106442 3.3 0.00106434 3.3 0.00106444 0 0.0010643599999999999 0 0.00106446 3.3 0.00106438 3.3 0.00106448 0 0.0010643999999999999 0 0.0010645 3.3 0.00106442 3.3 0.00106452 0 0.0010644399999999998 0 0.0010645399999999999 3.3 0.00106446 3.3 0.00106456 0 0.00106448 0 0.00106458 3.3 0.0010645 3.3 0.0010646 0 0.00106452 0 0.00106462 3.3 0.0010645399999999999 3.3 0.00106464 0 0.00106456 0 0.00106466 3.3 0.0010645799999999999 3.3 0.00106468 0 0.0010646 0 0.0010647 3.3 0.0010646199999999998 3.3 0.00106472 0 0.00106464 0 0.00106474 3.3 0.0010646599999999998 3.3 0.0010647599999999999 0 0.00106468 0 0.00106478 3.3 0.0010647 3.3 0.0010648 0 0.00106472 0 0.00106482 3.3 0.00106474 3.3 0.00106484 0 0.0010647599999999999 0 0.00106486 3.3 0.00106478 3.3 0.00106488 0 0.0010647999999999999 0 0.0010649 3.3 0.00106482 3.3 0.00106492 0 0.0010648399999999998 0 0.00106494 3.3 0.00106486 3.3 0.00106496 0 0.0010648799999999998 0 0.0010649799999999999 3.3 0.0010649 3.3 0.001065 0 0.00106492 0 0.00106502 3.3 0.00106494 3.3 0.00106504 0 0.00106496 0 0.00106506 3.3 0.0010649799999999999 3.3 0.00106508 0 0.001065 0 0.0010651 3.3 0.0010650199999999999 3.3 0.00106512 0 0.00106504 0 0.00106514 3.3 0.0010650599999999998 3.3 0.00106516 0 0.00106508 0 0.00106518 3.3 0.0010650999999999998 3.3 0.0010651999999999999 0 0.00106512 0 0.00106522 3.3 0.00106514 3.3 0.00106524 0 0.00106516 0 0.00106526 3.3 0.00106518 3.3 0.00106528 0 0.0010651999999999999 0 0.0010653 3.3 0.00106522 3.3 0.00106532 0 0.0010652399999999999 0 0.00106534 3.3 0.00106526 3.3 0.00106536 0 0.0010652799999999998 0 0.0010653799999999999 3.3 0.0010653 3.3 0.0010654 0 0.00106532 0 0.00106542 3.3 0.00106534 3.3 0.00106544 0 0.00106536 0 0.00106546 3.3 0.0010653799999999999 3.3 0.00106548 0 0.0010654 0 0.0010655 3.3 0.0010654199999999999 3.3 0.00106552 0 0.00106544 0 0.00106554 3.3 0.0010654599999999998 3.3 0.00106556 0 0.00106548 0 0.00106558 3.3 0.0010654999999999998 3.3 0.0010655999999999999 0 0.00106552 0 0.00106562 3.3 0.00106554 3.3 0.00106564 0 0.00106556 0 0.00106566 3.3 0.00106558 3.3 0.00106568 0 0.0010655999999999999 0 0.0010657 3.3 0.00106562 3.3 0.00106572 0 0.0010656399999999999 0 0.00106574 3.3 0.00106566 3.3 0.00106576 0 0.0010656799999999998 0 0.00106578 3.3 0.0010657 3.3 0.0010658 0 0.0010657199999999998 0 0.0010658199999999999 3.3 0.00106574 3.3 0.00106584 0 0.00106576 0 0.00106586 3.3 0.00106578 3.3 0.00106588 0 0.0010658 0 0.0010659 3.3 0.0010658199999999999 3.3 0.00106592 0 0.00106584 0 0.00106594 3.3 0.0010658599999999999 3.3 0.00106596 0 0.00106588 0 0.00106598 3.3 0.0010658999999999998 3.3 0.0010659999999999999 0 0.00106592 0 0.00106602 3.3 0.00106594 3.3 0.00106604 0 0.00106596 0 0.00106606 3.3 0.00106598 3.3 0.00106608 0 0.0010659999999999999 0 0.0010661 3.3 0.00106602 3.3 0.00106612 0 0.0010660399999999999 0 0.00106614 3.3 0.00106606 3.3 0.00106616 0 0.0010660799999999998 0 0.00106618 3.3 0.0010661 3.3 0.0010662 0 0.0010661199999999998 0 0.0010662199999999999 3.3 0.00106614 3.3 0.00106624 0 0.00106616 0 0.00106626 3.3 0.00106618 3.3 0.00106628 0 0.0010662 0 0.0010663 3.3 0.0010662199999999999 3.3 0.00106632 0 0.00106624 0 0.00106634 3.3 0.0010662599999999999 3.3 0.00106636 0 0.00106628 0 0.00106638 3.3 0.0010662999999999998 3.3 0.0010664 0 0.00106632 0 0.00106642 3.3 0.0010663399999999998 3.3 0.0010664399999999999 0 0.00106636 0 0.00106646 3.3 0.00106638 3.3 0.00106648 0 0.0010664 0 0.0010665 3.3 0.00106642 3.3 0.00106652 0 0.0010664399999999999 0 0.00106654 3.3 0.00106646 3.3 0.00106656 0 0.0010664799999999999 0 0.00106658 3.3 0.0010665 3.3 0.0010666 0 0.0010665199999999998 0 0.00106662 3.3 0.00106654 3.3 0.00106664 0 0.0010665599999999998 0 0.0010666599999999999 3.3 0.00106658 3.3 0.00106668 0 0.0010666 0 0.0010667 3.3 0.00106662 3.3 0.00106672 0 0.00106664 0 0.00106674 3.3 0.0010666599999999999 3.3 0.00106676 0 0.00106668 0 0.00106678 3.3 0.0010666999999999999 3.3 0.0010668 0 0.00106672 0 0.00106682 3.3 0.0010667399999999998 3.3 0.0010668399999999999 0 0.00106676 0 0.00106686 3.3 0.00106678 3.3 0.00106688 0 0.0010668 0 0.0010669 3.3 0.00106682 3.3 0.00106692 0 0.0010668399999999999 0 0.00106694 3.3 0.00106686 3.3 0.00106696 0 0.0010668799999999999 0 0.00106698 3.3 0.0010669 3.3 0.001067 0 0.0010669199999999998 0 0.00106702 3.3 0.00106694 3.3 0.00106704 0 0.0010669599999999998 0 0.0010670599999999999 3.3 0.00106698 3.3 0.00106708 0 0.001067 0 0.0010671 3.3 0.00106702 3.3 0.00106712 0 0.00106704 0 0.00106714 3.3 0.0010670599999999999 3.3 0.00106716 0 0.00106708 0 0.00106718 3.3 0.0010670999999999999 3.3 0.0010672 0 0.00106712 0 0.00106722 3.3 0.0010671399999999998 3.3 0.00106724 0 0.00106716 0 0.00106726 3.3 0.0010671799999999998 3.3 0.0010672799999999999 0 0.0010672 0 0.0010673 3.3 0.00106722 3.3 0.00106732 0 0.00106724 0 0.00106734 3.3 0.00106726 3.3 0.00106736 0 0.0010672799999999999 0 0.00106738 3.3 0.0010673 3.3 0.0010674 0 0.0010673199999999999 0 0.00106742 3.3 0.00106734 3.3 0.00106744 0 0.0010673599999999998 0 0.00106746 3.3 0.00106738 3.3 0.00106748 0 0.0010673999999999998 0 0.0010674999999999999 3.3 0.00106742 3.3 0.00106752 0 0.00106744 0 0.00106754 3.3 0.00106746 3.3 0.00106756 0 0.00106748 0 0.00106758 3.3 0.0010674999999999999 3.3 0.0010676 0 0.00106752 0 0.00106762 3.3 0.0010675399999999999 3.3 0.00106764 0 0.00106756 0 0.00106766 3.3 0.0010675799999999998 3.3 0.0010676799999999999 0 0.0010676 0 0.0010677 3.3 0.00106762 3.3 0.00106772 0 0.00106764 0 0.00106774 3.3 0.00106766 3.3 0.00106776 0 0.0010676799999999999 0 0.00106778 3.3 0.0010677 3.3 0.0010678 0 0.0010677199999999999 0 0.00106782 3.3 0.00106774 3.3 0.00106784 0 0.0010677599999999998 0 0.00106786 3.3 0.00106778 3.3 0.00106788 0 0.0010677999999999998 0 0.0010678999999999999 3.3 0.00106782 3.3 0.00106792 0 0.00106784 0 0.00106794 3.3 0.00106786 3.3 0.00106796 0 0.00106788 0 0.00106798 3.3 0.0010678999999999999 3.3 0.001068 0 0.00106792 0 0.00106802 3.3 0.0010679399999999999 3.3 0.00106804 0 0.00106796 0 0.00106806 3.3 0.0010679799999999998 3.3 0.00106808 0 0.001068 0 0.0010681 3.3 0.0010680199999999998 3.3 0.0010681199999999999 0 0.00106804 0 0.00106814 3.3 0.00106806 3.3 0.00106816 0 0.00106808 0 0.00106818 3.3 0.0010681 3.3 0.0010682 0 0.0010681199999999999 0 0.00106822 3.3 0.00106814 3.3 0.00106824 0 0.0010681599999999999 0 0.00106826 3.3 0.00106818 3.3 0.00106828 0 0.0010681999999999998 0 0.0010683 3.3 0.00106822 3.3 0.00106832 0 0.0010682399999999998 0 0.0010683399999999999 3.3 0.00106826 3.3 0.00106836 0 0.00106828 0 0.00106838 3.3 0.0010683 3.3 0.0010684 0 0.00106832 0 0.00106842 3.3 0.0010683399999999999 3.3 0.00106844 0 0.00106836 0 0.00106846 3.3 0.0010683799999999999 3.3 0.00106848 0 0.0010684 0 0.0010685 3.3 0.0010684199999999998 3.3 0.0010685199999999999 0 0.00106844 0 0.00106854 3.3 0.00106846 3.3 0.00106856 0 0.00106848 0 0.00106858 3.3 0.0010685 3.3 0.0010686 0 0.0010685199999999999 0 0.00106862 3.3 0.00106854 3.3 0.00106864 0 0.0010685599999999999 0 0.00106866 3.3 0.00106858 3.3 0.00106868 0 0.0010685999999999998 0 0.0010687 3.3 0.00106862 3.3 0.00106872 0 0.0010686399999999998 0 0.0010687399999999999 3.3 0.00106866 3.3 0.00106876 0 0.00106868 0 0.00106878 3.3 0.0010687 3.3 0.0010688 0 0.00106872 0 0.00106882 3.3 0.0010687399999999999 3.3 0.00106884 0 0.00106876 0 0.00106886 3.3 0.0010687799999999999 3.3 0.00106888 0 0.0010688 0 0.0010689 3.3 0.0010688199999999998 3.3 0.00106892 0 0.00106884 0 0.00106894 3.3 0.0010688599999999998 3.3 0.0010689599999999999 0 0.00106888 0 0.00106898 3.3 0.0010689 3.3 0.001069 0 0.00106892 0 0.00106902 3.3 0.00106894 3.3 0.00106904 0 0.0010689599999999999 0 0.00106906 3.3 0.00106898 3.3 0.00106908 0 0.0010689999999999999 0 0.0010691 3.3 0.00106902 3.3 0.00106912 0 0.0010690399999999998 0 0.0010691399999999999 3.3 0.00106906 3.3 0.00106916 0 0.00106908 0 0.00106918 3.3 0.0010691 3.3 0.0010692 0 0.00106912 0 0.00106922 3.3 0.0010691399999999999 3.3 0.00106924 0 0.00106916 0 0.00106926 3.3 0.0010691799999999999 3.3 0.00106928 0 0.0010692 0 0.0010693 3.3 0.0010692199999999998 3.3 0.00106932 0 0.00106924 0 0.00106934 3.3 0.0010692599999999998 3.3 0.0010693599999999999 0 0.00106928 0 0.00106938 3.3 0.0010693 3.3 0.0010694 0 0.00106932 0 0.00106942 3.3 0.00106934 3.3 0.00106944 0 0.0010693599999999999 0 0.00106946 3.3 0.00106938 3.3 0.00106948 0 0.0010693999999999999 0 0.0010695 3.3 0.00106942 3.3 0.00106952 0 0.0010694399999999998 0 0.00106954 3.3 0.00106946 3.3 0.00106956 0 0.0010694799999999998 0 0.0010695799999999999 3.3 0.0010695 3.3 0.0010696 0 0.00106952 0 0.00106962 3.3 0.00106954 3.3 0.00106964 0 0.00106956 0 0.00106966 3.3 0.0010695799999999999 3.3 0.00106968 0 0.0010696 0 0.0010697 3.3 0.0010696199999999999 3.3 0.00106972 0 0.00106964 0 0.00106974 3.3 0.0010696599999999998 3.3 0.00106976 0 0.00106968 0 0.00106978 3.3 0.0010696999999999998 3.3 0.0010697999999999999 0 0.00106972 0 0.00106982 3.3 0.00106974 3.3 0.00106984 0 0.00106976 0 0.00106986 3.3 0.00106978 3.3 0.00106988 0 0.0010697999999999999 0 0.0010699 3.3 0.00106982 3.3 0.00106992 0 0.0010698399999999999 0 0.00106994 3.3 0.00106986 3.3 0.00106996 0 0.0010698799999999998 0 0.0010699799999999999 3.3 0.0010699 3.3 0.00107 0 0.00106992 0 0.00107002 3.3 0.00106994 3.3 0.00107004 0 0.00106996 0 0.00107006 3.3 0.0010699799999999999 3.3 0.00107008 0 0.00107 0 0.0010701 3.3 0.0010700199999999999 3.3 0.00107012 0 0.00107004 0 0.00107014 3.3 0.0010700599999999998 3.3 0.00107016 0 0.00107008 0 0.00107018 3.3 0.0010700999999999998 3.3 0.0010701999999999999 0 0.00107012 0 0.00107022 3.3 0.00107014 3.3 0.00107024 0 0.00107016 0 0.00107026 3.3 0.00107018 3.3 0.00107028 0 0.0010701999999999999 0 0.0010703 3.3 0.00107022 3.3 0.00107032 0 0.0010702399999999999 0 0.00107034 3.3 0.00107026 3.3 0.00107036 0 0.0010702799999999998 0 0.00107038 3.3 0.0010703 3.3 0.0010704 0 0.0010703199999999998 0 0.0010704199999999999 3.3 0.00107034 3.3 0.00107044 0 0.00107036 0 0.00107046 3.3 0.00107038 3.3 0.00107048 0 0.0010704 0 0.0010705 3.3 0.0010704199999999999 3.3 0.00107052 0 0.00107044 0 0.00107054 3.3 0.0010704599999999999 3.3 0.00107056 0 0.00107048 0 0.00107058 3.3 0.0010704999999999998 3.3 0.0010706 0 0.00107052 0 0.00107062 3.3 0.0010705399999999998 3.3 0.0010706399999999999 0 0.00107056 0 0.00107066 3.3 0.00107058 3.3 0.00107068 0 0.0010706 0 0.0010707 3.3 0.00107062 3.3 0.00107072 0 0.0010706399999999999 0 0.00107074 3.3 0.00107066 3.3 0.00107076 0 0.0010706799999999999 0 0.00107078 3.3 0.0010707 3.3 0.0010708 0 0.0010707199999999998 0 0.0010708199999999999 3.3 0.00107074 3.3 0.00107084 0 0.00107076 0 0.00107086 3.3 0.00107078 3.3 0.00107088 0 0.0010708 0 0.0010709 3.3 0.0010708199999999999 3.3 0.00107092 0 0.00107084 0 0.00107094 3.3 0.0010708599999999999 3.3 0.00107096 0 0.00107088 0 0.00107098 3.3 0.0010708999999999998 3.3 0.001071 0 0.00107092 0 0.00107102 3.3 0.0010709399999999998 3.3 0.0010710399999999999 0 0.00107096 0 0.00107106 3.3 0.00107098 3.3 0.00107108 0 0.001071 0 0.0010711 3.3 0.00107102 3.3 0.00107112 0 0.0010710399999999999 0 0.00107114 3.3 0.00107106 3.3 0.00107116 0 0.0010710799999999999 0 0.00107118 3.3 0.0010711 3.3 0.0010712 0 0.0010711199999999998 0 0.00107122 3.3 0.00107114 3.3 0.00107124 0 0.0010711599999999998 0 0.0010712599999999999 3.3 0.00107118 3.3 0.00107128 0 0.0010712 0 0.0010713 3.3 0.00107122 3.3 0.00107132 0 0.00107124 0 0.00107134 3.3 0.0010712599999999999 3.3 0.00107136 0 0.00107128 0 0.00107138 3.3 0.0010712999999999999 3.3 0.0010714 0 0.00107132 0 0.00107142 3.3 0.0010713399999999998 3.3 0.00107144 0 0.00107136 0 0.00107146 3.3 0.0010713799999999998 3.3 0.0010714799999999999 0 0.0010714 0 0.0010715 3.3 0.00107142 3.3 0.00107152 0 0.00107144 0 0.00107154 3.3 0.00107146 3.3 0.00107156 0 0.0010714799999999999 0 0.00107158 3.3 0.0010715 3.3 0.0010716 0 0.0010715199999999999 0 0.00107162 3.3 0.00107154 3.3 0.00107164 0 0.0010715599999999998 0 0.0010716599999999999 3.3 0.00107158 3.3 0.00107168 0 0.0010716 0 0.0010717 3.3 0.00107162 3.3 0.00107172 0 0.00107164 0 0.00107174 3.3 0.0010716599999999999 3.3 0.00107176 0 0.00107168 0 0.00107178 3.3 0.0010716999999999999 3.3 0.0010718 0 0.00107172 0 0.00107182 3.3 0.0010717399999999998 3.3 0.00107184 0 0.00107176 0 0.00107186 3.3 0.0010717799999999998 3.3 0.0010718799999999999 0 0.0010718 0 0.0010719 3.3 0.00107182 3.3 0.00107192 0 0.00107184 0 0.00107194 3.3 0.00107186 3.3 0.00107196 0 0.0010718799999999999 0 0.00107198 3.3 0.0010719 3.3 0.001072 0 0.0010719199999999999 0 0.00107202 3.3 0.00107194 3.3 0.00107204 0 0.0010719599999999998 0 0.00107206 3.3 0.00107198 3.3 0.00107208 0 0.0010719999999999998 0 0.0010720999999999999 3.3 0.00107202 3.3 0.00107212 0 0.00107204 0 0.00107214 3.3 0.00107206 3.3 0.00107216 0 0.00107208 0 0.00107218 3.3 0.0010720999999999999 3.3 0.0010722 0 0.00107212 0 0.00107222 3.3 0.0010721399999999999 3.3 0.00107224 0 0.00107216 0 0.00107226 3.3 0.0010721799999999998 3.3 0.0010722799999999999 0 0.0010722 0 0.0010723 3.3 0.0010722199999999998 3.3 0.0010723199999999999 0 0.00107224 0 0.00107234 3.3 0.00107226 3.3 0.00107236 0 0.0010722799999999999 0 0.00107238 3.3 0.0010723 3.3 0.0010724 0 0.0010723199999999999 0 0.00107242 3.3 0.00107234 3.3 0.00107244 0 0.0010723599999999998 0 0.00107246 3.3 0.00107238 3.3 0.00107248 0 0.0010723999999999998 0 0.0010724999999999999 3.3 0.00107242 3.3 0.00107252 0 0.00107244 0 0.00107254 3.3 0.00107246 3.3 0.00107256 0 0.00107248 0 0.00107258 3.3 0.0010724999999999999 3.3 0.0010726 0 0.00107252 0 0.00107262 3.3 0.0010725399999999999 3.3 0.00107264 0 0.00107256 0 0.00107266 3.3 0.0010725799999999998 3.3 0.00107268 0 0.0010726 0 0.0010727 3.3 0.0010726199999999998 3.3 0.0010727199999999999 0 0.00107264 0 0.00107274 3.3 0.00107266 3.3 0.00107276 0 0.00107268 0 0.00107278 3.3 0.0010727 3.3 0.0010728 0 0.0010727199999999999 0 0.00107282 3.3 0.00107274 3.3 0.00107284 0 0.0010727599999999999 0 0.00107286 3.3 0.00107278 3.3 0.00107288 0 0.0010727999999999998 0 0.0010729 3.3 0.00107282 3.3 0.00107292 0 0.0010728399999999998 0 0.0010729399999999999 3.3 0.00107286 3.3 0.00107296 0 0.00107288 0 0.00107298 3.3 0.0010729 3.3 0.001073 0 0.00107292 0 0.00107302 3.3 0.0010729399999999999 3.3 0.00107304 0 0.00107296 0 0.00107306 3.3 0.0010729799999999999 3.3 0.00107308 0 0.001073 0 0.0010731 3.3 0.0010730199999999998 3.3 0.0010731199999999999 0 0.00107304 0 0.00107314 3.3 0.00107306 3.3 0.00107316 0 0.00107308 0 0.00107318 3.3 0.0010731 3.3 0.0010732 0 0.0010731199999999999 0 0.00107322 3.3 0.00107314 3.3 0.00107324 0 0.0010731599999999999 0 0.00107326 3.3 0.00107318 3.3 0.00107328 0 0.0010731999999999998 0 0.0010733 3.3 0.00107322 3.3 0.00107332 0 0.0010732399999999998 0 0.0010733399999999999 3.3 0.00107326 3.3 0.00107336 0 0.00107328 0 0.00107338 3.3 0.0010733 3.3 0.0010734 0 0.00107332 0 0.00107342 3.3 0.0010733399999999999 3.3 0.00107344 0 0.00107336 0 0.00107346 3.3 0.0010733799999999999 3.3 0.00107348 0 0.0010734 0 0.0010735 3.3 0.0010734199999999998 3.3 0.00107352 0 0.00107344 0 0.00107354 3.3 0.0010734599999999998 3.3 0.0010735599999999999 0 0.00107348 0 0.00107358 3.3 0.0010735 3.3 0.0010736 0 0.00107352 0 0.00107362 3.3 0.00107354 3.3 0.00107364 0 0.0010735599999999999 0 0.00107366 3.3 0.00107358 3.3 0.00107368 0 0.0010735999999999999 0 0.0010737 3.3 0.00107362 3.3 0.00107372 0 0.0010736399999999998 0 0.00107374 3.3 0.00107366 3.3 0.00107376 0 0.0010736799999999998 0 0.0010737799999999999 3.3 0.0010737 3.3 0.0010738 0 0.00107372 0 0.00107382 3.3 0.00107374 3.3 0.00107384 0 0.00107376 0 0.00107386 3.3 0.0010737799999999999 3.3 0.00107388 0 0.0010738 0 0.0010739 3.3 0.0010738199999999999 3.3 0.00107392 0 0.00107384 0 0.00107394 3.3 0.0010738599999999998 3.3 0.0010739599999999999 0 0.00107388 0 0.00107398 3.3 0.0010739 3.3 0.001074 0 0.00107392 0 0.00107402 3.3 0.00107394 3.3 0.00107404 0 0.0010739599999999999 0 0.00107406 3.3 0.00107398 3.3 0.00107408 0 0.0010739999999999999 0 0.0010741 3.3 0.00107402 3.3 0.00107412 0 0.0010740399999999998 0 0.00107414 3.3 0.00107406 3.3 0.00107416 0 0.0010740799999999998 0 0.0010741799999999999 3.3 0.0010741 3.3 0.0010742 0 0.00107412 0 0.00107422 3.3 0.00107414 3.3 0.00107424 0 0.00107416 0 0.00107426 3.3 0.0010741799999999999 3.3 0.00107428 0 0.0010742 0 0.0010743 3.3 0.0010742199999999999 3.3 0.00107432 0 0.00107424 0 0.00107434 3.3 0.0010742599999999998 3.3 0.00107436 0 0.00107428 0 0.00107438 3.3 0.0010742999999999998 3.3 0.0010743999999999999 0 0.00107432 0 0.00107442 3.3 0.00107434 3.3 0.00107444 0 0.00107436 0 0.00107446 3.3 0.00107438 3.3 0.00107448 0 0.0010743999999999999 0 0.0010745 3.3 0.00107442 3.3 0.00107452 0 0.0010744399999999999 0 0.00107454 3.3 0.00107446 3.3 0.00107456 0 0.0010744799999999998 0 0.00107458 3.3 0.0010745 3.3 0.0010746 0 0.0010745199999999998 0 0.0010746199999999999 3.3 0.00107454 3.3 0.00107464 0 0.00107456 0 0.00107466 3.3 0.00107458 3.3 0.00107468 0 0.0010746 0 0.0010747 3.3 0.0010746199999999999 3.3 0.00107472 0 0.00107464 0 0.00107474 3.3 0.0010746599999999999 3.3 0.00107476 0 0.00107468 0 0.00107478 3.3 0.0010746999999999998 3.3 0.0010747999999999999 0 0.00107472 0 0.00107482 3.3 0.00107474 3.3 0.00107484 0 0.00107476 0 0.00107486 3.3 0.00107478 3.3 0.00107488 0 0.0010747999999999999 0 0.0010749 3.3 0.00107482 3.3 0.00107492 0 0.0010748399999999999 0 0.00107494 3.3 0.00107486 3.3 0.00107496 0 0.0010748799999999998 0 0.00107498 3.3 0.0010749 3.3 0.001075 0 0.0010749199999999998 0 0.0010750199999999999 3.3 0.00107494 3.3 0.00107504 0 0.00107496 0 0.00107506 3.3 0.00107498 3.3 0.00107508 0 0.001075 0 0.0010751 3.3 0.0010750199999999999 3.3 0.00107512 0 0.00107504 0 0.00107514 3.3 0.0010750599999999999 3.3 0.00107516 0 0.00107508 0 0.00107518 3.3 0.0010750999999999998 3.3 0.0010752 0 0.00107512 0 0.00107522 3.3 0.0010751399999999998 3.3 0.0010752399999999999 0 0.00107516 0 0.00107526 3.3 0.00107518 3.3 0.00107528 0 0.0010752 0 0.0010753 3.3 0.00107522 3.3 0.00107532 0 0.0010752399999999999 0 0.00107534 3.3 0.00107526 3.3 0.00107536 0 0.0010752799999999999 0 0.00107538 3.3 0.0010753 3.3 0.0010754 0 0.0010753199999999998 0 0.00107542 3.3 0.00107534 3.3 0.00107544 0 0.0010753599999999998 0 0.0010754599999999999 3.3 0.00107538 3.3 0.00107548 0 0.0010754 0 0.0010755 3.3 0.00107542 3.3 0.00107552 0 0.00107544 0 0.00107554 3.3 0.0010754599999999999 3.3 0.00107556 0 0.00107548 0 0.00107558 3.3 0.0010754999999999999 3.3 0.0010756 0 0.00107552 0 0.00107562 3.3 0.0010755399999999998 3.3 0.0010756399999999999 0 0.00107556 0 0.00107566 3.3 0.00107558 3.3 0.00107568 0 0.0010756 0 0.0010757 3.3 0.00107562 3.3 0.00107572 0 0.0010756399999999999 0 0.00107574 3.3 0.00107566 3.3 0.00107576 0 0.0010756799999999999 0 0.00107578 3.3 0.0010757 3.3 0.0010758 0 0.0010757199999999998 0 0.00107582 3.3 0.00107574 3.3 0.00107584 0 0.0010757599999999998 0 0.0010758599999999999 3.3 0.00107578 3.3 0.00107588 0 0.0010758 0 0.0010759 3.3 0.00107582 3.3 0.00107592 0 0.00107584 0 0.00107594 3.3 0.0010758599999999999 3.3 0.00107596 0 0.00107588 0 0.00107598 3.3 0.0010758999999999999 3.3 0.001076 0 0.00107592 0 0.00107602 3.3 0.0010759399999999998 3.3 0.00107604 0 0.00107596 0 0.00107606 3.3 0.0010759799999999998 3.3 0.0010760799999999999 0 0.001076 0 0.0010761 3.3 0.00107602 3.3 0.00107612 0 0.00107604 0 0.00107614 3.3 0.00107606 3.3 0.00107616 0 0.0010760799999999999 0 0.00107618 3.3 0.0010761 3.3 0.0010762 0 0.0010761199999999999 0 0.00107622 3.3 0.00107614 3.3 0.00107624 0 0.0010761599999999998 0 0.0010762599999999999 3.3 0.00107618 3.3 0.00107628 0 0.0010762 0 0.0010763 3.3 0.00107622 3.3 0.00107632 0 0.00107624 0 0.00107634 3.3 0.0010762599999999999 3.3 0.00107636 0 0.00107628 0 0.00107638 3.3 0.0010762999999999999 3.3 0.0010764 0 0.00107632 0 0.00107642 3.3 0.0010763399999999998 3.3 0.00107644 0 0.00107636 0 0.00107646 3.3 0.0010763799999999998 3.3 0.0010764799999999999 0 0.0010764 0 0.0010765 3.3 0.00107642 3.3 0.00107652 0 0.00107644 0 0.00107654 3.3 0.00107646 3.3 0.00107656 0 0.0010764799999999999 0 0.00107658 3.3 0.0010765 3.3 0.0010766 0 0.0010765199999999999 0 0.00107662 3.3 0.00107654 3.3 0.00107664 0 0.0010765599999999998 0 0.00107666 3.3 0.00107658 3.3 0.00107668 0 0.0010765999999999998 0 0.0010766999999999999 3.3 0.00107662 3.3 0.00107672 0 0.00107664 0 0.00107674 3.3 0.00107666 3.3 0.00107676 0 0.00107668 0 0.00107678 3.3 0.0010766999999999999 3.3 0.0010768 0 0.00107672 0 0.00107682 3.3 0.0010767399999999999 3.3 0.00107684 0 0.00107676 0 0.00107686 3.3 0.0010767799999999998 3.3 0.00107688 0 0.0010768 0 0.0010769 3.3 0.0010768199999999998 3.3 0.0010769199999999999 0 0.00107684 0 0.00107694 3.3 0.00107686 3.3 0.00107696 0 0.00107688 0 0.00107698 3.3 0.0010769 3.3 0.001077 0 0.0010769199999999999 0 0.00107702 3.3 0.00107694 3.3 0.00107704 0 0.0010769599999999999 0 0.00107706 3.3 0.00107698 3.3 0.00107708 0 0.0010769999999999998 0 0.0010770999999999999 3.3 0.00107702 3.3 0.00107712 0 0.00107704 0 0.00107714 3.3 0.00107706 3.3 0.00107716 0 0.00107708 0 0.00107718 3.3 0.0010770999999999999 3.3 0.0010772 0 0.00107712 0 0.00107722 3.3 0.0010771399999999999 3.3 0.00107724 0 0.00107716 0 0.00107726 3.3 0.0010771799999999998 3.3 0.00107728 0 0.0010772 0 0.0010773 3.3 0.0010772199999999998 3.3 0.0010773199999999999 0 0.00107724 0 0.00107734 3.3 0.00107726 3.3 0.00107736 0 0.00107728 0 0.00107738 3.3 0.0010773 3.3 0.0010774 0 0.0010773199999999999 0 0.00107742 3.3 0.00107734 3.3 0.00107744 0 0.0010773599999999999 0 0.00107746 3.3 0.00107738 3.3 0.00107748 0 0.0010773999999999998 0 0.0010775 3.3 0.00107742 3.3 0.00107752 0 0.0010774399999999998 0 0.0010775399999999999 3.3 0.00107746 3.3 0.00107756 0 0.00107748 0 0.00107758 3.3 0.0010775 3.3 0.0010776 0 0.00107752 0 0.00107762 3.3 0.0010775399999999999 3.3 0.00107764 0 0.00107756 0 0.00107766 3.3 0.0010775799999999999 3.3 0.00107768 0 0.0010776 0 0.0010777 3.3 0.0010776199999999998 3.3 0.00107772 0 0.00107764 0 0.00107774 3.3 0.0010776599999999998 3.3 0.0010777599999999999 0 0.00107768 0 0.00107778 3.3 0.0010777 3.3 0.0010778 0 0.00107772 0 0.00107782 3.3 0.00107774 3.3 0.00107784 0 0.0010777599999999999 0 0.00107786 3.3 0.00107778 3.3 0.00107788 0 0.0010777999999999999 0 0.0010779 3.3 0.00107782 3.3 0.00107792 0 0.0010778399999999998 0 0.0010779399999999999 3.3 0.00107786 3.3 0.00107796 0 0.00107788 0 0.00107798 3.3 0.0010779 3.3 0.001078 0 0.00107792 0 0.00107802 3.3 0.0010779399999999999 3.3 0.00107804 0 0.00107796 0 0.00107806 3.3 0.0010779799999999999 3.3 0.00107808 0 0.001078 0 0.0010781 3.3 0.0010780199999999998 3.3 0.00107812 0 0.00107804 0 0.00107814 3.3 0.0010780599999999998 3.3 0.0010781599999999999 0 0.00107808 0 0.00107818 3.3 0.0010781 3.3 0.0010782 0 0.00107812 0 0.00107822 3.3 0.00107814 3.3 0.00107824 0 0.0010781599999999999 0 0.00107826 3.3 0.00107818 3.3 0.00107828 0 0.0010781999999999999 0 0.0010783 3.3 0.00107822 3.3 0.00107832 0 0.0010782399999999998 0 0.00107834 3.3 0.00107826 3.3 0.00107836 0 0.0010782799999999998 0 0.0010783799999999999 3.3 0.0010783 3.3 0.0010784 0 0.00107832 0 0.00107842 3.3 0.00107834 3.3 0.00107844 0 0.00107836 0 0.00107846 3.3 0.0010783799999999999 3.3 0.00107848 0 0.0010784 0 0.0010785 3.3 0.0010784199999999999 3.3 0.00107852 0 0.00107844 0 0.00107854 3.3 0.0010784599999999998 3.3 0.00107856 0 0.00107848 0 0.00107858 3.3 0.0010784999999999998 3.3 0.0010785999999999999 0 0.00107852 0 0.00107862 3.3 0.00107854 3.3 0.00107864 0 0.00107856 0 0.00107866 3.3 0.00107858 3.3 0.00107868 0 0.0010785999999999999 0 0.0010787 3.3 0.00107862 3.3 0.00107872 0 0.0010786399999999999 0 0.00107874 3.3 0.00107866 3.3 0.00107876 0 0.0010786799999999998 0 0.0010787799999999999 3.3 0.0010787 3.3 0.0010788 0 0.00107872 0 0.00107882 3.3 0.00107874 3.3 0.00107884 0 0.00107876 0 0.00107886 3.3 0.0010787799999999999 3.3 0.00107888 0 0.0010788 0 0.0010789 3.3 0.0010788199999999999 3.3 0.00107892 0 0.00107884 0 0.00107894 3.3 0.0010788599999999998 3.3 0.00107896 0 0.00107888 0 0.00107898 3.3 0.0010788999999999998 3.3 0.0010789999999999999 0 0.00107892 0 0.00107902 3.3 0.00107894 3.3 0.00107904 0 0.00107896 0 0.00107906 3.3 0.00107898 3.3 0.00107908 0 0.0010789999999999999 0 0.0010791 3.3 0.00107902 3.3 0.00107912 0 0.0010790399999999999 0 0.00107914 3.3 0.00107906 3.3 0.00107916 0 0.0010790799999999998 0 0.00107918 3.3 0.0010791 3.3 0.0010792 0 0.0010791199999999998 0 0.0010792199999999999 3.3 0.00107914 3.3 0.00107924 0 0.00107916 0 0.00107926 3.3 0.00107918 3.3 0.00107928 0 0.0010792 0 0.0010793 3.3 0.0010792199999999999 3.3 0.00107932 0 0.00107924 0 0.00107934 3.3 0.0010792599999999999 3.3 0.00107936 0 0.00107928 0 0.00107938 3.3 0.0010792999999999998 3.3 0.0010793999999999999 0 0.00107932 0 0.00107942 3.3 0.0010793399999999998 3.3 0.0010794399999999999 0 0.00107936 0 0.00107946 3.3 0.00107938 3.3 0.00107948 0 0.0010793999999999999 0 0.0010795 3.3 0.00107942 3.3 0.00107952 0 0.0010794399999999999 0 0.00107954 3.3 0.00107946 3.3 0.00107956 0 0.0010794799999999998 0 0.00107958 3.3 0.0010795 3.3 0.0010796 0 0.0010795199999999998 0 0.0010796199999999999 3.3 0.00107954 3.3 0.00107964 0 0.00107956 0 0.00107966 3.3 0.00107958 3.3 0.00107968 0 0.0010796 0 0.0010797 3.3 0.0010796199999999999 3.3 0.00107972 0 0.00107964 0 0.00107974 3.3 0.0010796599999999999 3.3 0.00107976 0 0.00107968 0 0.00107978 3.3 0.0010796999999999998 3.3 0.0010798 0 0.00107972 0 0.00107982 3.3 0.0010797399999999998 3.3 0.0010798399999999999 0 0.00107976 0 0.00107986 3.3 0.00107978 3.3 0.00107988 0 0.0010798 0 0.0010799 3.3 0.00107982 3.3 0.00107992 0 0.0010798399999999999 0 0.00107994 3.3 0.00107986 3.3 0.00107996 0 0.0010798799999999999 0 0.00107998 3.3 0.0010799 3.3 0.00108 0 0.0010799199999999998 0 0.00108002 3.3 0.00107994 3.3 0.00108004 0 0.0010799599999999998 0 0.0010800599999999999 3.3 0.00107998 3.3 0.00108008 0 0.00108 0 0.0010801 3.3 0.00108002 3.3 0.00108012 0 0.00108004 0 0.00108014 3.3 0.0010800599999999999 3.3 0.00108016 0 0.00108008 0 0.00108018 3.3 0.0010800999999999999 3.3 0.0010802 0 0.00108012 0 0.00108022 3.3 0.0010801399999999998 3.3 0.0010802399999999999 0 0.00108016 0 0.00108026 3.3 0.00108018 3.3 0.00108028 0 0.0010802 0 0.0010803 3.3 0.00108022 3.3 0.00108032 0 0.0010802399999999999 0 0.00108034 3.3 0.00108026 3.3 0.00108036 0 0.0010802799999999999 0 0.00108038 3.3 0.0010803 3.3 0.0010804 0 0.0010803199999999998 0 0.00108042 3.3 0.00108034 3.3 0.00108044 0 0.0010803599999999998 0 0.0010804599999999999 3.3 0.00108038 3.3 0.00108048 0 0.0010804 0 0.0010805 3.3 0.00108042 3.3 0.00108052 0 0.00108044 0 0.00108054 3.3 0.0010804599999999999 3.3 0.00108056 0 0.00108048 0 0.00108058 3.3 0.0010804999999999999 3.3 0.0010806 0 0.00108052 0 0.00108062 3.3 0.0010805399999999998 3.3 0.00108064 0 0.00108056 0 0.00108066 3.3 0.0010805799999999998 3.3 0.0010806799999999999 0 0.0010806 0 0.0010807 3.3 0.00108062 3.3 0.00108072 0 0.00108064 0 0.00108074 3.3 0.00108066 3.3 0.00108076 0 0.0010806799999999999 0 0.00108078 3.3 0.0010807 3.3 0.0010808 0 0.0010807199999999999 0 0.00108082 3.3 0.00108074 3.3 0.00108084 0 0.0010807599999999998 0 0.00108086 3.3 0.00108078 3.3 0.00108088 0 0.0010807999999999998 0 0.0010808999999999999 3.3 0.00108082 3.3 0.00108092 0 0.00108084 0 0.00108094 3.3 0.00108086 3.3 0.00108096 0 0.00108088 0 0.00108098 3.3 0.0010808999999999999 3.3 0.001081 0 0.00108092 0 0.00108102 3.3 0.0010809399999999999 3.3 0.00108104 0 0.00108096 0 0.00108106 3.3 0.0010809799999999998 3.3 0.0010810799999999999 0 0.001081 0 0.0010811 3.3 0.00108102 3.3 0.00108112 0 0.00108104 0 0.00108114 3.3 0.00108106 3.3 0.00108116 0 0.0010810799999999999 0 0.00108118 3.3 0.0010811 3.3 0.0010812 0 0.0010811199999999999 0 0.00108122 3.3 0.00108114 3.3 0.00108124 0 0.0010811599999999998 0 0.00108126 3.3 0.00108118 3.3 0.00108128 0 0.0010811999999999998 0 0.0010812999999999999 3.3 0.00108122 3.3 0.00108132 0 0.00108124 0 0.00108134 3.3 0.00108126 3.3 0.00108136 0 0.00108128 0 0.00108138 3.3 0.0010812999999999999 3.3 0.0010814 0 0.00108132 0 0.00108142 3.3 0.0010813399999999999 3.3 0.00108144 0 0.00108136 0 0.00108146 3.3 0.0010813799999999998 3.3 0.00108148 0 0.0010814 0 0.0010815 3.3 0.0010814199999999998 3.3 0.0010815199999999999 0 0.00108144 0 0.00108154 3.3 0.00108146 3.3 0.00108156 0 0.00108148 0 0.00108158 3.3 0.0010815 3.3 0.0010816 0 0.0010815199999999999 0 0.00108162 3.3 0.00108154 3.3 0.00108164 0 0.0010815599999999999 0 0.00108166 3.3 0.00108158 3.3 0.00108168 0 0.0010815999999999998 0 0.0010817 3.3 0.00108162 3.3 0.00108172 0 0.0010816399999999998 0 0.0010817399999999999 3.3 0.00108166 3.3 0.00108176 0 0.00108168 0 0.00108178 3.3 0.0010817 3.3 0.0010818 0 0.00108172 0 0.00108182 3.3 0.0010817399999999999 3.3 0.00108184 0 0.00108176 0 0.00108186 3.3 0.0010817799999999999 3.3 0.00108188 0 0.0010818 0 0.0010819 3.3 0.0010818199999999998 3.3 0.0010819199999999999 0 0.00108184 0 0.00108194 3.3 0.00108186 3.3 0.00108196 0 0.00108188 0 0.00108198 3.3 0.0010819 3.3 0.001082 0 0.0010819199999999999 0 0.00108202 3.3 0.00108194 3.3 0.00108204 0 0.0010819599999999999 0 0.00108206 3.3 0.00108198 3.3 0.00108208 0 0.0010819999999999998 0 0.0010821 3.3 0.00108202 3.3 0.00108212 0 0.0010820399999999998 0 0.0010821399999999999 3.3 0.00108206 3.3 0.00108216 0 0.00108208 0 0.00108218 3.3 0.0010821 3.3 0.0010822 0 0.00108212 0 0.00108222 3.3 0.0010821399999999999 3.3 0.00108224 0 0.00108216 0 0.00108226 3.3 0.0010821799999999999 3.3 0.00108228 0 0.0010822 0 0.0010823 3.3 0.0010822199999999998 3.3 0.00108232 0 0.00108224 0 0.00108234 3.3 0.0010822599999999998 3.3 0.0010823599999999999 0 0.00108228 0 0.00108238 3.3 0.0010823 3.3 0.0010824 0 0.00108232 0 0.00108242 3.3 0.00108234 3.3 0.00108244 0 0.0010823599999999999 0 0.00108246 3.3 0.00108238 3.3 0.00108248 0 0.0010823999999999999 0 0.0010825 3.3 0.00108242 3.3 0.00108252 0 0.0010824399999999998 0 0.0010825399999999999 3.3 0.00108246 3.3 0.00108256 0 0.0010824799999999998 0 0.0010825799999999999 3.3 0.0010825 3.3 0.0010826 0 0.00108252 0 0.00108262 3.3 0.0010825399999999999 3.3 0.00108264 0 0.00108256 0 0.00108266 3.3 0.0010825799999999999 3.3 0.00108268 0 0.0010826 0 0.0010827 3.3 0.0010826199999999998 3.3 0.00108272 0 0.00108264 0 0.00108274 3.3 0.0010826599999999998 3.3 0.0010827599999999999 0 0.00108268 0 0.00108278 3.3 0.0010827 3.3 0.0010828 0 0.00108272 0 0.00108282 3.3 0.00108274 3.3 0.00108284 0 0.0010827599999999999 0 0.00108286 3.3 0.00108278 3.3 0.00108288 0 0.0010827999999999999 0 0.0010829 3.3 0.00108282 3.3 0.00108292 0 0.0010828399999999998 0 0.00108294 3.3 0.00108286 3.3 0.00108296 0 0.0010828799999999998 0 0.0010829799999999999 3.3 0.0010829 3.3 0.001083 0 0.00108292 0 0.00108302 3.3 0.00108294 3.3 0.00108304 0 0.00108296 0 0.00108306 3.3 0.0010829799999999999 3.3 0.00108308 0 0.001083 0 0.0010831 3.3 0.0010830199999999999 3.3 0.00108312 0 0.00108304 0 0.00108314 3.3 0.0010830599999999998 3.3 0.00108316 0 0.00108308 0 0.00108318 3.3 0.0010830999999999998 3.3 0.0010831999999999999 0 0.00108312 0 0.00108322 3.3 0.00108314 3.3 0.00108324 0 0.00108316 0 0.00108326 3.3 0.00108318 3.3 0.00108328 0 0.0010831999999999999 0 0.0010833 3.3 0.00108322 3.3 0.00108332 0 0.0010832399999999999 0 0.00108334 3.3 0.00108326 3.3 0.00108336 0 0.0010832799999999998 0 0.0010833799999999999 3.3 0.0010833 3.3 0.0010834 0 0.00108332 0 0.00108342 3.3 0.00108334 3.3 0.00108344 0 0.00108336 0 0.00108346 3.3 0.0010833799999999999 3.3 0.00108348 0 0.0010834 0 0.0010835 3.3 0.0010834199999999999 3.3 0.00108352 0 0.00108344 0 0.00108354 3.3 0.0010834599999999998 3.3 0.00108356 0 0.00108348 0 0.00108358 3.3 0.0010834999999999998 3.3 0.0010835999999999999 0 0.00108352 0 0.00108362 3.3 0.00108354 3.3 0.00108364 0 0.00108356 0 0.00108366 3.3 0.00108358 3.3 0.00108368 0 0.0010835999999999999 0 0.0010837 3.3 0.00108362 3.3 0.00108372 0 0.0010836399999999999 0 0.00108374 3.3 0.00108366 3.3 0.00108376 0 0.0010836799999999998 0 0.00108378 3.3 0.0010837 3.3 0.0010838 0 0.0010837199999999998 0 0.0010838199999999999 3.3 0.00108374 3.3 0.00108384 0 0.00108376 0 0.00108386 3.3 0.00108378 3.3 0.00108388 0 0.0010838 0 0.0010839 3.3 0.0010838199999999999 3.3 0.00108392 0 0.00108384 0 0.00108394 3.3 0.0010838599999999999 3.3 0.00108396 0 0.00108388 0 0.00108398 3.3 0.0010838999999999998 3.3 0.001084 0 0.00108392 0 0.00108402 3.3 0.0010839399999999998 3.3 0.0010840399999999999 0 0.00108396 0 0.00108406 3.3 0.00108398 3.3 0.00108408 0 0.001084 0 0.0010841 3.3 0.00108402 3.3 0.00108412 0 0.0010840399999999999 0 0.00108414 3.3 0.00108406 3.3 0.00108416 0 0.0010840799999999999 0 0.00108418 3.3 0.0010841 3.3 0.0010842 0 0.0010841199999999998 0 0.0010842199999999999 3.3 0.00108414 3.3 0.00108424 0 0.00108416 0 0.00108426 3.3 0.00108418 3.3 0.00108428 0 0.0010842 0 0.0010843 3.3 0.0010842199999999999 3.3 0.00108432 0 0.00108424 0 0.00108434 3.3 0.0010842599999999999 3.3 0.00108436 0 0.00108428 0 0.00108438 3.3 0.0010842999999999998 3.3 0.0010844 0 0.00108432 0 0.00108442 3.3 0.0010843399999999998 3.3 0.0010844399999999999 0 0.00108436 0 0.00108446 3.3 0.00108438 3.3 0.00108448 0 0.0010844 0 0.0010845 3.3 0.00108442 3.3 0.00108452 0 0.0010844399999999999 0 0.00108454 3.3 0.00108446 3.3 0.00108456 0 0.0010844799999999999 0 0.00108458 3.3 0.0010845 3.3 0.0010846 0 0.0010845199999999998 0 0.00108462 3.3 0.00108454 3.3 0.00108464 0 0.0010845599999999998 0 0.0010846599999999999 3.3 0.00108458 3.3 0.00108468 0 0.0010846 0 0.0010847 3.3 0.00108462 3.3 0.00108472 0 0.00108464 0 0.00108474 3.3 0.0010846599999999999 3.3 0.00108476 0 0.00108468 0 0.00108478 3.3 0.0010846999999999999 3.3 0.0010848 0 0.00108472 0 0.00108482 3.3 0.0010847399999999998 3.3 0.00108484 0 0.00108476 0 0.00108486 3.3 0.0010847799999999998 3.3 0.0010848799999999999 0 0.0010848 0 0.0010849 3.3 0.00108482 3.3 0.00108492 0 0.00108484 0 0.00108494 3.3 0.00108486 3.3 0.00108496 0 0.0010848799999999999 0 0.00108498 3.3 0.0010849 3.3 0.001085 0 0.0010849199999999999 0 0.00108502 3.3 0.00108494 3.3 0.00108504 0 0.0010849599999999998 0 0.0010850599999999999 3.3 0.00108498 3.3 0.00108508 0 0.001085 0 0.0010851 3.3 0.00108502 3.3 0.00108512 0 0.00108504 0 0.00108514 3.3 0.0010850599999999999 3.3 0.00108516 0 0.00108508 0 0.00108518 3.3 0.0010850999999999999 3.3 0.0010852 0 0.00108512 0 0.00108522 3.3 0.0010851399999999998 3.3 0.00108524 0 0.00108516 0 0.00108526 3.3 0.0010851799999999998 3.3 0.0010852799999999999 0 0.0010852 0 0.0010853 3.3 0.00108522 3.3 0.00108532 0 0.00108524 0 0.00108534 3.3 0.00108526 3.3 0.00108536 0 0.0010852799999999999 0 0.00108538 3.3 0.0010853 3.3 0.0010854 0 0.0010853199999999999 0 0.00108542 3.3 0.00108534 3.3 0.00108544 0 0.0010853599999999998 0 0.00108546 3.3 0.00108538 3.3 0.00108548 0 0.0010853999999999998 0 0.0010854999999999999 3.3 0.00108542 3.3 0.00108552 0 0.00108544 0 0.00108554 3.3 0.00108546 3.3 0.00108556 0 0.00108548 0 0.00108558 3.3 0.0010854999999999999 3.3 0.0010856 0 0.00108552 0 0.00108562 3.3 0.0010855399999999999 3.3 0.00108564 0 0.00108556 0 0.00108566 3.3 0.0010855799999999998 3.3 0.00108568 0 0.0010856 0 0.0010857 3.3 0.0010856199999999998 3.3 0.0010857199999999999 0 0.00108564 0 0.00108574 3.3 0.00108566 3.3 0.00108576 0 0.00108568 0 0.00108578 3.3 0.0010857 3.3 0.0010858 0 0.0010857199999999999 0 0.00108582 3.3 0.00108574 3.3 0.00108584 0 0.0010857599999999999 0 0.00108586 3.3 0.00108578 3.3 0.00108588 0 0.0010857999999999998 0 0.0010858999999999999 3.3 0.00108582 3.3 0.00108592 0 0.00108584 0 0.00108594 3.3 0.00108586 3.3 0.00108596 0 0.00108588 0 0.00108598 3.3 0.0010858999999999999 3.3 0.001086 0 0.00108592 0 0.00108602 3.3 0.0010859399999999999 3.3 0.00108604 0 0.00108596 0 0.00108606 3.3 0.0010859799999999998 3.3 0.00108608 0 0.001086 0 0.0010861 3.3 0.0010860199999999998 3.3 0.0010861199999999999 0 0.00108604 0 0.00108614 3.3 0.00108606 3.3 0.00108616 0 0.00108608 0 0.00108618 3.3 0.0010861 3.3 0.0010862 0 0.0010861199999999999 0 0.00108622 3.3 0.00108614 3.3 0.00108624 0 0.0010861599999999999 0 0.00108626 3.3 0.00108618 3.3 0.00108628 0 0.0010861999999999998 0 0.0010863 3.3 0.00108622 3.3 0.00108632 0 0.0010862399999999998 0 0.0010863399999999999 3.3 0.00108626 3.3 0.00108636 0 0.00108628 0 0.00108638 3.3 0.0010863 3.3 0.0010864 0 0.00108632 0 0.00108642 3.3 0.0010863399999999999 3.3 0.00108644 0 0.00108636 0 0.00108646 3.3 0.0010863799999999999 3.3 0.00108648 0 0.0010864 0 0.0010865 3.3 0.0010864199999999998 3.3 0.0010865199999999999 0 0.00108644 0 0.00108654 3.3 0.00108646 3.3 0.00108656 0 0.00108648 0 0.00108658 3.3 0.0010865 3.3 0.0010866 0 0.0010865199999999999 0 0.00108662 3.3 0.00108654 3.3 0.00108664 0 0.0010865599999999999 0 0.00108666 3.3 0.00108658 3.3 0.00108668 0 0.0010865999999999998 0 0.0010867 3.3 0.00108662 3.3 0.00108672 0 0.0010866399999999998 0 0.0010867399999999999 3.3 0.00108666 3.3 0.00108676 0 0.00108668 0 0.00108678 3.3 0.0010867 3.3 0.0010868 0 0.00108672 0 0.00108682 3.3 0.0010867399999999999 3.3 0.00108684 0 0.00108676 0 0.00108686 3.3 0.0010867799999999999 3.3 0.00108688 0 0.0010868 0 0.0010869 3.3 0.0010868199999999998 3.3 0.00108692 0 0.00108684 0 0.00108694 3.3 0.0010868599999999998 3.3 0.0010869599999999999 0 0.00108688 0 0.00108698 3.3 0.0010869 3.3 0.001087 0 0.00108692 0 0.00108702 3.3 0.00108694 3.3 0.00108704 0 0.0010869599999999999 0 0.00108706 3.3 0.00108698 3.3 0.00108708 0 0.0010869999999999999 0 0.0010871 3.3 0.00108702 3.3 0.00108712 0 0.0010870399999999998 0 0.00108714 3.3 0.00108706 3.3 0.00108716 0 0.0010870799999999998 0 0.0010871799999999999 3.3 0.0010871 3.3 0.0010872 0 0.00108712 0 0.00108722 3.3 0.00108714 3.3 0.00108724 0 0.00108716 0 0.00108726 3.3 0.0010871799999999999 3.3 0.00108728 0 0.0010872 0 0.0010873 3.3 0.0010872199999999999 3.3 0.00108732 0 0.00108724 0 0.00108734 3.3 0.0010872599999999998 3.3 0.0010873599999999999 0 0.00108728 0 0.00108738 3.3 0.0010873 3.3 0.0010874 0 0.00108732 0 0.00108742 3.3 0.00108734 3.3 0.00108744 0 0.0010873599999999999 0 0.00108746 3.3 0.00108738 3.3 0.00108748 0 0.0010873999999999999 0 0.0010875 3.3 0.00108742 3.3 0.00108752 0 0.0010874399999999998 0 0.00108754 3.3 0.00108746 3.3 0.00108756 0 0.0010874799999999998 0 0.0010875799999999999 3.3 0.0010875 3.3 0.0010876 0 0.00108752 0 0.00108762 3.3 0.00108754 3.3 0.00108764 0 0.00108756 0 0.00108766 3.3 0.0010875799999999999 3.3 0.00108768 0 0.0010876 0 0.0010877 3.3 0.0010876199999999999 3.3 0.00108772 0 0.00108764 0 0.00108774 3.3 0.0010876599999999998 3.3 0.00108776 0 0.00108768 0 0.00108778 3.3 0.0010876999999999998 3.3 0.0010877999999999999 0 0.00108772 0 0.00108782 3.3 0.00108774 3.3 0.00108784 0 0.00108776 0 0.00108786 3.3 0.00108778 3.3 0.00108788 0 0.0010877999999999999 0 0.0010879 3.3 0.00108782 3.3 0.00108792 0 0.0010878399999999999 0 0.00108794 3.3 0.00108786 3.3 0.00108796 0 0.0010878799999999998 0 0.00108798 3.3 0.0010879 3.3 0.001088 0 0.0010879199999999998 0 0.0010880199999999999 3.3 0.00108794 3.3 0.00108804 0 0.00108796 0 0.00108806 3.3 0.00108798 3.3 0.00108808 0 0.001088 0 0.0010881 3.3 0.0010880199999999999 3.3 0.00108812 0 0.00108804 0 0.00108814 3.3 0.0010880599999999999 3.3 0.00108816 0 0.00108808 0 0.00108818 3.3 0.0010880999999999998 3.3 0.0010881999999999999 0 0.00108812 0 0.00108822 3.3 0.00108814 3.3 0.00108824 0 0.00108816 0 0.00108826 3.3 0.00108818 3.3 0.00108828 0 0.0010881999999999999 0 0.0010883 3.3 0.00108822 3.3 0.00108832 0 0.0010882399999999999 0 0.00108834 3.3 0.00108826 3.3 0.00108836 0 0.0010882799999999998 0 0.00108838 3.3 0.0010883 3.3 0.0010884 0 0.0010883199999999998 0 0.0010884199999999999 3.3 0.00108834 3.3 0.00108844 0 0.00108836 0 0.00108846 3.3 0.00108838 3.3 0.00108848 0 0.0010884 0 0.0010885 3.3 0.0010884199999999999 3.3 0.00108852 0 0.00108844 0 0.00108854 3.3 0.0010884599999999999 3.3 0.00108856 0 0.00108848 0 0.00108858 3.3 0.0010884999999999998 3.3 0.0010886 0 0.00108852 0 0.00108862 3.3 0.0010885399999999998 3.3 0.0010886399999999999 0 0.00108856 0 0.00108866 3.3 0.00108858 3.3 0.00108868 0 0.0010886 0 0.0010887 3.3 0.00108862 3.3 0.00108872 0 0.0010886399999999999 0 0.00108874 3.3 0.00108866 3.3 0.00108876 0 0.0010886799999999999 0 0.00108878 3.3 0.0010887 3.3 0.0010888 0 0.0010887199999999998 0 0.00108882 3.3 0.00108874 3.3 0.00108884 0 0.0010887599999999998 0 0.0010888599999999999 3.3 0.00108878 3.3 0.00108888 0 0.0010888 0 0.0010889 3.3 0.00108882 3.3 0.00108892 0 0.00108884 0 0.00108894 3.3 0.0010888599999999999 3.3 0.00108896 0 0.00108888 0 0.00108898 3.3 0.0010888999999999999 3.3 0.001089 0 0.00108892 0 0.00108902 3.3 0.0010889399999999998 3.3 0.0010890399999999999 0 0.00108896 0 0.00108906 3.3 0.00108898 3.3 0.00108908 0 0.001089 0 0.0010891 3.3 0.00108902 3.3 0.00108912 0 0.0010890399999999999 0 0.00108914 3.3 0.00108906 3.3 0.00108916 0 0.0010890799999999999 0 0.00108918 3.3 0.0010891 3.3 0.0010892 0 0.0010891199999999998 0 0.00108922 3.3 0.00108914 3.3 0.00108924 0 0.0010891599999999998 0 0.0010892599999999999 3.3 0.00108918 3.3 0.00108928 0 0.0010892 0 0.0010893 3.3 0.00108922 3.3 0.00108932 0 0.00108924 0 0.00108934 3.3 0.0010892599999999999 3.3 0.00108936 0 0.00108928 0 0.00108938 3.3 0.0010892999999999999 3.3 0.0010894 0 0.00108932 0 0.00108942 3.3 0.0010893399999999998 3.3 0.00108944 0 0.00108936 0 0.00108946 3.3 0.0010893799999999998 3.3 0.0010894799999999999 0 0.0010894 0 0.0010895 3.3 0.00108942 3.3 0.00108952 0 0.00108944 0 0.00108954 3.3 0.00108946 3.3 0.00108956 0 0.0010894799999999999 0 0.00108958 3.3 0.0010895 3.3 0.0010896 0 0.0010895199999999999 0 0.00108962 3.3 0.00108954 3.3 0.00108964 0 0.0010895599999999998 0 0.0010896599999999999 3.3 0.00108958 3.3 0.00108968 0 0.0010895999999999998 0 0.0010896999999999999 3.3 0.00108962 3.3 0.00108972 0 0.00108964 0 0.00108974 3.3 0.0010896599999999999 3.3 0.00108976 0 0.00108968 0 0.00108978 3.3 0.0010896999999999999 3.3 0.0010898 0 0.00108972 0 0.00108982 3.3 0.0010897399999999998 3.3 0.00108984 0 0.00108976 0 0.00108986 3.3 0.0010897799999999998 3.3 0.0010898799999999999 0 0.0010898 0 0.0010899 3.3 0.00108982 3.3 0.00108992 0 0.00108984 0 0.00108994 3.3 0.00108986 3.3 0.00108996 0 0.0010898799999999999 0 0.00108998 3.3 0.0010899 3.3 0.00109 0 0.0010899199999999999 0 0.00109002 3.3 0.00108994 3.3 0.00109004 0 0.0010899599999999998 0 0.00109006 3.3 0.00108998 3.3 0.00109008 0 0.0010899999999999998 0 0.0010900999999999999 3.3 0.00109002 3.3 0.00109012 0 0.00109004 0 0.00109014 3.3 0.00109006 3.3 0.00109016 0 0.00109008 0 0.00109018 3.3 0.0010900999999999999 3.3 0.0010902 0 0.00109012 0 0.00109022 3.3 0.0010901399999999999 3.3 0.00109024 0 0.00109016 0 0.00109026 3.3 0.0010901799999999998 3.3 0.00109028 0 0.0010902 0 0.0010903 3.3 0.0010902199999999998 3.3 0.0010903199999999999 0 0.00109024 0 0.00109034 3.3 0.00109026 3.3 0.00109036 0 0.00109028 0 0.00109038 3.3 0.0010903 3.3 0.0010904 0 0.0010903199999999999 0 0.00109042 3.3 0.00109034 3.3 0.00109044 0 0.0010903599999999999 0 0.00109046 3.3 0.00109038 3.3 0.00109048 0 0.0010903999999999998 0 0.0010904999999999999 3.3 0.00109042 3.3 0.00109052 0 0.00109044 0 0.00109054 3.3 0.00109046 3.3 0.00109056 0 0.00109048 0 0.00109058 3.3 0.0010904999999999999 3.3 0.0010906 0 0.00109052 0 0.00109062 3.3 0.0010905399999999999 3.3 0.00109064 0 0.00109056 0 0.00109066 3.3 0.0010905799999999998 3.3 0.00109068 0 0.0010906 0 0.0010907 3.3 0.0010906199999999998 3.3 0.0010907199999999999 0 0.00109064 0 0.00109074 3.3 0.00109066 3.3 0.00109076 0 0.00109068 0 0.00109078 3.3 0.0010907 3.3 0.0010908 0 0.0010907199999999999 0 0.00109082 3.3 0.00109074 3.3 0.00109084 0 0.0010907599999999999 0 0.00109086 3.3 0.00109078 3.3 0.00109088 0 0.0010907999999999998 0 0.0010909 3.3 0.00109082 3.3 0.00109092 0 0.0010908399999999998 0 0.0010909399999999999 3.3 0.00109086 3.3 0.00109096 0 0.00109088 0 0.00109098 3.3 0.0010909 3.3 0.001091 0 0.00109092 0 0.00109102 3.3 0.0010909399999999999 3.3 0.00109104 0 0.00109096 0 0.00109106 3.3 0.0010909799999999999 3.3 0.00109108 0 0.001091 0 0.0010911 3.3 0.0010910199999999998 3.3 0.00109112 0 0.00109104 0 0.00109114 3.3 0.0010910599999999998 3.3 0.0010911599999999999 0 0.00109108 0 0.00109118 3.3 0.0010911 3.3 0.0010912 0 0.00109112 0 0.00109122 3.3 0.00109114 3.3 0.00109124 0 0.0010911599999999999 0 0.00109126 3.3 0.00109118 3.3 0.00109128 0 0.0010911999999999999 0 0.0010913 3.3 0.00109122 3.3 0.00109132 0 0.0010912399999999998 0 0.0010913399999999999 3.3 0.00109126 3.3 0.00109136 0 0.00109128 0 0.00109138 3.3 0.0010913 3.3 0.0010914 0 0.00109132 0 0.00109142 3.3 0.0010913399999999999 3.3 0.00109144 0 0.00109136 0 0.00109146 3.3 0.0010913799999999999 3.3 0.00109148 0 0.0010914 0 0.0010915 3.3 0.0010914199999999998 3.3 0.00109152 0 0.00109144 0 0.00109154 3.3 0.0010914599999999998 3.3 0.0010915599999999999 0 0.00109148 0 0.00109158 3.3 0.0010915 3.3 0.0010916 0 0.00109152 0 0.00109162 3.3 0.00109154 3.3 0.00109164 0 0.0010915599999999999 0 0.00109166 3.3 0.00109158 3.3 0.00109168 0 0.0010915999999999999 0 0.0010917 3.3 0.00109162 3.3 0.00109172 0 0.0010916399999999998 0 0.00109174 3.3 0.00109166 3.3 0.00109176 0 0.0010916799999999998 0 0.0010917799999999999 3.3 0.0010917 3.3 0.0010918 0 0.00109172 0 0.00109182 3.3 0.00109174 3.3 0.00109184 0 0.00109176 0 0.00109186 3.3 0.0010917799999999999 3.3 0.00109188 0 0.0010918 0 0.0010919 3.3 0.0010918199999999999 3.3 0.00109192 0 0.00109184 0 0.00109194 3.3 0.0010918599999999998 3.3 0.00109196 0 0.00109188 0 0.00109198 3.3 0.0010918999999999998 3.3 0.0010919999999999999 0 0.00109192 0 0.00109202 3.3 0.00109194 3.3 0.00109204 0 0.00109196 0 0.00109206 3.3 0.00109198 3.3 0.00109208 0 0.0010919999999999999 0 0.0010921 3.3 0.00109202 3.3 0.00109212 0 0.0010920399999999999 0 0.00109214 3.3 0.00109206 3.3 0.00109216 0 0.0010920799999999998 0 0.0010921799999999999 3.3 0.0010921 3.3 0.0010922 0 0.00109212 0 0.00109222 3.3 0.00109214 3.3 0.00109224 0 0.00109216 0 0.00109226 3.3 0.0010921799999999999 3.3 0.00109228 0 0.0010922 0 0.0010923 3.3 0.0010922199999999999 3.3 0.00109232 0 0.00109224 0 0.00109234 3.3 0.0010922599999999998 3.3 0.00109236 0 0.00109228 0 0.00109238 3.3 0.0010922999999999998 3.3 0.0010923999999999999 0 0.00109232 0 0.00109242 3.3 0.00109234 3.3 0.00109244 0 0.00109236 0 0.00109246 3.3 0.00109238 3.3 0.00109248 0 0.0010923999999999999 0 0.0010925 3.3 0.00109242 3.3 0.00109252 0 0.0010924399999999999 0 0.00109254 3.3 0.00109246 3.3 0.00109256 0 0.0010924799999999998 0 0.00109258 3.3 0.0010925 3.3 0.0010926 0 0.0010925199999999998 0 0.0010926199999999999 3.3 0.00109254 3.3 0.00109264 0 0.00109256 0 0.00109266 3.3 0.00109258 3.3 0.00109268 0 0.0010926 0 0.0010927 3.3 0.0010926199999999999 3.3 0.00109272 0 0.00109264 0 0.00109274 3.3 0.0010926599999999999 3.3 0.00109276 0 0.00109268 0 0.00109278 3.3 0.0010926999999999998 3.3 0.0010927999999999999 0 0.00109272 0 0.00109282 3.3 0.0010927399999999998 3.3 0.0010928399999999999 0 0.00109276 0 0.00109286 3.3 0.00109278 3.3 0.00109288 0 0.0010927999999999999 0 0.0010929 3.3 0.00109282 3.3 0.00109292 0 0.0010928399999999999 0 0.00109294 3.3 0.00109286 3.3 0.00109296 0 0.0010928799999999998 0 0.00109298 3.3 0.0010929 3.3 0.001093 0 0.0010929199999999998 0 0.0010930199999999999 3.3 0.00109294 3.3 0.00109304 0 0.00109296 0 0.00109306 3.3 0.00109298 3.3 0.00109308 0 0.001093 0 0.0010931 3.3 0.0010930199999999999 3.3 0.00109312 0 0.00109304 0 0.00109314 3.3 0.0010930599999999999 3.3 0.00109316 0 0.00109308 0 0.00109318 3.3 0.0010930999999999998 3.3 0.0010932 0 0.00109312 0 0.00109322 3.3 0.0010931399999999998 3.3 0.0010932399999999999 0 0.00109316 0 0.00109326 3.3 0.00109318 3.3 0.00109328 0 0.0010932 0 0.0010933 3.3 0.00109322 3.3 0.00109332 0 0.0010932399999999999 0 0.00109334 3.3 0.00109326 3.3 0.00109336 0 0.0010932799999999999 0 0.00109338 3.3 0.0010933 3.3 0.0010934 0 0.0010933199999999998 0 0.00109342 3.3 0.00109334 3.3 0.00109344 0 0.0010933599999999998 0 0.0010934599999999999 3.3 0.00109338 3.3 0.00109348 0 0.0010934 0 0.0010935 3.3 0.00109342 3.3 0.00109352 0 0.00109344 0 0.00109354 3.3 0.0010934599999999999 3.3 0.00109356 0 0.00109348 0 0.00109358 3.3 0.0010934999999999999 3.3 0.0010936 0 0.00109352 0 0.00109362 3.3 0.0010935399999999998 3.3 0.0010936399999999999 0 0.00109356 0 0.00109366 3.3 0.00109358 3.3 0.00109368 0 0.0010936 0 0.0010937 3.3 0.00109362 3.3 0.00109372 0 0.0010936399999999999 0 0.00109374 3.3 0.00109366 3.3 0.00109376 0 0.0010936799999999999 0 0.00109378 3.3 0.0010937 3.3 0.0010938 0 0.0010937199999999998 0 0.00109382 3.3 0.00109374 3.3 0.00109384 0 0.0010937599999999998 0 0.0010938599999999999 3.3 0.00109378 3.3 0.00109388 0 0.0010938 0 0.0010939 3.3 0.00109382 3.3 0.00109392 0 0.00109384 0 0.00109394 3.3 0.0010938599999999999 3.3 0.00109396 0 0.00109388 0 0.00109398 3.3 0.0010938999999999999 3.3 0.001094 0 0.00109392 0 0.00109402 3.3 0.0010939399999999998 3.3 0.00109404 0 0.00109396 0 0.00109406 3.3 0.0010939799999999998 3.3 0.0010940799999999999 0 0.001094 0 0.0010941 3.3 0.00109402 3.3 0.00109412 0 0.00109404 0 0.00109414 3.3 0.00109406 3.3 0.00109416 0 0.0010940799999999999 0 0.00109418 3.3 0.0010941 3.3 0.0010942 0 0.0010941199999999999 0 0.00109422 3.3 0.00109414 3.3 0.00109424 0 0.0010941599999999998 0 0.00109426 3.3 0.00109418 3.3 0.00109428 0 0.0010941999999999998 0 0.0010942999999999999 3.3 0.00109422 3.3 0.00109432 0 0.00109424 0 0.00109434 3.3 0.00109426 3.3 0.00109436 0 0.00109428 0 0.00109438 3.3 0.0010942999999999999 3.3 0.0010944 0 0.00109432 0 0.00109442 3.3 0.0010943399999999999 3.3 0.00109444 0 0.00109436 0 0.00109446 3.3 0.0010943799999999998 3.3 0.0010944799999999999 0 0.0010944 0 0.0010945 3.3 0.00109442 3.3 0.00109452 0 0.00109444 0 0.00109454 3.3 0.00109446 3.3 0.00109456 0 0.0010944799999999999 0 0.00109458 3.3 0.0010945 3.3 0.0010946 0 0.0010945199999999999 0 0.00109462 3.3 0.00109454 3.3 0.00109464 0 0.0010945599999999998 0 0.00109466 3.3 0.00109458 3.3 0.00109468 0 0.0010945999999999998 0 0.0010946999999999999 3.3 0.00109462 3.3 0.00109472 0 0.00109464 0 0.00109474 3.3 0.00109466 3.3 0.00109476 0 0.00109468 0 0.00109478 3.3 0.0010946999999999999 3.3 0.0010948 0 0.00109472 0 0.00109482 3.3 0.0010947399999999999 3.3 0.00109484 0 0.00109476 0 0.00109486 3.3 0.0010947799999999998 3.3 0.00109488 0 0.0010948 0 0.0010949 3.3 0.0010948199999999998 3.3 0.0010949199999999999 0 0.00109484 0 0.00109494 3.3 0.00109486 3.3 0.00109496 0 0.00109488 0 0.00109498 3.3 0.0010949 3.3 0.001095 0 0.0010949199999999999 0 0.00109502 3.3 0.00109494 3.3 0.00109504 0 0.0010949599999999999 0 0.00109506 3.3 0.00109498 3.3 0.00109508 0 0.0010949999999999998 0 0.0010951 3.3 0.00109502 3.3 0.00109512 0 0.0010950399999999998 0 0.0010951399999999999 3.3 0.00109506 3.3 0.00109516 0 0.00109508 0 0.00109518 3.3 0.0010951 3.3 0.0010952 0 0.00109512 0 0.00109522 3.3 0.0010951399999999999 3.3 0.00109524 0 0.00109516 0 0.00109526 3.3 0.0010951799999999999 3.3 0.00109528 0 0.0010952 0 0.0010953 3.3 0.0010952199999999998 3.3 0.0010953199999999999 0 0.00109524 0 0.00109534 3.3 0.00109526 3.3 0.00109536 0 0.00109528 0 0.00109538 3.3 0.0010953 3.3 0.0010954 0 0.0010953199999999999 0 0.00109542 3.3 0.00109534 3.3 0.00109544 0 0.0010953599999999999 0 0.00109546 3.3 0.00109538 3.3 0.00109548 0 0.0010953999999999998 0 0.0010955 3.3 0.00109542 3.3 0.00109552 0 0.0010954399999999998 0 0.0010955399999999999 3.3 0.00109546 3.3 0.00109556 0 0.00109548 0 0.00109558 3.3 0.0010955 3.3 0.0010956 0 0.00109552 0 0.00109562 3.3 0.0010955399999999999 3.3 0.00109564 0 0.00109556 0 0.00109566 3.3 0.0010955799999999999 3.3 0.00109568 0 0.0010956 0 0.0010957 3.3 0.0010956199999999998 3.3 0.00109572 0 0.00109564 0 0.00109574 3.3 0.0010956599999999998 3.3 0.0010957599999999999 0 0.00109568 0 0.00109578 3.3 0.0010957 3.3 0.0010958 0 0.00109572 0 0.00109582 3.3 0.00109574 3.3 0.00109584 0 0.0010957599999999999 0 0.00109586 3.3 0.00109578 3.3 0.00109588 0 0.0010957999999999999 0 0.0010959 3.3 0.00109582 3.3 0.00109592 0 0.0010958399999999998 0 0.00109594 3.3 0.00109586 3.3 0.00109596 0 0.0010958799999999998 0 0.0010959799999999999 3.3 0.0010959 3.3 0.001096 0 0.00109592 0 0.00109602 3.3 0.00109594 3.3 0.00109604 0 0.00109596 0 0.00109606 3.3 0.0010959799999999999 3.3 0.00109608 0 0.001096 0 0.0010961 3.3 0.0010960199999999999 3.3 0.00109612 0 0.00109604 0 0.00109614 3.3 0.0010960599999999998 3.3 0.0010961599999999999 0 0.00109608 0 0.00109618 3.3 0.0010961 3.3 0.0010962 0 0.00109612 0 0.00109622 3.3 0.00109614 3.3 0.00109624 0 0.0010961599999999999 0 0.00109626 3.3 0.00109618 3.3 0.00109628 0 0.0010961999999999999 0 0.0010963 3.3 0.00109622 3.3 0.00109632 0 0.0010962399999999998 0 0.00109634 3.3 0.00109626 3.3 0.00109636 0 0.0010962799999999998 0 0.0010963799999999999 3.3 0.0010963 3.3 0.0010964 0 0.00109632 0 0.00109642 3.3 0.00109634 3.3 0.00109644 0 0.00109636 0 0.00109646 3.3 0.0010963799999999999 3.3 0.00109648 0 0.0010964 0 0.0010965 3.3 0.0010964199999999999 3.3 0.00109652 0 0.00109644 0 0.00109654 3.3 0.0010964599999999998 3.3 0.00109656 0 0.00109648 0 0.00109658 3.3 0.0010964999999999998 3.3 0.0010965999999999999 0 0.00109652 0 0.00109662 3.3 0.00109654 3.3 0.00109664 0 0.00109656 0 0.00109666 3.3 0.00109658 3.3 0.00109668 0 0.0010965999999999999 0 0.0010967 3.3 0.00109662 3.3 0.00109672 0 0.0010966399999999999 0 0.00109674 3.3 0.00109666 3.3 0.00109676 0 0.0010966799999999998 0 0.0010967799999999999 3.3 0.0010967 3.3 0.0010968 0 0.0010967199999999998 0 0.0010968199999999999 3.3 0.00109674 3.3 0.00109684 0 0.00109676 0 0.00109686 3.3 0.0010967799999999999 3.3 0.00109688 0 0.0010968 0 0.0010969 3.3 0.0010968199999999999 3.3 0.00109692 0 0.00109684 0 0.00109694 3.3 0.0010968599999999998 3.3 0.00109696 0 0.00109688 0 0.00109698 3.3 0.0010968999999999998 3.3 0.0010969999999999999 0 0.00109692 0 0.00109702 3.3 0.00109694 3.3 0.00109704 0 0.00109696 0 0.00109706 3.3 0.00109698 3.3 0.00109708 0 0.0010969999999999999 0 0.0010971 3.3 0.00109702 3.3 0.00109712 0 0.0010970399999999999 0 0.00109714 3.3 0.00109706 3.3 0.00109716 0 0.0010970799999999998 0 0.00109718 3.3 0.0010971 3.3 0.0010972 0 0.0010971199999999998 0 0.0010972199999999999 3.3 0.00109714 3.3 0.00109724 0 0.00109716 0 0.00109726 3.3 0.00109718 3.3 0.00109728 0 0.0010972 0 0.0010973 3.3 0.0010972199999999999 3.3 0.00109732 0 0.00109724 0 0.00109734 3.3 0.0010972599999999999 3.3 0.00109736 0 0.00109728 0 0.00109738 3.3 0.0010972999999999998 3.3 0.0010974 0 0.00109732 0 0.00109742 3.3 0.0010973399999999998 3.3 0.0010974399999999999 0 0.00109736 0 0.00109746 3.3 0.00109738 3.3 0.00109748 0 0.0010974 0 0.0010975 3.3 0.00109742 3.3 0.00109752 0 0.0010974399999999999 0 0.00109754 3.3 0.00109746 3.3 0.00109756 0 0.0010974799999999999 0 0.00109758 3.3 0.0010975 3.3 0.0010976 0 0.0010975199999999998 0 0.0010976199999999999 3.3 0.00109754 3.3 0.00109764 0 0.00109756 0 0.00109766 3.3 0.00109758 3.3 0.00109768 0 0.0010976 0 0.0010977 3.3 0.0010976199999999999 3.3 0.00109772 0 0.00109764 0 0.00109774 3.3 0.0010976599999999999 3.3 0.00109776 0 0.00109768 0 0.00109778 3.3 0.0010976999999999998 3.3 0.0010978 0 0.00109772 0 0.00109782 3.3 0.0010977399999999998 3.3 0.0010978399999999999 0 0.00109776 0 0.00109786 3.3 0.00109778 3.3 0.00109788 0 0.0010978 0 0.0010979 3.3 0.00109782 3.3 0.00109792 0 0.0010978399999999999 0 0.00109794 3.3 0.00109786 3.3 0.00109796 0 0.0010978799999999999 0 0.00109798 3.3 0.0010979 3.3 0.001098 0 0.0010979199999999998 0 0.00109802 3.3 0.00109794 3.3 0.00109804 0 0.0010979599999999998 0 0.0010980599999999999 3.3 0.00109798 3.3 0.00109808 0 0.001098 0 0.0010981 3.3 0.00109802 3.3 0.00109812 0 0.00109804 0 0.00109814 3.3 0.0010980599999999999 3.3 0.00109816 0 0.00109808 0 0.00109818 3.3 0.0010980999999999999 3.3 0.0010982 0 0.00109812 0 0.00109822 3.3 0.0010981399999999998 3.3 0.00109824 0 0.00109816 0 0.00109826 3.3 0.0010981799999999998 3.3 0.0010982799999999999 0 0.0010982 0 0.0010983 3.3 0.00109822 3.3 0.00109832 0 0.00109824 0 0.00109834 3.3 0.00109826 3.3 0.00109836 0 0.0010982799999999999 0 0.00109838 3.3 0.0010983 3.3 0.0010984 0 0.0010983199999999999 0 0.00109842 3.3 0.00109834 3.3 0.00109844 0 0.0010983599999999998 0 0.0010984599999999999 3.3 0.00109838 3.3 0.00109848 0 0.0010984 0 0.0010985 3.3 0.00109842 3.3 0.00109852 0 0.00109844 0 0.00109854 3.3 0.0010984599999999999 3.3 0.00109856 0 0.00109848 0 0.00109858 3.3 0.0010984999999999999 3.3 0.0010986 0 0.00109852 0 0.00109862 3.3 0.0010985399999999998 3.3 0.00109864 0 0.00109856 0 0.00109866 3.3 0.0010985799999999998 3.3 0.0010986799999999999 0 0.0010986 0 0.0010987 3.3 0.00109862 3.3 0.00109872 0 0.00109864 0 0.00109874 3.3 0.00109866 3.3 0.00109876 0 0.0010986799999999999 0 0.00109878 3.3 0.0010987 3.3 0.0010988 0 0.0010987199999999999 0 0.00109882 3.3 0.00109874 3.3 0.00109884 0 0.0010987599999999998 0 0.00109886 3.3 0.00109878 3.3 0.00109888 0 0.0010987999999999998 0 0.0010988999999999999 3.3 0.00109882 3.3 0.00109892 0 0.00109884 0 0.00109894 3.3 0.00109886 3.3 0.00109896 0 0.00109888 0 0.00109898 3.3 0.0010988999999999999 3.3 0.001099 0 0.00109892 0 0.00109902 3.3 0.0010989399999999999 3.3 0.00109904 0 0.00109896 0 0.00109906 3.3 0.0010989799999999998 3.3 0.00109908 0 0.001099 0 0.0010991 3.3 0.0010990199999999998 3.3 0.0010991199999999999 0 0.00109904 0 0.00109914 3.3 0.00109906 3.3 0.00109916 0 0.00109908 0 0.00109918 3.3 0.0010991 3.3 0.0010992 0 0.0010991199999999999 0 0.00109922 3.3 0.00109914 3.3 0.00109924 0 0.0010991599999999999 0 0.00109926 3.3 0.00109918 3.3 0.00109928 0 0.0010991999999999998 0 0.0010992999999999999 3.3 0.00109922 3.3 0.00109932 0 0.00109924 0 0.00109934 3.3 0.00109926 3.3 0.00109936 0 0.00109928 0 0.00109938 3.3 0.0010992999999999999 3.3 0.0010994 0 0.00109932 0 0.00109942 3.3 0.0010993399999999999 3.3 0.00109944 0 0.00109936 0 0.00109946 3.3 0.0010993799999999998 3.3 0.00109948 0 0.0010994 0 0.0010995 3.3 0.0010994199999999998 3.3 0.0010995199999999999 0 0.00109944 0 0.00109954 3.3 0.00109946 3.3 0.00109956 0 0.00109948 0 0.00109958 3.3 0.0010995 3.3 0.0010996 0 0.0010995199999999999 0 0.00109962 3.3 0.00109954 3.3 0.00109964 0 0.0010995599999999999 0 0.00109966 3.3 0.00109958 3.3 0.00109968 0 0.0010995999999999998 0 0.0010997 3.3 0.00109962 3.3 0.00109972 0 0.0010996399999999998 0 0.0010997399999999999 3.3 0.00109966 3.3 0.00109976 0 0.00109968 0 0.00109978 3.3 0.0010997 3.3 0.0010998 0 0.00109972 0 0.00109982 3.3 0.0010997399999999999 3.3 0.00109984 0 0.00109976 0 0.00109986 3.3 0.0010997799999999999 3.3 0.00109988 0 0.0010998 0 0.0010999 3.3 0.0010998199999999998 3.3 0.0010999199999999999 0 0.00109984 0 0.00109994 3.3 0.0010998599999999998 3.3 0.0010999599999999999 0 0.00109988 0 0.00109998 3.3 0.0010999 3.3 0.0011 0 0.0010999199999999999 0 0.00110002 3.3 0.00109994 3.3 0.00110004 0 0.0010999599999999999 0 0.00110006 3.3 0.00109998 3.3 0.00110008 0 0.0010999999999999998 0 0.0011001 3.3 0.00110002 3.3 0.00110012 0 0.0011000399999999998 0 0.0011001399999999999 3.3 0.00110006 3.3 0.00110016 0 0.00110008 0 0.00110018 3.3 0.0011001 3.3 0.0011002 0 0.00110012 0 0.00110022 3.3 0.0011001399999999999 3.3 0.00110024 0 0.00110016 0 0.00110026 3.3 0.0011001799999999999 3.3 0.00110028 0 0.0011002 0 0.0011003 3.3 0.0011002199999999998 3.3 0.00110032 0 0.00110024 0 0.00110034 3.3 0.0011002599999999998 3.3 0.0011003599999999999 0 0.00110028 0 0.00110038 3.3 0.0011003 3.3 0.0011004 0 0.00110032 0 0.00110042 3.3 0.00110034 3.3 0.00110044 0 0.0011003599999999999 0 0.00110046 3.3 0.00110038 3.3 0.00110048 0 0.0011003999999999999 0 0.0011005 3.3 0.00110042 3.3 0.00110052 0 0.0011004399999999998 0 0.00110054 3.3 0.00110046 3.3 0.00110056 0 0.0011004799999999998 0 0.0011005799999999999 3.3 0.0011005 3.3 0.0011006 0 0.00110052 0 0.00110062 3.3 0.00110054 3.3 0.00110064 0 0.00110056 0 0.00110066 3.3 0.0011005799999999999 3.3 0.00110068 0 0.0011006 0 0.0011007 3.3 0.0011006199999999999 3.3 0.00110072 0 0.00110064 0 0.00110074 3.3 0.0011006599999999998 3.3 0.0011007599999999999 0 0.00110068 0 0.00110078 3.3 0.0011007 3.3 0.0011008 0 0.00110072 0 0.00110082 3.3 0.00110074 3.3 0.00110084 0 0.0011007599999999999 0 0.00110086 3.3 0.00110078 3.3 0.00110088 0 0.0011007999999999999 0 0.0011009 3.3 0.00110082 3.3 0.00110092 0 0.0011008399999999998 0 0.00110094 3.3 0.00110086 3.3 0.00110096 0 0.0011008799999999998 0 0.0011009799999999999 3.3 0.0011009 3.3 0.001101 0 0.00110092 0 0.00110102 3.3 0.00110094 3.3 0.00110104 0 0.00110096 0 0.00110106 3.3 0.0011009799999999999 3.3 0.00110108 0 0.001101 0 0.0011011 3.3 0.0011010199999999999 3.3 0.00110112 0 0.00110104 0 0.00110114 3.3 0.0011010599999999998 3.3 0.00110116 0 0.00110108 0 0.00110118 3.3 0.0011010999999999998 3.3 0.0011011999999999999 0 0.00110112 0 0.00110122 3.3 0.00110114 3.3 0.00110124 0 0.00110116 0 0.00110126 3.3 0.00110118 3.3 0.00110128 0 0.0011011999999999999 0 0.0011013 3.3 0.00110122 3.3 0.00110132 0 0.0011012399999999999 0 0.00110134 3.3 0.00110126 3.3 0.00110136 0 0.0011012799999999998 0 0.00110138 3.3 0.0011013 3.3 0.0011014 0 0.0011013199999999998 0 0.0011014199999999999 3.3 0.00110134 3.3 0.00110144 0 0.00110136 0 0.00110146 3.3 0.00110138 3.3 0.00110148 0 0.0011014 0 0.0011015 3.3 0.0011014199999999999 3.3 0.00110152 0 0.00110144 0 0.00110154 3.3 0.0011014599999999999 3.3 0.00110156 0 0.00110148 0 0.00110158 3.3 0.0011014999999999998 3.3 0.0011015999999999999 0 0.00110152 0 0.00110162 3.3 0.00110154 3.3 0.00110164 0 0.00110156 0 0.00110166 3.3 0.00110158 3.3 0.00110168 0 0.0011015999999999999 0 0.0011017 3.3 0.00110162 3.3 0.00110172 0 0.0011016399999999999 0 0.00110174 3.3 0.00110166 3.3 0.00110176 0 0.0011016799999999998 0 0.00110178 3.3 0.0011017 3.3 0.0011018 0 0.0011017199999999998 0 0.0011018199999999999 3.3 0.00110174 3.3 0.00110184 0 0.00110176 0 0.00110186 3.3 0.00110178 3.3 0.00110188 0 0.0011018 0 0.0011019 3.3 0.0011018199999999999 3.3 0.00110192 0 0.00110184 0 0.00110194 3.3 0.0011018599999999999 3.3 0.00110196 0 0.00110188 0 0.00110198 3.3 0.0011018999999999998 3.3 0.001102 0 0.00110192 0 0.00110202 3.3 0.0011019399999999998 3.3 0.0011020399999999999 0 0.00110196 0 0.00110206 3.3 0.00110198 3.3 0.00110208 0 0.001102 0 0.0011021 3.3 0.00110202 3.3 0.00110212 0 0.0011020399999999999 0 0.00110214 3.3 0.00110206 3.3 0.00110216 0 0.0011020799999999999 0 0.00110218 3.3 0.0011021 3.3 0.0011022 0 0.0011021199999999998 0 0.00110222 3.3 0.00110214 3.3 0.00110224 0 0.0011021599999999998 0 0.0011022599999999999 3.3 0.00110218 3.3 0.00110228 0 0.0011022 0 0.0011023 3.3 0.00110222 3.3 0.00110232 0 0.00110224 0 0.00110234 3.3 0.0011022599999999999 3.3 0.00110236 0 0.00110228 0 0.00110238 3.3 0.0011022999999999999 3.3 0.0011024 0 0.00110232 0 0.00110242 3.3 0.0011023399999999998 3.3 0.0011024399999999999 0 0.00110236 0 0.00110246 3.3 0.00110238 3.3 0.00110248 0 0.0011024 0 0.0011025 3.3 0.00110242 3.3 0.00110252 0 0.0011024399999999999 0 0.00110254 3.3 0.00110246 3.3 0.00110256 0 0.0011024799999999999 0 0.00110258 3.3 0.0011025 3.3 0.0011026 0 0.0011025199999999998 0 0.00110262 3.3 0.00110254 3.3 0.00110264 0 0.0011025599999999998 0 0.0011026599999999999 3.3 0.00110258 3.3 0.00110268 0 0.0011026 0 0.0011027 3.3 0.00110262 3.3 0.00110272 0 0.00110264 0 0.00110274 3.3 0.0011026599999999999 3.3 0.00110276 0 0.00110268 0 0.00110278 3.3 0.0011026999999999999 3.3 0.0011028 0 0.00110272 0 0.00110282 3.3 0.0011027399999999998 3.3 0.00110284 0 0.00110276 0 0.00110286 3.3 0.0011027799999999998 3.3 0.0011028799999999999 0 0.0011028 0 0.0011029 3.3 0.00110282 3.3 0.00110292 0 0.00110284 0 0.00110294 3.3 0.00110286 3.3 0.00110296 0 0.0011028799999999999 0 0.00110298 3.3 0.0011029 3.3 0.001103 0 0.0011029199999999999 0 0.00110302 3.3 0.00110294 3.3 0.00110304 0 0.0011029599999999998 0 0.0011030599999999999 3.3 0.00110298 3.3 0.00110308 0 0.0011029999999999998 0 0.0011030999999999999 3.3 0.00110302 3.3 0.00110312 0 0.00110304 0 0.00110314 3.3 0.0011030599999999999 3.3 0.00110316 0 0.00110308 0 0.00110318 3.3 0.0011030999999999999 3.3 0.0011032 0 0.00110312 0 0.00110322 3.3 0.0011031399999999998 3.3 0.00110324 0 0.00110316 0 0.00110326 3.3 0.0011031799999999998 3.3 0.0011032799999999999 0 0.0011032 0 0.0011033 3.3 0.00110322 3.3 0.00110332 0 0.00110324 0 0.00110334 3.3 0.00110326 3.3 0.00110336 0 0.0011032799999999999 0 0.00110338 3.3 0.0011033 3.3 0.0011034 0 0.0011033199999999999 0 0.00110342 3.3 0.00110334 3.3 0.00110344 0 0.0011033599999999998 0 0.00110346 3.3 0.00110338 3.3 0.00110348 0 0.0011033999999999998 0 0.0011034999999999999 3.3 0.00110342 3.3 0.00110352 0 0.00110344 0 0.00110354 3.3 0.00110346 3.3 0.00110356 0 0.00110348 0 0.00110358 3.3 0.0011034999999999999 3.3 0.0011036 0 0.00110352 0 0.00110362 3.3 0.0011035399999999999 3.3 0.00110364 0 0.00110356 0 0.00110366 3.3 0.0011035799999999998 3.3 0.00110368 0 0.0011036 0 0.0011037 3.3 0.0011036199999999998 3.3 0.0011037199999999999 0 0.00110364 0 0.00110374 3.3 0.00110366 3.3 0.00110376 0 0.00110368 0 0.00110378 3.3 0.0011037 3.3 0.0011038 0 0.0011037199999999999 0 0.00110382 3.3 0.00110374 3.3 0.00110384 0 0.0011037599999999999 0 0.00110386 3.3 0.00110378 3.3 0.00110388 0 0.0011037999999999998 0 0.0011038999999999999 3.3 0.00110382 3.3 0.00110392 0 0.00110384 0 0.00110394 3.3 0.00110386 3.3 0.00110396 0 0.00110388 0 0.00110398 3.3 0.0011038999999999999 3.3 0.001104 0 0.00110392 0 0.00110402 3.3 0.0011039399999999999 3.3 0.00110404 0 0.00110396 0 0.00110406 3.3 0.0011039799999999998 3.3 0.00110408 0 0.001104 0 0.0011041 3.3 0.0011040199999999998 3.3 0.0011041199999999999 0 0.00110404 0 0.00110414 3.3 0.00110406 3.3 0.00110416 0 0.00110408 0 0.00110418 3.3 0.0011041 3.3 0.0011042 0 0.0011041199999999999 0 0.00110422 3.3 0.00110414 3.3 0.00110424 0 0.0011041599999999999 0 0.00110426 3.3 0.00110418 3.3 0.00110428 0 0.0011041999999999998 0 0.0011043 3.3 0.00110422 3.3 0.00110432 0 0.0011042399999999998 0 0.0011043399999999999 3.3 0.00110426 3.3 0.00110436 0 0.00110428 0 0.00110438 3.3 0.0011043 3.3 0.0011044 0 0.00110432 0 0.00110442 3.3 0.0011043399999999999 3.3 0.00110444 0 0.00110436 0 0.00110446 3.3 0.0011043799999999999 3.3 0.00110448 0 0.0011044 0 0.0011045 3.3 0.0011044199999999998 3.3 0.00110452 0 0.00110444 0 0.00110454 3.3 0.0011044599999999998 3.3 0.0011045599999999999 0 0.00110448 0 0.00110458 3.3 0.0011045 3.3 0.0011046 0 0.00110452 0 0.00110462 3.3 0.00110454 3.3 0.00110464 0 0.0011045599999999999 0 0.00110466 3.3 0.00110458 3.3 0.00110468 0 0.0011045999999999999 0 0.0011047 3.3 0.00110462 3.3 0.00110472 0 0.0011046399999999998 0 0.0011047399999999999 3.3 0.00110466 3.3 0.00110476 0 0.00110468 0 0.00110478 3.3 0.0011047 3.3 0.0011048 0 0.00110472 0 0.00110482 3.3 0.0011047399999999999 3.3 0.00110484 0 0.00110476 0 0.00110486 3.3 0.0011047799999999999 3.3 0.00110488 0 0.0011048 0 0.0011049 3.3 0.0011048199999999998 3.3 0.00110492 0 0.00110484 0 0.00110494 3.3 0.0011048599999999998 3.3 0.0011049599999999999 0 0.00110488 0 0.00110498 3.3 0.0011049 3.3 0.001105 0 0.00110492 0 0.00110502 3.3 0.00110494 3.3 0.00110504 0 0.0011049599999999999 0 0.00110506 3.3 0.00110498 3.3 0.00110508 0 0.0011049999999999999 0 0.0011051 3.3 0.00110502 3.3 0.00110512 0 0.0011050399999999998 0 0.00110514 3.3 0.00110506 3.3 0.00110516 0 0.0011050799999999998 0 0.0011051799999999999 3.3 0.0011051 3.3 0.0011052 0 0.00110512 0 0.00110522 3.3 0.00110514 3.3 0.00110524 0 0.00110516 0 0.00110526 3.3 0.0011051799999999999 3.3 0.00110528 0 0.0011052 0 0.0011053 3.3 0.0011052199999999999 3.3 0.00110532 0 0.00110524 0 0.00110534 3.3 0.0011052599999999998 3.3 0.00110536 0 0.00110528 0 0.00110538 3.3 0.0011052999999999998 3.3 0.0011053999999999999 0 0.00110532 0 0.00110542 3.3 0.00110534 3.3 0.00110544 0 0.00110536 0 0.00110546 3.3 0.00110538 3.3 0.00110548 0 0.0011053999999999999 0 0.0011055 3.3 0.00110542 3.3 0.00110552 0 0.0011054399999999999 0 0.00110554 3.3 0.00110546 3.3 0.00110556 0 0.0011054799999999998 0 0.0011055799999999999 3.3 0.0011055 3.3 0.0011056 0 0.00110552 0 0.00110562 3.3 0.00110554 3.3 0.00110564 0 0.00110556 0 0.00110566 3.3 0.0011055799999999999 3.3 0.00110568 0 0.0011056 0 0.0011057 3.3 0.0011056199999999999 3.3 0.00110572 0 0.00110564 0 0.00110574 3.3 0.0011056599999999998 3.3 0.00110576 0 0.00110568 0 0.00110578 3.3 0.0011056999999999998 3.3 0.0011057999999999999 0 0.00110572 0 0.00110582 3.3 0.00110574 3.3 0.00110584 0 0.00110576 0 0.00110586 3.3 0.00110578 3.3 0.00110588 0 0.0011057999999999999 0 0.0011059 3.3 0.00110582 3.3 0.00110592 0 0.0011058399999999999 0 0.00110594 3.3 0.00110586 3.3 0.00110596 0 0.0011058799999999998 0 0.00110598 3.3 0.0011059 3.3 0.001106 0 0.0011059199999999998 0 0.0011060199999999999 3.3 0.00110594 3.3 0.00110604 0 0.00110596 0 0.00110606 3.3 0.00110598 3.3 0.00110608 0 0.001106 0 0.0011061 3.3 0.0011060199999999999 3.3 0.00110612 0 0.00110604 0 0.00110614 3.3 0.0011060599999999999 3.3 0.00110616 0 0.00110608 0 0.00110618 3.3 0.0011060999999999998 3.3 0.0011062 0 0.00110612 0 0.00110622 3.3 0.0011061399999999998 3.3 0.0011062399999999999 0 0.00110616 0 0.00110626 3.3 0.00110618 3.3 0.00110628 0 0.0011062 0 0.0011063 3.3 0.00110622 3.3 0.00110632 0 0.0011062399999999999 0 0.00110634 3.3 0.00110626 3.3 0.00110636 0 0.0011062799999999999 0 0.00110638 3.3 0.0011063 3.3 0.0011064 0 0.0011063199999999998 0 0.0011064199999999999 3.3 0.00110634 3.3 0.00110644 0 0.00110636 0 0.00110646 3.3 0.00110638 3.3 0.00110648 0 0.0011064 0 0.0011065 3.3 0.0011064199999999999 3.3 0.00110652 0 0.00110644 0 0.00110654 3.3 0.0011064599999999999 3.3 0.00110656 0 0.00110648 0 0.00110658 3.3 0.0011064999999999998 3.3 0.0011066 0 0.00110652 0 0.00110662 3.3 0.0011065399999999998 3.3 0.0011066399999999999 0 0.00110656 0 0.00110666 3.3 0.00110658 3.3 0.00110668 0 0.0011066 0 0.0011067 3.3 0.00110662 3.3 0.00110672 0 0.0011066399999999999 0 0.00110674 3.3 0.00110666 3.3 0.00110676 0 0.0011066799999999999 0 0.00110678 3.3 0.0011067 3.3 0.0011068 0 0.0011067199999999998 0 0.00110682 3.3 0.00110674 3.3 0.00110684 0 0.0011067599999999998 0 0.0011068599999999999 3.3 0.00110678 3.3 0.00110688 0 0.0011068 0 0.0011069 3.3 0.00110682 3.3 0.00110692 0 0.00110684 0 0.00110694 3.3 0.0011068599999999999 3.3 0.00110696 0 0.00110688 0 0.00110698 3.3 0.0011068999999999999 3.3 0.001107 0 0.00110692 0 0.00110702 3.3 0.0011069399999999998 3.3 0.0011070399999999999 0 0.00110696 0 0.00110706 3.3 0.0011069799999999998 3.3 0.0011070799999999999 0 0.001107 0 0.0011071 3.3 0.00110702 3.3 0.00110712 0 0.0011070399999999999 0 0.00110714 3.3 0.00110706 3.3 0.00110716 0 0.0011070799999999999 0 0.00110718 3.3 0.0011071 3.3 0.0011072 0 0.0011071199999999998 0 0.00110722 3.3 0.00110714 3.3 0.00110724 0 0.0011071599999999998 0 0.0011072599999999999 3.3 0.00110718 3.3 0.00110728 0 0.0011072 0 0.0011073 3.3 0.00110722 3.3 0.00110732 0 0.00110724 0 0.00110734 3.3 0.0011072599999999999 3.3 0.00110736 0 0.00110728 0 0.00110738 3.3 0.0011072999999999999 3.3 0.0011074 0 0.00110732 0 0.00110742 3.3 0.0011073399999999998 3.3 0.00110744 0 0.00110736 0 0.00110746 3.3 0.0011073799999999998 3.3 0.0011074799999999999 0 0.0011074 0 0.0011075 3.3 0.00110742 3.3 0.00110752 0 0.00110744 0 0.00110754 3.3 0.00110746 3.3 0.00110756 0 0.0011074799999999999 0 0.00110758 3.3 0.0011075 3.3 0.0011076 0 0.0011075199999999999 0 0.00110762 3.3 0.00110754 3.3 0.00110764 0 0.0011075599999999998 0 0.00110766 3.3 0.00110758 3.3 0.00110768 0 0.0011075999999999998 0 0.0011076999999999999 3.3 0.00110762 3.3 0.00110772 0 0.00110764 0 0.00110774 3.3 0.00110766 3.3 0.00110776 0 0.00110768 0 0.00110778 3.3 0.0011076999999999999 3.3 0.0011078 0 0.00110772 0 0.00110782 3.3 0.0011077399999999999 3.3 0.00110784 0 0.00110776 0 0.00110786 3.3 0.0011077799999999998 3.3 0.0011078799999999999 0 0.0011078 0 0.0011079 3.3 0.00110782 3.3 0.00110792 0 0.00110784 0 0.00110794 3.3 0.00110786 3.3 0.00110796 0 0.0011078799999999999 0 0.00110798 3.3 0.0011079 3.3 0.001108 0 0.0011079199999999999 0 0.00110802 3.3 0.00110794 3.3 0.00110804 0 0.0011079599999999998 0 0.00110806 3.3 0.00110798 3.3 0.00110808 0 0.0011079999999999998 0 0.0011080999999999999 3.3 0.00110802 3.3 0.00110812 0 0.00110804 0 0.00110814 3.3 0.00110806 3.3 0.00110816 0 0.00110808 0 0.00110818 3.3 0.0011080999999999999 3.3 0.0011082 0 0.00110812 0 0.00110822 3.3 0.0011081399999999999 3.3 0.00110824 0 0.00110816 0 0.00110826 3.3 0.0011081799999999998 3.3 0.00110828 0 0.0011082 0 0.0011083 3.3 0.0011082199999999998 3.3 0.0011083199999999999 0 0.00110824 0 0.00110834 3.3 0.00110826 3.3 0.00110836 0 0.00110828 0 0.00110838 3.3 0.0011083 3.3 0.0011084 0 0.0011083199999999999 0 0.00110842 3.3 0.00110834 3.3 0.00110844 0 0.0011083599999999999 0 0.00110846 3.3 0.00110838 3.3 0.00110848 0 0.0011083999999999998 0 0.0011085 3.3 0.00110842 3.3 0.00110852 0 0.0011084399999999998 0 0.0011085399999999999 3.3 0.00110846 3.3 0.00110856 0 0.00110848 0 0.00110858 3.3 0.0011085 3.3 0.0011086 0 0.00110852 0 0.00110862 3.3 0.0011085399999999999 3.3 0.00110864 0 0.00110856 0 0.00110866 3.3 0.0011085799999999999 3.3 0.00110868 0 0.0011086 0 0.0011087 3.3 0.0011086199999999998 3.3 0.0011087199999999999 0 0.00110864 0 0.00110874 3.3 0.00110866 3.3 0.00110876 0 0.00110868 0 0.00110878 3.3 0.0011087 3.3 0.0011088 0 0.0011087199999999999 0 0.00110882 3.3 0.00110874 3.3 0.00110884 0 0.0011087599999999999 0 0.00110886 3.3 0.00110878 3.3 0.00110888 0 0.0011087999999999998 0 0.0011089 3.3 0.00110882 3.3 0.00110892 0 0.0011088399999999998 0 0.0011089399999999999 3.3 0.00110886 3.3 0.00110896 0 0.00110888 0 0.00110898 3.3 0.0011089 3.3 0.001109 0 0.00110892 0 0.00110902 3.3 0.0011089399999999999 3.3 0.00110904 0 0.00110896 0 0.00110906 3.3 0.0011089799999999999 3.3 0.00110908 0 0.001109 0 0.0011091 3.3 0.0011090199999999998 3.3 0.00110912 0 0.00110904 0 0.00110914 3.3 0.0011090599999999998 3.3 0.0011091599999999999 0 0.00110908 0 0.00110918 3.3 0.0011091 3.3 0.0011092 0 0.00110912 0 0.00110922 3.3 0.00110914 3.3 0.00110924 0 0.0011091599999999999 0 0.00110926 3.3 0.00110918 3.3 0.00110928 0 0.0011091999999999999 0 0.0011093 3.3 0.00110922 3.3 0.00110932 0 0.0011092399999999998 0 0.00110934 3.3 0.00110926 3.3 0.00110936 0 0.0011092799999999998 0 0.0011093799999999999 3.3 0.0011093 3.3 0.0011094 0 0.00110932 0 0.00110942 3.3 0.00110934 3.3 0.00110944 0 0.00110936 0 0.00110946 3.3 0.0011093799999999999 3.3 0.00110948 0 0.0011094 0 0.0011095 3.3 0.0011094199999999999 3.3 0.00110952 0 0.00110944 0 0.00110954 3.3 0.0011094599999999998 3.3 0.0011095599999999999 0 0.00110948 0 0.00110958 3.3 0.0011095 3.3 0.0011096 0 0.00110952 0 0.00110962 3.3 0.00110954 3.3 0.00110964 0 0.0011095599999999999 0 0.00110966 3.3 0.00110958 3.3 0.00110968 0 0.0011095999999999999 0 0.0011097 3.3 0.00110962 3.3 0.00110972 0 0.0011096399999999998 0 0.00110974 3.3 0.00110966 3.3 0.00110976 0 0.0011096799999999998 0 0.0011097799999999999 3.3 0.0011097 3.3 0.0011098 0 0.00110972 0 0.00110982 3.3 0.00110974 3.3 0.00110984 0 0.00110976 0 0.00110986 3.3 0.0011097799999999999 3.3 0.00110988 0 0.0011098 0 0.0011099 3.3 0.0011098199999999999 3.3 0.00110992 0 0.00110984 0 0.00110994 3.3 0.0011098599999999998 3.3 0.00110996 0 0.00110988 0 0.00110998 3.3 0.0011098999999999998 3.3 0.0011099999999999999 0 0.00110992 0 0.00111002 3.3 0.00110994 3.3 0.00111004 0 0.00110996 0 0.00111006 3.3 0.00110998 3.3 0.00111008 0 0.0011099999999999999 0 0.0011101 3.3 0.00111002 3.3 0.00111012 0 0.0011100399999999999 0 0.00111014 3.3 0.00111006 3.3 0.00111016 0 0.0011100799999999998 0 0.0011101799999999999 3.3 0.0011101 3.3 0.0011102 0 0.0011101199999999998 0 0.0011102199999999999 3.3 0.00111014 3.3 0.00111024 0 0.00111016 0 0.00111026 3.3 0.0011101799999999999 3.3 0.00111028 0 0.0011102 0 0.0011103 3.3 0.0011102199999999999 3.3 0.00111032 0 0.00111024 0 0.00111034 3.3 0.0011102599999999998 3.3 0.00111036 0 0.00111028 0 0.00111038 3.3 0.0011102999999999998 3.3 0.0011103999999999999 0 0.00111032 0 0.00111042 3.3 0.00111034 3.3 0.00111044 0 0.00111036 0 0.00111046 3.3 0.00111038 3.3 0.00111048 0 0.0011103999999999999 0 0.0011105 3.3 0.00111042 3.3 0.00111052 0 0.0011104399999999999 0 0.00111054 3.3 0.00111046 3.3 0.00111056 0 0.0011104799999999998 0 0.00111058 3.3 0.0011105 3.3 0.0011106 0 0.0011105199999999998 0 0.0011106199999999999 3.3 0.00111054 3.3 0.00111064 0 0.00111056 0 0.00111066 3.3 0.00111058 3.3 0.00111068 0 0.0011106 0 0.0011107 3.3 0.0011106199999999999 3.3 0.00111072 0 0.00111064 0 0.00111074 3.3 0.0011106599999999999 3.3 0.00111076 0 0.00111068 0 0.00111078 3.3 0.0011106999999999998 3.3 0.0011108 0 0.00111072 0 0.00111082 3.3 0.0011107399999999998 3.3 0.0011108399999999999 0 0.00111076 0 0.00111086 3.3 0.00111078 3.3 0.00111088 0 0.0011108 0 0.0011109 3.3 0.00111082 3.3 0.00111092 0 0.0011108399999999999 0 0.00111094 3.3 0.00111086 3.3 0.00111096 0 0.0011108799999999999 0 0.00111098 3.3 0.0011109 3.3 0.001111 0 0.0011109199999999998 0 0.0011110199999999999 3.3 0.00111094 3.3 0.00111104 0 0.00111096 0 0.00111106 3.3 0.00111098 3.3 0.00111108 0 0.001111 0 0.0011111 3.3 0.0011110199999999999 3.3 0.00111112 0 0.00111104 0 0.00111114 3.3 0.0011110599999999999 3.3 0.00111116 0 0.00111108 0 0.00111118 3.3 0.0011110999999999998 3.3 0.0011112 0 0.00111112 0 0.00111122 3.3 0.0011111399999999998 3.3 0.0011112399999999999 0 0.00111116 0 0.00111126 3.3 0.00111118 3.3 0.00111128 0 0.0011112 0 0.0011113 3.3 0.00111122 3.3 0.00111132 0 0.0011112399999999999 0 0.00111134 3.3 0.00111126 3.3 0.00111136 0 0.0011112799999999999 0 0.00111138 3.3 0.0011113 3.3 0.0011114 0 0.0011113199999999998 0 0.00111142 3.3 0.00111134 3.3 0.00111144 0 0.0011113599999999998 0 0.0011114599999999999 3.3 0.00111138 3.3 0.00111148 0 0.0011114 0 0.0011115 3.3 0.00111142 3.3 0.00111152 0 0.00111144 0 0.00111154 3.3 0.0011114599999999999 3.3 0.00111156 0 0.00111148 0 0.00111158 3.3 0.0011114999999999999 3.3 0.0011116 0 0.00111152 0 0.00111162 3.3 0.0011115399999999998 3.3 0.00111164 0 0.00111156 0 0.00111166 3.3 0.0011115799999999998 3.3 0.0011116799999999999 0 0.0011116 0 0.0011117 3.3 0.00111162 3.3 0.00111172 0 0.00111164 0 0.00111174 3.3 0.00111166 3.3 0.00111176 0 0.0011116799999999999 0 0.00111178 3.3 0.0011117 3.3 0.0011118 0 0.0011117199999999999 0 0.00111182 3.3 0.00111174 3.3 0.00111184 0 0.0011117599999999998 0 0.0011118599999999999 3.3 0.00111178 3.3 0.00111188 0 0.0011118 0 0.0011119 3.3 0.00111182 3.3 0.00111192 0 0.00111184 0 0.00111194 3.3 0.0011118599999999999 3.3 0.00111196 0 0.00111188 0 0.00111198 3.3 0.0011118999999999999 3.3 0.001112 0 0.00111192 0 0.00111202 3.3 0.0011119399999999998 3.3 0.00111204 0 0.00111196 0 0.00111206 3.3 0.0011119799999999998 3.3 0.0011120799999999999 0 0.001112 0 0.0011121 3.3 0.00111202 3.3 0.00111212 0 0.00111204 0 0.00111214 3.3 0.00111206 3.3 0.00111216 0 0.0011120799999999999 0 0.00111218 3.3 0.0011121 3.3 0.0011122 0 0.0011121199999999999 0 0.00111222 3.3 0.00111214 3.3 0.00111224 0 0.0011121599999999998 0 0.00111226 3.3 0.00111218 3.3 0.00111228 0 0.0011121999999999998 0 0.0011122999999999999 3.3 0.00111222 3.3 0.00111232 0 0.00111224 0 0.00111234 3.3 0.00111226 3.3 0.00111236 0 0.00111228 0 0.00111238 3.3 0.0011122999999999999 3.3 0.0011124 0 0.00111232 0 0.00111242 3.3 0.0011123399999999999 3.3 0.00111244 0 0.00111236 0 0.00111246 3.3 0.0011123799999999998 3.3 0.00111248 0 0.0011124 0 0.0011125 3.3 0.0011124199999999998 3.3 0.0011125199999999999 0 0.00111244 0 0.00111254 3.3 0.00111246 3.3 0.00111256 0 0.00111248 0 0.00111258 3.3 0.0011125 3.3 0.0011126 0 0.0011125199999999999 0 0.00111262 3.3 0.00111254 3.3 0.00111264 0 0.0011125599999999999 0 0.00111266 3.3 0.00111258 3.3 0.00111268 0 0.0011125999999999998 0 0.0011126999999999999 3.3 0.00111262 3.3 0.00111272 0 0.00111264 0 0.00111274 3.3 0.00111266 3.3 0.00111276 0 0.00111268 0 0.00111278 3.3 0.0011126999999999999 3.3 0.0011128 0 0.00111272 0 0.00111282 3.3 0.0011127399999999999 3.3 0.00111284 0 0.00111276 0 0.00111286 3.3 0.0011127799999999998 3.3 0.00111288 0 0.0011128 0 0.0011129 3.3 0.0011128199999999998 3.3 0.0011129199999999999 0 0.00111284 0 0.00111294 3.3 0.00111286 3.3 0.00111296 0 0.00111288 0 0.00111298 3.3 0.0011129 3.3 0.001113 0 0.0011129199999999999 0 0.00111302 3.3 0.00111294 3.3 0.00111304 0 0.0011129599999999999 0 0.00111306 3.3 0.00111298 3.3 0.00111308 0 0.0011129999999999998 0 0.0011131 3.3 0.00111302 3.3 0.00111312 0 0.0011130399999999998 0 0.0011131399999999999 3.3 0.00111306 3.3 0.00111316 0 0.00111308 0 0.00111318 3.3 0.0011131 3.3 0.0011132 0 0.00111312 0 0.00111322 3.3 0.0011131399999999999 3.3 0.00111324 0 0.00111316 0 0.00111326 3.3 0.0011131799999999999 3.3 0.00111328 0 0.0011132 0 0.0011133 3.3 0.0011132199999999998 3.3 0.0011133199999999999 0 0.00111324 0 0.00111334 3.3 0.0011132599999999998 3.3 0.0011133599999999999 0 0.00111328 0 0.00111338 3.3 0.0011133 3.3 0.0011134 0 0.0011133199999999999 0 0.00111342 3.3 0.00111334 3.3 0.00111344 0 0.0011133599999999999 0 0.00111346 3.3 0.00111338 3.3 0.00111348 0 0.0011133999999999998 0 0.0011135 3.3 0.00111342 3.3 0.00111352 0 0.0011134399999999998 0 0.0011135399999999999 3.3 0.00111346 3.3 0.00111356 0 0.00111348 0 0.00111358 3.3 0.0011135 3.3 0.0011136 0 0.00111352 0 0.00111362 3.3 0.0011135399999999999 3.3 0.00111364 0 0.00111356 0 0.00111366 3.3 0.0011135799999999999 3.3 0.00111368 0 0.0011136 0 0.0011137 3.3 0.0011136199999999998 3.3 0.00111372 0 0.00111364 0 0.00111374 3.3 0.0011136599999999998 3.3 0.0011137599999999999 0 0.00111368 0 0.00111378 3.3 0.0011137 3.3 0.0011138 0 0.00111372 0 0.00111382 3.3 0.00111374 3.3 0.00111384 0 0.0011137599999999999 0 0.00111386 3.3 0.00111378 3.3 0.00111388 0 0.0011137999999999999 0 0.0011139 3.3 0.00111382 3.3 0.00111392 0 0.0011138399999999998 0 0.00111394 3.3 0.00111386 3.3 0.00111396 0 0.0011138799999999998 0 0.0011139799999999999 3.3 0.0011139 3.3 0.001114 0 0.00111392 0 0.00111402 3.3 0.00111394 3.3 0.00111404 0 0.00111396 0 0.00111406 3.3 0.0011139799999999999 3.3 0.00111408 0 0.001114 0 0.0011141 3.3 0.0011140199999999999 3.3 0.00111412 0 0.00111404 0 0.00111414 3.3 0.0011140599999999998 3.3 0.0011141599999999999 0 0.00111408 0 0.00111418 3.3 0.0011140999999999998 3.3 0.0011141999999999999 0 0.00111412 0 0.00111422 3.3 0.00111414 3.3 0.00111424 0 0.0011141599999999999 0 0.00111426 3.3 0.00111418 3.3 0.00111428 0 0.0011141999999999999 0 0.0011143 3.3 0.00111422 3.3 0.00111432 0 0.0011142399999999998 0 0.00111434 3.3 0.00111426 3.3 0.00111436 0 0.0011142799999999998 0 0.0011143799999999999 3.3 0.0011143 3.3 0.0011144 0 0.00111432 0 0.00111442 3.3 0.00111434 3.3 0.00111444 0 0.00111436 0 0.00111446 3.3 0.0011143799999999999 3.3 0.00111448 0 0.0011144 0 0.0011145 3.3 0.0011144199999999999 3.3 0.00111452 0 0.00111444 0 0.00111454 3.3 0.0011144599999999998 3.3 0.00111456 0 0.00111448 0 0.00111458 3.3 0.0011144999999999998 3.3 0.0011145999999999999 0 0.00111452 0 0.00111462 3.3 0.00111454 3.3 0.00111464 0 0.00111456 0 0.00111466 3.3 0.00111458 3.3 0.00111468 0 0.0011145999999999999 0 0.0011147 3.3 0.00111462 3.3 0.00111472 0 0.0011146399999999999 0 0.00111474 3.3 0.00111466 3.3 0.00111476 0 0.0011146799999999998 0 0.00111478 3.3 0.0011147 3.3 0.0011148 0 0.0011147199999999998 0 0.0011148199999999999 3.3 0.00111474 3.3 0.00111484 0 0.00111476 0 0.00111486 3.3 0.00111478 3.3 0.00111488 0 0.0011148 0 0.0011149 3.3 0.0011148199999999999 3.3 0.00111492 0 0.00111484 0 0.00111494 3.3 0.0011148599999999999 3.3 0.00111496 0 0.00111488 0 0.00111498 3.3 0.0011148999999999998 3.3 0.0011149999999999999 0 0.00111492 0 0.00111502 3.3 0.00111494 3.3 0.00111504 0 0.00111496 0 0.00111506 3.3 0.00111498 3.3 0.00111508 0 0.0011149999999999999 0 0.0011151 3.3 0.00111502 3.3 0.00111512 0 0.0011150399999999999 0 0.00111514 3.3 0.00111506 3.3 0.00111516 0 0.0011150799999999998 0 0.00111518 3.3 0.0011151 3.3 0.0011152 0 0.0011151199999999998 0 0.0011152199999999999 3.3 0.00111514 3.3 0.00111524 0 0.00111516 0 0.00111526 3.3 0.00111518 3.3 0.00111528 0 0.0011152 0 0.0011153 3.3 0.0011152199999999999 3.3 0.00111532 0 0.00111524 0 0.00111534 3.3 0.0011152599999999999 3.3 0.00111536 0 0.00111528 0 0.00111538 3.3 0.0011152999999999998 3.3 0.0011154 0 0.00111532 0 0.00111542 3.3 0.0011153399999999998 3.3 0.0011154399999999999 0 0.00111536 0 0.00111546 3.3 0.00111538 3.3 0.00111548 0 0.0011154 0 0.0011155 3.3 0.00111542 3.3 0.00111552 0 0.0011154399999999999 0 0.00111554 3.3 0.00111546 3.3 0.00111556 0 0.0011154799999999999 0 0.00111558 3.3 0.0011155 3.3 0.0011156 0 0.0011155199999999998 0 0.00111562 3.3 0.00111554 3.3 0.00111564 0 0.0011155599999999998 0 0.0011156599999999999 3.3 0.00111558 3.3 0.00111568 0 0.0011156 0 0.0011157 3.3 0.00111562 3.3 0.00111572 0 0.00111564 0 0.00111574 3.3 0.0011156599999999999 3.3 0.00111576 0 0.00111568 0 0.00111578 3.3 0.0011156999999999999 3.3 0.0011158 0 0.00111572 0 0.00111582 3.3 0.0011157399999999998 3.3 0.0011158399999999999 0 0.00111576 0 0.00111586 3.3 0.00111578 3.3 0.00111588 0 0.0011158 0 0.0011159 3.3 0.00111582 3.3 0.00111592 0 0.0011158399999999999 0 0.00111594 3.3 0.00111586 3.3 0.00111596 0 0.0011158799999999999 0 0.00111598 3.3 0.0011159 3.3 0.001116 0 0.0011159199999999998 0 0.00111602 3.3 0.00111594 3.3 0.00111604 0 0.0011159599999999998 0 0.0011160599999999999 3.3 0.00111598 3.3 0.00111608 0 0.001116 0 0.0011161 3.3 0.00111602 3.3 0.00111612 0 0.00111604 0 0.00111614 3.3 0.0011160599999999999 3.3 0.00111616 0 0.00111608 0 0.00111618 3.3 0.0011160999999999999 3.3 0.0011162 0 0.00111612 0 0.00111622 3.3 0.0011161399999999998 3.3 0.00111624 0 0.00111616 0 0.00111626 3.3 0.0011161799999999998 3.3 0.0011162799999999999 0 0.0011162 0 0.0011163 3.3 0.00111622 3.3 0.00111632 0 0.00111624 0 0.00111634 3.3 0.00111626 3.3 0.00111636 0 0.0011162799999999999 0 0.00111638 3.3 0.0011163 3.3 0.0011164 0 0.0011163199999999999 0 0.00111642 3.3 0.00111634 3.3 0.00111644 0 0.0011163599999999998 0 0.00111646 3.3 0.00111638 3.3 0.00111648 0 0.0011163999999999998 0 0.0011164999999999999 3.3 0.00111642 3.3 0.00111652 0 0.00111644 0 0.00111654 3.3 0.00111646 3.3 0.00111656 0 0.00111648 0 0.00111658 3.3 0.0011164999999999999 3.3 0.0011166 0 0.00111652 0 0.00111662 3.3 0.0011165399999999999 3.3 0.00111664 0 0.00111656 0 0.00111666 3.3 0.0011165799999999998 3.3 0.0011166799999999999 0 0.0011166 0 0.0011167 3.3 0.00111662 3.3 0.00111672 0 0.00111664 0 0.00111674 3.3 0.00111666 3.3 0.00111676 0 0.0011166799999999999 0 0.00111678 3.3 0.0011167 3.3 0.0011168 0 0.0011167199999999999 0 0.00111682 3.3 0.00111674 3.3 0.00111684 0 0.0011167599999999998 0 0.00111686 3.3 0.00111678 3.3 0.00111688 0 0.0011167999999999998 0 0.0011168999999999999 3.3 0.00111682 3.3 0.00111692 0 0.00111684 0 0.00111694 3.3 0.00111686 3.3 0.00111696 0 0.00111688 0 0.00111698 3.3 0.0011168999999999999 3.3 0.001117 0 0.00111692 0 0.00111702 3.3 0.0011169399999999999 3.3 0.00111704 0 0.00111696 0 0.00111706 3.3 0.0011169799999999998 3.3 0.00111708 0 0.001117 0 0.0011171 3.3 0.0011170199999999998 3.3 0.0011171199999999999 0 0.00111704 0 0.00111714 3.3 0.00111706 3.3 0.00111716 0 0.00111708 0 0.00111718 3.3 0.0011171 3.3 0.0011172 0 0.0011171199999999999 0 0.00111722 3.3 0.00111714 3.3 0.00111724 0 0.0011171599999999999 0 0.00111726 3.3 0.00111718 3.3 0.00111728 0 0.0011171999999999998 0 0.0011172999999999999 3.3 0.00111722 3.3 0.00111732 0 0.0011172399999999998 0 0.0011173399999999999 3.3 0.00111726 3.3 0.00111736 0 0.00111728 0 0.00111738 3.3 0.0011172999999999999 3.3 0.0011174 0 0.00111732 0 0.00111742 3.3 0.0011173399999999999 3.3 0.00111744 0 0.00111736 0 0.00111746 3.3 0.0011173799999999998 3.3 0.00111748 0 0.0011174 0 0.0011175 3.3 0.0011174199999999998 3.3 0.0011175199999999999 0 0.00111744 0 0.00111754 3.3 0.00111746 3.3 0.00111756 0 0.00111748 0 0.00111758 3.3 0.0011175 3.3 0.0011176 0 0.0011175199999999999 0 0.00111762 3.3 0.00111754 3.3 0.00111764 0 0.0011175599999999999 0 0.00111766 3.3 0.00111758 3.3 0.00111768 0 0.0011175999999999998 0 0.0011177 3.3 0.00111762 3.3 0.00111772 0 0.0011176399999999998 0 0.0011177399999999999 3.3 0.00111766 3.3 0.00111776 0 0.00111768 0 0.00111778 3.3 0.0011177 3.3 0.0011178 0 0.00111772 0 0.00111782 3.3 0.0011177399999999999 3.3 0.00111784 0 0.00111776 0 0.00111786 3.3 0.0011177799999999999 3.3 0.00111788 0 0.0011178 0 0.0011179 3.3 0.0011178199999999998 3.3 0.00111792 0 0.00111784 0 0.00111794 3.3 0.0011178599999999998 3.3 0.0011179599999999999 0 0.00111788 0 0.00111798 3.3 0.0011179 3.3 0.001118 0 0.00111792 0 0.00111802 3.3 0.00111794 3.3 0.00111804 0 0.0011179599999999999 0 0.00111806 3.3 0.00111798 3.3 0.00111808 0 0.0011179999999999999 0 0.0011181 3.3 0.00111802 3.3 0.00111812 0 0.0011180399999999998 0 0.0011181399999999999 3.3 0.00111806 3.3 0.00111816 0 0.00111808 0 0.00111818 3.3 0.0011181 3.3 0.0011182 0 0.00111812 0 0.00111822 3.3 0.0011181399999999999 3.3 0.00111824 0 0.00111816 0 0.00111826 3.3 0.0011181799999999999 3.3 0.00111828 0 0.0011182 0 0.0011183 3.3 0.0011182199999999998 3.3 0.00111832 0 0.00111824 0 0.00111834 3.3 0.0011182599999999998 3.3 0.0011183599999999999 0 0.00111828 0 0.00111838 3.3 0.0011183 3.3 0.0011184 0 0.00111832 0 0.00111842 3.3 0.00111834 3.3 0.00111844 0 0.0011183599999999999 0 0.00111846 3.3 0.00111838 3.3 0.00111848 0 0.0011183999999999999 0 0.0011185 3.3 0.00111842 3.3 0.00111852 0 0.0011184399999999998 0 0.00111854 3.3 0.00111846 3.3 0.00111856 0 0.0011184799999999998 0 0.0011185799999999999 3.3 0.0011185 3.3 0.0011186 0 0.00111852 0 0.00111862 3.3 0.00111854 3.3 0.00111864 0 0.00111856 0 0.00111866 3.3 0.0011185799999999999 3.3 0.00111868 0 0.0011186 0 0.0011187 3.3 0.0011186199999999999 3.3 0.00111872 0 0.00111864 0 0.00111874 3.3 0.0011186599999999998 3.3 0.00111876 0 0.00111868 0 0.00111878 3.3 0.0011186999999999998 3.3 0.0011187999999999999 0 0.00111872 0 0.00111882 3.3 0.00111874 3.3 0.00111884 0 0.00111876 0 0.00111886 3.3 0.00111878 3.3 0.00111888 0 0.0011187999999999999 0 0.0011189 3.3 0.00111882 3.3 0.00111892 0 0.0011188399999999999 0 0.00111894 3.3 0.00111886 3.3 0.00111896 0 0.0011188799999999998 0 0.0011189799999999999 3.3 0.0011189 3.3 0.001119 0 0.00111892 0 0.00111902 3.3 0.00111894 3.3 0.00111904 0 0.00111896 0 0.00111906 3.3 0.0011189799999999999 3.3 0.00111908 0 0.001119 0 0.0011191 3.3 0.0011190199999999999 3.3 0.00111912 0 0.00111904 0 0.00111914 3.3 0.0011190599999999998 3.3 0.00111916 0 0.00111908 0 0.00111918 3.3 0.0011190999999999998 3.3 0.0011191999999999999 0 0.00111912 0 0.00111922 3.3 0.00111914 3.3 0.00111924 0 0.00111916 0 0.00111926 3.3 0.00111918 3.3 0.00111928 0 0.0011191999999999999 0 0.0011193 3.3 0.00111922 3.3 0.00111932 0 0.0011192399999999999 0 0.00111934 3.3 0.00111926 3.3 0.00111936 0 0.0011192799999999998 0 0.00111938 3.3 0.0011193 3.3 0.0011194 0 0.0011193199999999998 0 0.0011194199999999999 3.3 0.00111934 3.3 0.00111944 0 0.00111936 0 0.00111946 3.3 0.00111938 3.3 0.00111948 0 0.0011194 0 0.0011195 3.3 0.0011194199999999999 3.3 0.00111952 0 0.00111944 0 0.00111954 3.3 0.0011194599999999999 3.3 0.00111956 0 0.00111948 0 0.00111958 3.3 0.0011194999999999998 3.3 0.0011196 0 0.00111952 0 0.00111962 3.3 0.0011195399999999998 3.3 0.0011196399999999999 0 0.00111956 0 0.00111966 3.3 0.00111958 3.3 0.00111968 0 0.0011196 0 0.0011197 3.3 0.00111962 3.3 0.00111972 0 0.0011196399999999999 0 0.00111974 3.3 0.00111966 3.3 0.00111976 0 0.0011196799999999999 0 0.00111978 3.3 0.0011197 3.3 0.0011198 0 0.0011197199999999998 0 0.0011198199999999999 3.3 0.00111974 3.3 0.00111984 0 0.00111976 0 0.00111986 3.3 0.00111978 3.3 0.00111988 0 0.0011198 0 0.0011199 3.3 0.0011198199999999999 3.3 0.00111992 0 0.00111984 0 0.00111994 3.3 0.0011198599999999999 3.3 0.00111996 0 0.00111988 0 0.00111998 3.3 0.0011198999999999998 3.3 0.00112 0 0.00111992 0 0.00112002 3.3 0.0011199399999999998 3.3 0.0011200399999999999 0 0.00111996 0 0.00112006 3.3 0.00111998 3.3 0.00112008 0 0.00112 0 0.0011201 3.3 0.00112002 3.3 0.00112012 0 0.0011200399999999999 0 0.00112014 3.3 0.00112006 3.3 0.00112016 0 0.0011200799999999999 0 0.00112018 3.3 0.0011201 3.3 0.0011202 0 0.0011201199999999998 0 0.00112022 3.3 0.00112014 3.3 0.00112024 0 0.0011201599999999998 0 0.0011202599999999999 3.3 0.00112018 3.3 0.00112028 0 0.0011202 0 0.0011203 3.3 0.00112022 3.3 0.00112032 0 0.00112024 0 0.00112034 3.3 0.0011202599999999999 3.3 0.00112036 0 0.00112028 0 0.00112038 3.3 0.0011202999999999999 3.3 0.0011204 0 0.00112032 0 0.00112042 3.3 0.0011203399999999998 3.3 0.0011204399999999999 0 0.00112036 0 0.00112046 3.3 0.0011203799999999998 3.3 0.0011204799999999999 0 0.0011204 0 0.0011205 3.3 0.00112042 3.3 0.00112052 0 0.0011204399999999999 0 0.00112054 3.3 0.00112046 3.3 0.00112056 0 0.0011204799999999999 0 0.00112058 3.3 0.0011205 3.3 0.0011206 0 0.0011205199999999998 0 0.00112062 3.3 0.00112054 3.3 0.00112064 0 0.0011205599999999998 0 0.0011206599999999999 3.3 0.00112058 3.3 0.00112068 0 0.0011206 0 0.0011207 3.3 0.00112062 3.3 0.00112072 0 0.00112064 0 0.00112074 3.3 0.0011206599999999999 3.3 0.00112076 0 0.00112068 0 0.00112078 3.3 0.0011206999999999999 3.3 0.0011208 0 0.00112072 0 0.00112082 3.3 0.0011207399999999998 3.3 0.00112084 0 0.00112076 0 0.00112086 3.3 0.0011207799999999998 3.3 0.0011208799999999999 0 0.0011208 0 0.0011209 3.3 0.00112082 3.3 0.00112092 0 0.00112084 0 0.00112094 3.3 0.00112086 3.3 0.00112096 0 0.0011208799999999999 0 0.00112098 3.3 0.0011209 3.3 0.001121 0 0.0011209199999999999 0 0.00112102 3.3 0.00112094 3.3 0.00112104 0 0.0011209599999999998 0 0.00112106 3.3 0.00112098 3.3 0.00112108 0 0.0011209999999999998 0 0.0011210999999999999 3.3 0.00112102 3.3 0.00112112 0 0.00112104 0 0.00112114 3.3 0.00112106 3.3 0.00112116 0 0.00112108 0 0.00112118 3.3 0.0011210999999999999 3.3 0.0011212 0 0.00112112 0 0.00112122 3.3 0.0011211399999999999 3.3 0.00112124 0 0.00112116 0 0.00112126 3.3 0.0011211799999999998 3.3 0.0011212799999999999 0 0.0011212 0 0.0011213 3.3 0.00112122 3.3 0.00112132 0 0.00112124 0 0.00112134 3.3 0.00112126 3.3 0.00112136 0 0.0011212799999999999 0 0.00112138 3.3 0.0011213 3.3 0.0011214 0 0.0011213199999999999 0 0.00112142 3.3 0.00112134 3.3 0.00112144 0 0.0011213599999999998 0 0.00112146 3.3 0.00112138 3.3 0.00112148 0 0.0011213999999999998 0 0.0011214999999999999 3.3 0.00112142 3.3 0.00112152 0 0.00112144 0 0.00112154 3.3 0.00112146 3.3 0.00112156 0 0.00112148 0 0.00112158 3.3 0.0011214999999999999 3.3 0.0011216 0 0.00112152 0 0.00112162 3.3 0.0011215399999999999 3.3 0.00112164 0 0.00112156 0 0.00112166 3.3 0.0011215799999999998 3.3 0.00112168 0 0.0011216 0 0.0011217 3.3 0.0011216199999999998 3.3 0.0011217199999999999 0 0.00112164 0 0.00112174 3.3 0.00112166 3.3 0.00112176 0 0.00112168 0 0.00112178 3.3 0.0011217 3.3 0.0011218 0 0.0011217199999999999 0 0.00112182 3.3 0.00112174 3.3 0.00112184 0 0.0011217599999999999 0 0.00112186 3.3 0.00112178 3.3 0.00112188 0 0.0011217999999999998 0 0.0011219 3.3 0.00112182 3.3 0.00112192 0 0.0011218399999999998 0 0.0011219399999999999 3.3 0.00112186 3.3 0.00112196 0 0.00112188 0 0.00112198 3.3 0.0011219 3.3 0.001122 0 0.00112192 0 0.00112202 3.3 0.0011219399999999999 3.3 0.00112204 0 0.00112196 0 0.00112206 3.3 0.0011219799999999999 3.3 0.00112208 0 0.001122 0 0.0011221 3.3 0.0011220199999999998 3.3 0.0011221199999999999 0 0.00112204 0 0.00112214 3.3 0.00112206 3.3 0.00112216 0 0.00112208 0 0.00112218 3.3 0.0011221 3.3 0.0011222 0 0.0011221199999999999 0 0.00112222 3.3 0.00112214 3.3 0.00112224 0 0.0011221599999999999 0 0.00112226 3.3 0.00112218 3.3 0.00112228 0 0.0011221999999999998 0 0.0011223 3.3 0.00112222 3.3 0.00112232 0 0.0011222399999999998 0 0.0011223399999999999 3.3 0.00112226 3.3 0.00112236 0 0.00112228 0 0.00112238 3.3 0.0011223 3.3 0.0011224 0 0.00112232 0 0.00112242 3.3 0.0011223399999999999 3.3 0.00112244 0 0.00112236 0 0.00112246 3.3 0.0011223799999999999 3.3 0.00112248 0 0.0011224 0 0.0011225 3.3 0.0011224199999999998 3.3 0.00112252 0 0.00112244 0 0.00112254 3.3 0.0011224599999999998 3.3 0.0011225599999999999 0 0.00112248 0 0.00112258 3.3 0.0011225 3.3 0.0011226 0 0.00112252 0 0.00112262 3.3 0.00112254 3.3 0.00112264 0 0.0011225599999999999 0 0.00112266 3.3 0.00112258 3.3 0.00112268 0 0.0011225999999999999 0 0.0011227 3.3 0.00112262 3.3 0.00112272 0 0.0011226399999999998 0 0.00112274 3.3 0.00112266 3.3 0.00112276 0 0.0011226799999999998 0 0.0011227799999999999 3.3 0.0011227 3.3 0.0011228 0 0.00112272 0 0.00112282 3.3 0.00112274 3.3 0.00112284 0 0.00112276 0 0.00112286 3.3 0.0011227799999999999 3.3 0.00112288 0 0.0011228 0 0.0011229 3.3 0.0011228199999999999 3.3 0.00112292 0 0.00112284 0 0.00112294 3.3 0.0011228599999999998 3.3 0.0011229599999999999 0 0.00112288 0 0.00112298 3.3 0.0011229 3.3 0.001123 0 0.00112292 0 0.00112302 3.3 0.00112294 3.3 0.00112304 0 0.0011229599999999999 0 0.00112306 3.3 0.00112298 3.3 0.00112308 0 0.0011229999999999999 0 0.0011231 3.3 0.00112302 3.3 0.00112312 0 0.0011230399999999998 0 0.00112314 3.3 0.00112306 3.3 0.00112316 0 0.0011230799999999998 0 0.0011231799999999999 3.3 0.0011231 3.3 0.0011232 0 0.00112312 0 0.00112322 3.3 0.00112314 3.3 0.00112324 0 0.00112316 0 0.00112326 3.3 0.0011231799999999999 3.3 0.00112328 0 0.0011232 0 0.0011233 3.3 0.0011232199999999999 3.3 0.00112332 0 0.00112324 0 0.00112334 3.3 0.0011232599999999998 3.3 0.00112336 0 0.00112328 0 0.00112338 3.3 0.0011232999999999998 3.3 0.0011233999999999999 0 0.00112332 0 0.00112342 3.3 0.00112334 3.3 0.00112344 0 0.00112336 0 0.00112346 3.3 0.00112338 3.3 0.00112348 0 0.0011233999999999999 0 0.0011235 3.3 0.00112342 3.3 0.00112352 0 0.0011234399999999999 0 0.00112354 3.3 0.00112346 3.3 0.00112356 0 0.0011234799999999998 0 0.0011235799999999999 3.3 0.0011235 3.3 0.0011236 0 0.0011235199999999998 0 0.0011236199999999999 3.3 0.00112354 3.3 0.00112364 0 0.00112356 0 0.00112366 3.3 0.0011235799999999999 3.3 0.00112368 0 0.0011236 0 0.0011237 3.3 0.0011236199999999999 3.3 0.00112372 0 0.00112364 0 0.00112374 3.3 0.0011236599999999998 3.3 0.00112376 0 0.00112368 0 0.00112378 3.3 0.0011236999999999998 3.3 0.0011237999999999999 0 0.00112372 0 0.00112382 3.3 0.00112374 3.3 0.00112384 0 0.00112376 0 0.00112386 3.3 0.00112378 3.3 0.00112388 0 0.0011237999999999999 0 0.0011239 3.3 0.00112382 3.3 0.00112392 0 0.0011238399999999999 0 0.00112394 3.3 0.00112386 3.3 0.00112396 0 0.0011238799999999998 0 0.00112398 3.3 0.0011239 3.3 0.001124 0 0.0011239199999999998 0 0.0011240199999999999 3.3 0.00112394 3.3 0.00112404 0 0.00112396 0 0.00112406 3.3 0.00112398 3.3 0.00112408 0 0.001124 0 0.0011241 3.3 0.0011240199999999999 3.3 0.00112412 0 0.00112404 0 0.00112414 3.3 0.0011240599999999999 3.3 0.00112416 0 0.00112408 0 0.00112418 3.3 0.0011240999999999998 3.3 0.0011242 0 0.00112412 0 0.00112422 3.3 0.0011241399999999998 3.3 0.0011242399999999999 0 0.00112416 0 0.00112426 3.3 0.00112418 3.3 0.00112428 0 0.0011242 0 0.0011243 3.3 0.00112422 3.3 0.00112432 0 0.0011242399999999999 0 0.00112434 3.3 0.00112426 3.3 0.00112436 0 0.0011242799999999999 0 0.00112438 3.3 0.0011243 3.3 0.0011244 0 0.0011243199999999998 0 0.0011244199999999999 3.3 0.00112434 3.3 0.00112444 0 0.0011243599999999998 0 0.0011244599999999999 3.3 0.00112438 3.3 0.00112448 0 0.0011244 0 0.0011245 3.3 0.0011244199999999999 3.3 0.00112452 0 0.00112444 0 0.00112454 3.3 0.0011244599999999999 3.3 0.00112456 0 0.00112448 0 0.00112458 3.3 0.0011244999999999998 3.3 0.0011246 0 0.00112452 0 0.00112462 3.3 0.0011245399999999998 3.3 0.0011246399999999999 0 0.00112456 0 0.00112466 3.3 0.00112458 3.3 0.00112468 0 0.0011246 0 0.0011247 3.3 0.00112462 3.3 0.00112472 0 0.0011246399999999999 0 0.00112474 3.3 0.00112466 3.3 0.00112476 0 0.0011246799999999999 0 0.00112478 3.3 0.0011247 3.3 0.0011248 0 0.0011247199999999998 0 0.00112482 3.3 0.00112474 3.3 0.00112484 0 0.0011247599999999998 0 0.0011248599999999999 3.3 0.00112478 3.3 0.00112488 0 0.0011248 0 0.0011249 3.3 0.00112482 3.3 0.00112492 0 0.00112484 0 0.00112494 3.3 0.0011248599999999999 3.3 0.00112496 0 0.00112488 0 0.00112498 3.3 0.0011248999999999999 3.3 0.001125 0 0.00112492 0 0.00112502 3.3 0.0011249399999999998 3.3 0.00112504 0 0.00112496 0 0.00112506 3.3 0.0011249799999999998 3.3 0.0011250799999999999 0 0.001125 0 0.0011251 3.3 0.00112502 3.3 0.00112512 0 0.00112504 0 0.00112514 3.3 0.00112506 3.3 0.00112516 0 0.0011250799999999999 0 0.00112518 3.3 0.0011251 3.3 0.0011252 0 0.0011251199999999999 0 0.00112522 3.3 0.00112514 3.3 0.00112524 0 0.0011251599999999998 0 0.0011252599999999999 3.3 0.00112518 3.3 0.00112528 0 0.0011252 0 0.0011253 3.3 0.00112522 3.3 0.00112532 0 0.00112524 0 0.00112534 3.3 0.0011252599999999999 3.3 0.00112536 0 0.00112528 0 0.00112538 3.3 0.0011252999999999999 3.3 0.0011254 0 0.00112532 0 0.00112542 3.3 0.0011253399999999998 3.3 0.00112544 0 0.00112536 0 0.00112546 3.3 0.0011253799999999998 3.3 0.0011254799999999999 0 0.0011254 0 0.0011255 3.3 0.00112542 3.3 0.00112552 0 0.00112544 0 0.00112554 3.3 0.00112546 3.3 0.00112556 0 0.0011254799999999999 0 0.00112558 3.3 0.0011255 3.3 0.0011256 0 0.0011255199999999999 0 0.00112562 3.3 0.00112554 3.3 0.00112564 0 0.0011255599999999998 0 0.00112566 3.3 0.00112558 3.3 0.00112568 0 0.0011255999999999998 0 0.0011256999999999999 3.3 0.00112562 3.3 0.00112572 0 0.00112564 0 0.00112574 3.3 0.00112566 3.3 0.00112576 0 0.00112568 0 0.00112578 3.3 0.0011256999999999999 3.3 0.0011258 0 0.00112572 0 0.00112582 3.3 0.0011257399999999999 3.3 0.00112584 0 0.00112576 0 0.00112586 3.3 0.0011257799999999998 3.3 0.00112588 0 0.0011258 0 0.0011259 3.3 0.0011258199999999998 3.3 0.0011259199999999999 0 0.00112584 0 0.00112594 3.3 0.00112586 3.3 0.00112596 0 0.00112588 0 0.00112598 3.3 0.0011259 3.3 0.001126 0 0.0011259199999999999 0 0.00112602 3.3 0.00112594 3.3 0.00112604 0 0.0011259599999999999 0 0.00112606 3.3 0.00112598 3.3 0.00112608 0 0.0011259999999999998 0 0.0011260999999999999 3.3 0.00112602 3.3 0.00112612 0 0.00112604 0 0.00112614 3.3 0.00112606 3.3 0.00112616 0 0.00112608 0 0.00112618 3.3 0.0011260999999999999 3.3 0.0011262 0 0.00112612 0 0.00112622 3.3 0.0011261399999999999 3.3 0.00112624 0 0.00112616 0 0.00112626 3.3 0.0011261799999999998 3.3 0.00112628 0 0.0011262 0 0.0011263 3.3 0.0011262199999999998 3.3 0.0011263199999999999 0 0.00112624 0 0.00112634 3.3 0.00112626 3.3 0.00112636 0 0.00112628 0 0.00112638 3.3 0.0011263 3.3 0.0011264 0 0.0011263199999999999 0 0.00112642 3.3 0.00112634 3.3 0.00112644 0 0.0011263599999999999 0 0.00112646 3.3 0.00112638 3.3 0.00112648 0 0.0011263999999999998 0 0.0011265 3.3 0.00112642 3.3 0.00112652 0 0.0011264399999999998 0 0.0011265399999999999 3.3 0.00112646 3.3 0.00112656 0 0.00112648 0 0.00112658 3.3 0.0011265 3.3 0.0011266 0 0.00112652 0 0.00112662 3.3 0.0011265399999999999 3.3 0.00112664 0 0.00112656 0 0.00112666 3.3 0.0011265799999999999 3.3 0.00112668 0 0.0011266 0 0.0011267 3.3 0.0011266199999999998 3.3 0.00112672 0 0.00112664 0 0.00112674 3.3 0.0011266599999999998 3.3 0.0011267599999999999 0 0.00112668 0 0.00112678 3.3 0.0011267 3.3 0.0011268 0 0.00112672 0 0.00112682 3.3 0.00112674 3.3 0.00112684 0 0.0011267599999999999 0 0.00112686 3.3 0.00112678 3.3 0.00112688 0 0.0011267999999999999 0 0.0011269 3.3 0.00112682 3.3 0.00112692 0 0.0011268399999999998 0 0.0011269399999999999 3.3 0.00112686 3.3 0.00112696 0 0.00112688 0 0.00112698 3.3 0.0011269 3.3 0.001127 0 0.00112692 0 0.00112702 3.3 0.0011269399999999999 3.3 0.00112704 0 0.00112696 0 0.00112706 3.3 0.0011269799999999999 3.3 0.00112708 0 0.001127 0 0.0011271 3.3 0.0011270199999999998 3.3 0.00112712 0 0.00112704 0 0.00112714 3.3 0.0011270599999999998 3.3 0.0011271599999999999 0 0.00112708 0 0.00112718 3.3 0.0011271 3.3 0.0011272 0 0.00112712 0 0.00112722 3.3 0.00112714 3.3 0.00112724 0 0.0011271599999999999 0 0.00112726 3.3 0.00112718 3.3 0.00112728 0 0.0011271999999999999 0 0.0011273 3.3 0.00112722 3.3 0.00112732 0 0.0011272399999999998 0 0.00112734 3.3 0.00112726 3.3 0.00112736 0 0.0011272799999999998 0 0.0011273799999999999 3.3 0.0011273 3.3 0.0011274 0 0.00112732 0 0.00112742 3.3 0.00112734 3.3 0.00112744 0 0.00112736 0 0.00112746 3.3 0.0011273799999999999 3.3 0.00112748 0 0.0011274 0 0.0011275 3.3 0.0011274199999999999 3.3 0.00112752 0 0.00112744 0 0.00112754 3.3 0.0011274599999999998 3.3 0.0011275599999999999 0 0.00112748 0 0.00112758 3.3 0.0011274999999999998 3.3 0.0011275999999999999 0 0.00112752 0 0.00112762 3.3 0.00112754 3.3 0.00112764 0 0.0011275599999999999 0 0.00112766 3.3 0.00112758 3.3 0.00112768 0 0.0011275999999999999 0 0.0011277 3.3 0.00112762 3.3 0.00112772 0 0.0011276399999999998 0 0.00112774 3.3 0.00112766 3.3 0.00112776 0 0.0011276799999999998 0 0.0011277799999999999 3.3 0.0011277 3.3 0.0011278 0 0.00112772 0 0.00112782 3.3 0.00112774 3.3 0.00112784 0 0.00112776 0 0.00112786 3.3 0.0011277799999999999 3.3 0.00112788 0 0.0011278 0 0.0011279 3.3 0.0011278199999999999 3.3 0.00112792 0 0.00112784 0 0.00112794 3.3 0.0011278599999999998 3.3 0.00112796 0 0.00112788 0 0.00112798 3.3 0.0011278999999999998 3.3 0.0011279999999999999 0 0.00112792 0 0.00112802 3.3 0.00112794 3.3 0.00112804 0 0.00112796 0 0.00112806 3.3 0.00112798 3.3 0.00112808 0 0.0011279999999999999 0 0.0011281 3.3 0.00112802 3.3 0.00112812 0 0.0011280399999999999 0 0.00112814 3.3 0.00112806 3.3 0.00112816 0 0.0011280799999999998 0 0.00112818 3.3 0.0011281 3.3 0.0011282 0 0.0011281199999999998 0 0.0011282199999999999 3.3 0.00112814 3.3 0.00112824 0 0.00112816 0 0.00112826 3.3 0.00112818 3.3 0.00112828 0 0.0011282 0 0.0011283 3.3 0.0011282199999999999 3.3 0.00112832 0 0.00112824 0 0.00112834 3.3 0.0011282599999999999 3.3 0.00112836 0 0.00112828 0 0.00112838 3.3 0.0011282999999999998 3.3 0.0011283999999999999 0 0.00112832 0 0.00112842 3.3 0.00112834 3.3 0.00112844 0 0.00112836 0 0.00112846 3.3 0.00112838 3.3 0.00112848 0 0.0011283999999999999 0 0.0011285 3.3 0.00112842 3.3 0.00112852 0 0.0011284399999999999 0 0.00112854 3.3 0.00112846 3.3 0.00112856 0 0.0011284799999999998 0 0.00112858 3.3 0.0011285 3.3 0.0011286 0 0.0011285199999999998 0 0.0011286199999999999 3.3 0.00112854 3.3 0.00112864 0 0.00112856 0 0.00112866 3.3 0.00112858 3.3 0.00112868 0 0.0011286 0 0.0011287 3.3 0.0011286199999999999 3.3 0.00112872 0 0.00112864 0 0.00112874 3.3 0.0011286599999999999 3.3 0.00112876 0 0.00112868 0 0.00112878 3.3 0.0011286999999999998 3.3 0.0011288 0 0.00112872 0 0.00112882 3.3 0.0011287399999999998 3.3 0.0011288399999999999 0 0.00112876 0 0.00112886 3.3 0.00112878 3.3 0.00112888 0 0.0011288 0 0.0011289 3.3 0.00112882 3.3 0.00112892 0 0.0011288399999999999 0 0.00112894 3.3 0.00112886 3.3 0.00112896 0 0.0011288799999999999 0 0.00112898 3.3 0.0011289 3.3 0.001129 0 0.0011289199999999998 0 0.00112902 3.3 0.00112894 3.3 0.00112904 0 0.0011289599999999998 0 0.0011290599999999999 3.3 0.00112898 3.3 0.00112908 0 0.001129 0 0.0011291 3.3 0.00112902 3.3 0.00112912 0 0.00112904 0 0.00112914 3.3 0.0011290599999999999 3.3 0.00112916 0 0.00112908 0 0.00112918 3.3 0.0011290999999999999 3.3 0.0011292 0 0.00112912 0 0.00112922 3.3 0.0011291399999999998 3.3 0.0011292399999999999 0 0.00112916 0 0.00112926 3.3 0.00112918 3.3 0.00112928 0 0.0011292 0 0.0011293 3.3 0.00112922 3.3 0.00112932 0 0.0011292399999999999 0 0.00112934 3.3 0.00112926 3.3 0.00112936 0 0.0011292799999999999 0 0.00112938 3.3 0.0011293 3.3 0.0011294 0 0.0011293199999999998 0 0.00112942 3.3 0.00112934 3.3 0.00112944 0 0.0011293599999999998 0 0.0011294599999999999 3.3 0.00112938 3.3 0.00112948 0 0.0011294 0 0.0011295 3.3 0.00112942 3.3 0.00112952 0 0.00112944 0 0.00112954 3.3 0.0011294599999999999 3.3 0.00112956 0 0.00112948 0 0.00112958 3.3 0.0011294999999999999 3.3 0.0011296 0 0.00112952 0 0.00112962 3.3 0.0011295399999999998 3.3 0.00112964 0 0.00112956 0 0.00112966 3.3 0.0011295799999999998 3.3 0.0011296799999999999 0 0.0011296 0 0.0011297 3.3 0.00112962 3.3 0.00112972 0 0.00112964 0 0.00112974 3.3 0.00112966 3.3 0.00112976 0 0.0011296799999999999 0 0.00112978 3.3 0.0011297 3.3 0.0011298 0 0.0011297199999999999 0 0.00112982 3.3 0.00112974 3.3 0.00112984 0 0.0011297599999999998 0 0.00112986 3.3 0.00112978 3.3 0.00112988 0 0.0011297999999999998 0 0.0011298999999999999 3.3 0.00112982 3.3 0.00112992 0 0.00112984 0 0.00112994 3.3 0.00112986 3.3 0.00112996 0 0.00112988 0 0.00112998 3.3 0.0011298999999999999 3.3 0.00113 0 0.00112992 0 0.00113002 3.3 0.0011299399999999999 3.3 0.00113004 0 0.00112996 0 0.00113006 3.3 0.0011299799999999998 3.3 0.0011300799999999999 0 0.00113 0 0.0011301 3.3 0.00113002 3.3 0.00113012 0 0.00113004 0 0.00113014 3.3 0.00113006 3.3 0.00113016 0 0.0011300799999999999 0 0.00113018 3.3 0.0011301 3.3 0.0011302 0 0.0011301199999999999 0 0.00113022 3.3 0.00113014 3.3 0.00113024 0 0.0011301599999999998 0 0.00113026 3.3 0.00113018 3.3 0.00113028 0 0.0011301999999999998 0 0.0011302999999999999 3.3 0.00113022 3.3 0.00113032 0 0.00113024 0 0.00113034 3.3 0.00113026 3.3 0.00113036 0 0.00113028 0 0.00113038 3.3 0.0011302999999999999 3.3 0.0011304 0 0.00113032 0 0.00113042 3.3 0.0011303399999999999 3.3 0.00113044 0 0.00113036 0 0.00113046 3.3 0.0011303799999999998 3.3 0.00113048 0 0.0011304 0 0.0011305 3.3 0.0011304199999999998 3.3 0.0011305199999999999 0 0.00113044 0 0.00113054 3.3 0.00113046 3.3 0.00113056 0 0.00113048 0 0.00113058 3.3 0.0011305 3.3 0.0011306 0 0.0011305199999999999 0 0.00113062 3.3 0.00113054 3.3 0.00113064 0 0.0011305599999999999 0 0.00113066 3.3 0.00113058 3.3 0.00113068 0 0.0011305999999999998 0 0.0011306999999999999 3.3 0.00113062 3.3 0.00113072 0 0.0011306399999999998 0 0.0011307399999999999 3.3 0.00113066 3.3 0.00113076 0 0.00113068 0 0.00113078 3.3 0.0011306999999999999 3.3 0.0011308 0 0.00113072 0 0.00113082 3.3 0.0011307399999999999 3.3 0.00113084 0 0.00113076 0 0.00113086 3.3 0.0011307799999999998 3.3 0.00113088 0 0.0011308 0 0.0011309 3.3 0.0011308199999999998 3.3 0.0011309199999999999 0 0.00113084 0 0.00113094 3.3 0.00113086 3.3 0.00113096 0 0.00113088 0 0.00113098 3.3 0.0011309 3.3 0.001131 0 0.0011309199999999999 0 0.00113102 3.3 0.00113094 3.3 0.00113104 0 0.0011309599999999999 0 0.00113106 3.3 0.00113098 3.3 0.00113108 0 0.0011309999999999998 0 0.0011311 3.3 0.00113102 3.3 0.00113112 0 0.0011310399999999998 0 0.0011311399999999999 3.3 0.00113106 3.3 0.00113116 0 0.00113108 0 0.00113118 3.3 0.0011311 3.3 0.0011312 0 0.00113112 0 0.00113122 3.3 0.0011311399999999999 3.3 0.00113124 0 0.00113116 0 0.00113126 3.3 0.0011311799999999999 3.3 0.00113128 0 0.0011312 0 0.0011313 3.3 0.0011312199999999998 3.3 0.00113132 0 0.00113124 0 0.00113134 3.3 0.0011312599999999998 3.3 0.0011313599999999999 0 0.00113128 0 0.00113138 3.3 0.0011313 3.3 0.0011314 0 0.00113132 0 0.00113142 3.3 0.00113134 3.3 0.00113144 0 0.0011313599999999999 0 0.00113146 3.3 0.00113138 3.3 0.00113148 0 0.0011313999999999999 0 0.0011315 3.3 0.00113142 3.3 0.00113152 0 0.0011314399999999998 0 0.0011315399999999999 3.3 0.00113146 3.3 0.00113156 0 0.0011314799999999998 0 0.0011315799999999999 3.3 0.0011315 3.3 0.0011316 0 0.00113152 0 0.00113162 3.3 0.0011315399999999999 3.3 0.00113164 0 0.00113156 0 0.00113166 3.3 0.0011315799999999999 3.3 0.00113168 0 0.0011316 0 0.0011317 3.3 0.0011316199999999998 3.3 0.00113172 0 0.00113164 0 0.00113174 3.3 0.0011316599999999998 3.3 0.0011317599999999999 0 0.00113168 0 0.00113178 3.3 0.0011317 3.3 0.0011318 0 0.00113172 0 0.00113182 3.3 0.00113174 3.3 0.00113184 0 0.0011317599999999999 0 0.00113186 3.3 0.00113178 3.3 0.00113188 0 0.0011317999999999999 0 0.0011319 3.3 0.00113182 3.3 0.00113192 0 0.0011318399999999998 0 0.00113194 3.3 0.00113186 3.3 0.00113196 0 0.0011318799999999998 0 0.0011319799999999999 3.3 0.0011319 3.3 0.001132 0 0.00113192 0 0.00113202 3.3 0.00113194 3.3 0.00113204 0 0.00113196 0 0.00113206 3.3 0.0011319799999999999 3.3 0.00113208 0 0.001132 0 0.0011321 3.3 0.0011320199999999999 3.3 0.00113212 0 0.00113204 0 0.00113214 3.3 0.0011320599999999998 3.3 0.00113216 0 0.00113208 0 0.00113218 3.3 0.0011320999999999998 3.3 0.0011321999999999999 0 0.00113212 0 0.00113222 3.3 0.00113214 3.3 0.00113224 0 0.00113216 0 0.00113226 3.3 0.00113218 3.3 0.00113228 0 0.0011321999999999999 0 0.0011323 3.3 0.00113222 3.3 0.00113232 0 0.0011322399999999999 0 0.00113234 3.3 0.00113226 3.3 0.00113236 0 0.0011322799999999998 0 0.0011323799999999999 3.3 0.0011323 3.3 0.0011324 0 0.00113232 0 0.00113242 3.3 0.00113234 3.3 0.00113244 0 0.00113236 0 0.00113246 3.3 0.0011323799999999999 3.3 0.00113248 0 0.0011324 0 0.0011325 3.3 0.0011324199999999999 3.3 0.00113252 0 0.00113244 0 0.00113254 3.3 0.0011324599999999998 3.3 0.00113256 0 0.00113248 0 0.00113258 3.3 0.0011324999999999998 3.3 0.0011325999999999999 0 0.00113252 0 0.00113262 3.3 0.00113254 3.3 0.00113264 0 0.00113256 0 0.00113266 3.3 0.00113258 3.3 0.00113268 0 0.0011325999999999999 0 0.0011327 3.3 0.00113262 3.3 0.00113272 0 0.0011326399999999999 0 0.00113274 3.3 0.00113266 3.3 0.00113276 0 0.0011326799999999998 0 0.00113278 3.3 0.0011327 3.3 0.0011328 0 0.0011327199999999998 0 0.0011328199999999999 3.3 0.00113274 3.3 0.00113284 0 0.00113276 0 0.00113286 3.3 0.00113278 3.3 0.00113288 0 0.0011328 0 0.0011329 3.3 0.0011328199999999999 3.3 0.00113292 0 0.00113284 0 0.00113294 3.3 0.0011328599999999999 3.3 0.00113296 0 0.00113288 0 0.00113298 3.3 0.0011328999999999998 3.3 0.001133 0 0.00113292 0 0.00113302 3.3 0.0011329399999999998 3.3 0.0011330399999999999 0 0.00113296 0 0.00113306 3.3 0.00113298 3.3 0.00113308 0 0.001133 0 0.0011331 3.3 0.00113302 3.3 0.00113312 0 0.0011330399999999999 0 0.00113314 3.3 0.00113306 3.3 0.00113316 0 0.0011330799999999999 0 0.00113318 3.3 0.0011331 3.3 0.0011332 0 0.0011331199999999998 0 0.0011332199999999999 3.3 0.00113314 3.3 0.00113324 0 0.00113316 0 0.00113326 3.3 0.00113318 3.3 0.00113328 0 0.0011332 0 0.0011333 3.3 0.0011332199999999999 3.3 0.00113332 0 0.00113324 0 0.00113334 3.3 0.0011332599999999999 3.3 0.00113336 0 0.00113328 0 0.00113338 3.3 0.0011332999999999998 3.3 0.0011334 0 0.00113332 0 0.00113342 3.3 0.0011333399999999998 3.3 0.0011334399999999999 0 0.00113336 0 0.00113346 3.3 0.00113338 3.3 0.00113348 0 0.0011334 0 0.0011335 3.3 0.00113342 3.3 0.00113352 0 0.0011334399999999999 0 0.00113354 3.3 0.00113346 3.3 0.00113356 0 0.0011334799999999999 0 0.00113358 3.3 0.0011335 3.3 0.0011336 0 0.0011335199999999998 0 0.00113362 3.3 0.00113354 3.3 0.00113364 0 0.0011335599999999998 0 0.0011336599999999999 3.3 0.00113358 3.3 0.00113368 0 0.0011336 0 0.0011337 3.3 0.00113362 3.3 0.00113372 0 0.00113364 0 0.00113374 3.3 0.0011336599999999999 3.3 0.00113376 0 0.00113368 0 0.00113378 3.3 0.0011336999999999999 3.3 0.0011338 0 0.00113372 0 0.00113382 3.3 0.0011337399999999998 3.3 0.0011338399999999999 0 0.00113376 0 0.00113386 3.3 0.0011337799999999998 3.3 0.0011338799999999999 0 0.0011338 0 0.0011339 3.3 0.00113382 3.3 0.00113392 0 0.0011338399999999999 0 0.00113394 3.3 0.00113386 3.3 0.00113396 0 0.0011338799999999999 0 0.00113398 3.3 0.0011339 3.3 0.001134 0 0.0011339199999999998 0 0.00113402 3.3 0.00113394 3.3 0.00113404 0 0.0011339599999999998 0 0.0011340599999999999 3.3 0.00113398 3.3 0.00113408 0 0.001134 0 0.0011341 3.3 0.00113402 3.3 0.00113412 0 0.00113404 0 0.00113414 3.3 0.0011340599999999999 3.3 0.00113416 0 0.00113408 0 0.00113418 3.3 0.0011340999999999999 3.3 0.0011342 0 0.00113412 0 0.00113422 3.3 0.0011341399999999998 3.3 0.00113424 0 0.00113416 0 0.00113426 3.3 0.0011341799999999998 3.3 0.0011342799999999999 0 0.0011342 0 0.0011343 3.3 0.00113422 3.3 0.00113432 0 0.00113424 0 0.00113434 3.3 0.00113426 3.3 0.00113436 0 0.0011342799999999999 0 0.00113438 3.3 0.0011343 3.3 0.0011344 0 0.0011343199999999999 0 0.00113442 3.3 0.00113434 3.3 0.00113444 0 0.0011343599999999998 0 0.00113446 3.3 0.00113438 3.3 0.00113448 0 0.0011343999999999998 0 0.0011344999999999999 3.3 0.00113442 3.3 0.00113452 0 0.00113444 0 0.00113454 3.3 0.00113446 3.3 0.00113456 0 0.00113448 0 0.00113458 3.3 0.0011344999999999999 3.3 0.0011346 0 0.00113452 0 0.00113462 3.3 0.0011345399999999999 3.3 0.00113464 0 0.00113456 0 0.00113466 3.3 0.0011345799999999998 3.3 0.0011346799999999999 0 0.0011346 0 0.0011347 3.3 0.0011346199999999998 3.3 0.0011347199999999999 0 0.00113464 0 0.00113474 3.3 0.00113466 3.3 0.00113476 0 0.0011346799999999999 0 0.00113478 3.3 0.0011347 3.3 0.0011348 0 0.0011347199999999999 0 0.00113482 3.3 0.00113474 3.3 0.00113484 0 0.0011347599999999998 0 0.00113486 3.3 0.00113478 3.3 0.00113488 0 0.0011347999999999998 0 0.0011348999999999999 3.3 0.00113482 3.3 0.00113492 0 0.00113484 0 0.00113494 3.3 0.00113486 3.3 0.00113496 0 0.00113488 0 0.00113498 3.3 0.0011348999999999999 3.3 0.001135 0 0.00113492 0 0.00113502 3.3 0.0011349399999999999 3.3 0.00113504 0 0.00113496 0 0.00113506 3.3 0.0011349799999999998 3.3 0.00113508 0 0.001135 0 0.0011351 3.3 0.0011350199999999998 3.3 0.0011351199999999999 0 0.00113504 0 0.00113514 3.3 0.00113506 3.3 0.00113516 0 0.00113508 0 0.00113518 3.3 0.0011351 3.3 0.0011352 0 0.0011351199999999999 0 0.00113522 3.3 0.00113514 3.3 0.00113524 0 0.0011351599999999999 0 0.00113526 3.3 0.00113518 3.3 0.00113528 0 0.0011351999999999998 0 0.0011353 3.3 0.00113522 3.3 0.00113532 0 0.0011352399999999998 0 0.0011353399999999999 3.3 0.00113526 3.3 0.00113536 0 0.00113528 0 0.00113538 3.3 0.0011353 3.3 0.0011354 0 0.00113532 0 0.00113542 3.3 0.0011353399999999999 3.3 0.00113544 0 0.00113536 0 0.00113546 3.3 0.0011353799999999999 3.3 0.00113548 0 0.0011354 0 0.0011355 3.3 0.0011354199999999998 3.3 0.0011355199999999999 0 0.00113544 0 0.00113554 3.3 0.00113546 3.3 0.00113556 0 0.00113548 0 0.00113558 3.3 0.0011355 3.3 0.0011356 0 0.0011355199999999999 0 0.00113562 3.3 0.00113554 3.3 0.00113564 0 0.0011355599999999999 0 0.00113566 3.3 0.00113558 3.3 0.00113568 0 0.0011355999999999998 0 0.0011357 3.3 0.00113562 3.3 0.00113572 0 0.0011356399999999998 0 0.0011357399999999999 3.3 0.00113566 3.3 0.00113576 0 0.00113568 0 0.00113578 3.3 0.0011357 3.3 0.0011358 0 0.00113572 0 0.00113582 3.3 0.0011357399999999999 3.3 0.00113584 0 0.00113576 0 0.00113586 3.3 0.0011357799999999999 3.3 0.00113588 0 0.0011358 0 0.0011359 3.3 0.0011358199999999998 3.3 0.00113592 0 0.00113584 0 0.00113594 3.3 0.0011358599999999998 3.3 0.0011359599999999999 0 0.00113588 0 0.00113598 3.3 0.0011359 3.3 0.001136 0 0.00113592 0 0.00113602 3.3 0.00113594 3.3 0.00113604 0 0.0011359599999999999 0 0.00113606 3.3 0.00113598 3.3 0.00113608 0 0.0011359999999999999 0 0.0011361 3.3 0.00113602 3.3 0.00113612 0 0.0011360399999999998 0 0.00113614 3.3 0.00113606 3.3 0.00113616 0 0.0011360799999999998 0 0.0011361799999999999 3.3 0.0011361 3.3 0.0011362 0 0.00113612 0 0.00113622 3.3 0.00113614 3.3 0.00113624 0 0.00113616 0 0.00113626 3.3 0.0011361799999999999 3.3 0.00113628 0 0.0011362 0 0.0011363 3.3 0.0011362199999999999 3.3 0.00113632 0 0.00113624 0 0.00113634 3.3 0.0011362599999999998 3.3 0.0011363599999999999 0 0.00113628 0 0.00113638 3.3 0.0011363 3.3 0.0011364 0 0.00113632 0 0.00113642 3.3 0.00113634 3.3 0.00113644 0 0.0011363599999999999 0 0.00113646 3.3 0.00113638 3.3 0.00113648 0 0.0011363999999999999 0 0.0011365 3.3 0.00113642 3.3 0.00113652 0 0.0011364399999999998 0 0.00113654 3.3 0.00113646 3.3 0.00113656 0 0.0011364799999999998 0 0.0011365799999999999 3.3 0.0011365 3.3 0.0011366 0 0.00113652 0 0.00113662 3.3 0.00113654 3.3 0.00113664 0 0.00113656 0 0.00113666 3.3 0.0011365799999999999 3.3 0.00113668 0 0.0011366 0 0.0011367 3.3 0.0011366199999999999 3.3 0.00113672 0 0.00113664 0 0.00113674 3.3 0.0011366599999999998 3.3 0.00113676 0 0.00113668 0 0.00113678 3.3 0.0011366999999999998 3.3 0.0011367999999999999 0 0.00113672 0 0.00113682 3.3 0.00113674 3.3 0.00113684 0 0.00113676 0 0.00113686 3.3 0.00113678 3.3 0.00113688 0 0.0011367999999999999 0 0.0011369 3.3 0.00113682 3.3 0.00113692 0 0.0011368399999999999 0 0.00113694 3.3 0.00113686 3.3 0.00113696 0 0.0011368799999999998 0 0.00113698 3.3 0.0011369 3.3 0.001137 0 0.0011369199999999998 0 0.0011370199999999999 3.3 0.00113694 3.3 0.00113704 0 0.00113696 0 0.00113706 3.3 0.00113698 3.3 0.00113708 0 0.001137 0 0.0011371 3.3 0.0011370199999999999 3.3 0.00113712 0 0.00113704 0 0.00113714 3.3 0.0011370599999999999 3.3 0.00113716 0 0.00113708 0 0.00113718 3.3 0.0011370999999999998 3.3 0.0011371999999999999 0 0.00113712 0 0.00113722 3.3 0.00113714 3.3 0.00113724 0 0.00113716 0 0.00113726 3.3 0.00113718 3.3 0.00113728 0 0.0011371999999999999 0 0.0011373 3.3 0.00113722 3.3 0.00113732 0 0.0011372399999999999 0 0.00113734 3.3 0.00113726 3.3 0.00113736 0 0.0011372799999999998 0 0.00113738 3.3 0.0011373 3.3 0.0011374 0 0.0011373199999999998 0 0.0011374199999999999 3.3 0.00113734 3.3 0.00113744 0 0.00113736 0 0.00113746 3.3 0.00113738 3.3 0.00113748 0 0.0011374 0 0.0011375 3.3 0.0011374199999999999 3.3 0.00113752 0 0.00113744 0 0.00113754 3.3 0.0011374599999999999 3.3 0.00113756 0 0.00113748 0 0.00113758 3.3 0.0011374999999999998 3.3 0.0011376 0 0.00113752 0 0.00113762 3.3 0.0011375399999999998 3.3 0.0011376399999999999 0 0.00113756 0 0.00113766 3.3 0.00113758 3.3 0.00113768 0 0.0011376 0 0.0011377 3.3 0.00113762 3.3 0.00113772 0 0.0011376399999999999 0 0.00113774 3.3 0.00113766 3.3 0.00113776 0 0.0011376799999999999 0 0.00113778 3.3 0.0011377 3.3 0.0011378 0 0.0011377199999999998 0 0.0011378199999999999 3.3 0.00113774 3.3 0.00113784 0 0.0011377599999999998 0 0.0011378599999999999 3.3 0.00113778 3.3 0.00113788 0 0.0011378 0 0.0011379 3.3 0.0011378199999999999 3.3 0.00113792 0 0.00113784 0 0.00113794 3.3 0.0011378599999999999 3.3 0.00113796 0 0.00113788 0 0.00113798 3.3 0.0011378999999999998 3.3 0.001138 0 0.00113792 0 0.00113802 3.3 0.0011379399999999998 3.3 0.0011380399999999999 0 0.00113796 0 0.00113806 3.3 0.00113798 3.3 0.00113808 0 0.001138 0 0.0011381 3.3 0.00113802 3.3 0.00113812 0 0.0011380399999999999 0 0.00113814 3.3 0.00113806 3.3 0.00113816 0 0.0011380799999999999 0 0.00113818 3.3 0.0011381 3.3 0.0011382 0 0.0011381199999999998 0 0.00113822 3.3 0.00113814 3.3 0.00113824 0 0.0011381599999999998 0 0.0011382599999999999 3.3 0.00113818 3.3 0.00113828 0 0.0011382 0 0.0011383 3.3 0.00113822 3.3 0.00113832 0 0.00113824 0 0.00113834 3.3 0.0011382599999999999 3.3 0.00113836 0 0.00113828 0 0.00113838 3.3 0.0011382999999999999 3.3 0.0011384 0 0.00113832 0 0.00113842 3.3 0.0011383399999999998 3.3 0.00113844 0 0.00113836 0 0.00113846 3.3 0.0011383799999999998 3.3 0.0011384799999999999 0 0.0011384 0 0.0011385 3.3 0.00113842 3.3 0.00113852 0 0.00113844 0 0.00113854 3.3 0.00113846 3.3 0.00113856 0 0.0011384799999999999 0 0.00113858 3.3 0.0011385 3.3 0.0011386 0 0.0011385199999999999 0 0.00113862 3.3 0.00113854 3.3 0.00113864 0 0.0011385599999999998 0 0.0011386599999999999 3.3 0.00113858 3.3 0.00113868 0 0.0011386 0 0.0011387 3.3 0.00113862 3.3 0.00113872 0 0.00113864 0 0.00113874 3.3 0.0011386599999999999 3.3 0.00113876 0 0.00113868 0 0.00113878 3.3 0.0011386999999999999 3.3 0.0011388 0 0.00113872 0 0.00113882 3.3 0.0011387399999999998 3.3 0.00113884 0 0.00113876 0 0.00113886 3.3 0.0011387799999999998 3.3 0.0011388799999999999 0 0.0011388 0 0.0011389 3.3 0.00113882 3.3 0.00113892 0 0.00113884 0 0.00113894 3.3 0.00113886 3.3 0.00113896 0 0.0011388799999999999 0 0.00113898 3.3 0.0011389 3.3 0.001139 0 0.0011389199999999999 0 0.00113902 3.3 0.00113894 3.3 0.00113904 0 0.0011389599999999998 0 0.00113906 3.3 0.00113898 3.3 0.00113908 0 0.0011389999999999998 0 0.0011390999999999999 3.3 0.00113902 3.3 0.00113912 0 0.00113904 0 0.00113914 3.3 0.00113906 3.3 0.00113916 0 0.00113908 0 0.00113918 3.3 0.0011390999999999999 3.3 0.0011392 0 0.00113912 0 0.00113922 3.3 0.0011391399999999999 3.3 0.00113924 0 0.00113916 0 0.00113926 3.3 0.0011391799999999998 3.3 0.00113928 0 0.0011392 0 0.0011393 3.3 0.0011392199999999998 3.3 0.0011393199999999999 0 0.00113924 0 0.00113934 3.3 0.00113926 3.3 0.00113936 0 0.00113928 0 0.00113938 3.3 0.0011393 3.3 0.0011394 0 0.0011393199999999999 0 0.00113942 3.3 0.00113934 3.3 0.00113944 0 0.0011393599999999999 0 0.00113946 3.3 0.00113938 3.3 0.00113948 0 0.0011393999999999998 0 0.0011394999999999999 3.3 0.00113942 3.3 0.00113952 0 0.00113944 0 0.00113954 3.3 0.00113946 3.3 0.00113956 0 0.00113948 0 0.00113958 3.3 0.0011394999999999999 3.3 0.0011396 0 0.00113952 0 0.00113962 3.3 0.0011395399999999999 3.3 0.00113964 0 0.00113956 0 0.00113966 3.3 0.0011395799999999998 3.3 0.00113968 0 0.0011396 0 0.0011397 3.3 0.0011396199999999998 3.3 0.0011397199999999999 0 0.00113964 0 0.00113974 3.3 0.00113966 3.3 0.00113976 0 0.00113968 0 0.00113978 3.3 0.0011397 3.3 0.0011398 0 0.0011397199999999999 0 0.00113982 3.3 0.00113974 3.3 0.00113984 0 0.0011397599999999999 0 0.00113986 3.3 0.00113978 3.3 0.00113988 0 0.0011397999999999998 0 0.0011399 3.3 0.00113982 3.3 0.00113992 0 0.0011398399999999998 0 0.0011399399999999999 3.3 0.00113986 3.3 0.00113996 0 0.00113988 0 0.00113998 3.3 0.0011399 3.3 0.00114 0 0.00113992 0 0.00114002 3.3 0.0011399399999999999 3.3 0.00114004 0 0.00113996 0 0.00114006 3.3 0.0011399799999999999 3.3 0.00114008 0 0.00114 0 0.0011401 3.3 0.0011400199999999998 3.3 0.00114012 0 0.00114004 0 0.00114014 3.3 0.0011400599999999998 3.3 0.0011401599999999999 0 0.00114008 0 0.00114018 3.3 0.0011401 3.3 0.0011402 0 0.00114012 0 0.00114022 3.3 0.00114014 3.3 0.00114024 0 0.0011401599999999999 0 0.00114026 3.3 0.00114018 3.3 0.00114028 0 0.0011401999999999999 0 0.0011403 3.3 0.00114022 3.3 0.00114032 0 0.0011402399999999998 0 0.0011403399999999999 3.3 0.00114026 3.3 0.00114036 0 0.00114028 0 0.00114038 3.3 0.0011403 3.3 0.0011404 0 0.00114032 0 0.00114042 3.3 0.0011403399999999999 3.3 0.00114044 0 0.00114036 0 0.00114046 3.3 0.0011403799999999999 3.3 0.00114048 0 0.0011404 0 0.0011405 3.3 0.0011404199999999998 3.3 0.00114052 0 0.00114044 0 0.00114054 3.3 0.0011404599999999998 3.3 0.0011405599999999999 0 0.00114048 0 0.00114058 3.3 0.0011405 3.3 0.0011406 0 0.00114052 0 0.00114062 3.3 0.00114054 3.3 0.00114064 0 0.0011405599999999999 0 0.00114066 3.3 0.00114058 3.3 0.00114068 0 0.0011405999999999999 0 0.0011407 3.3 0.00114062 3.3 0.00114072 0 0.0011406399999999998 0 0.00114074 3.3 0.00114066 3.3 0.00114076 0 0.0011406799999999998 0 0.0011407799999999999 3.3 0.0011407 3.3 0.0011408 0 0.00114072 0 0.00114082 3.3 0.00114074 3.3 0.00114084 0 0.00114076 0 0.00114086 3.3 0.0011407799999999999 3.3 0.00114088 0 0.0011408 0 0.0011409 3.3 0.0011408199999999999 3.3 0.00114092 0 0.00114084 0 0.00114094 3.3 0.0011408599999999998 3.3 0.0011409599999999999 0 0.00114088 0 0.00114098 3.3 0.0011408999999999998 3.3 0.0011409999999999999 0 0.00114092 0 0.00114102 3.3 0.00114094 3.3 0.00114104 0 0.0011409599999999999 0 0.00114106 3.3 0.00114098 3.3 0.00114108 0 0.0011409999999999999 0 0.0011411 3.3 0.00114102 3.3 0.00114112 0 0.0011410399999999998 0 0.00114114 3.3 0.00114106 3.3 0.00114116 0 0.0011410799999999998 0 0.0011411799999999999 3.3 0.0011411 3.3 0.0011412 0 0.00114112 0 0.00114122 3.3 0.00114114 3.3 0.00114124 0 0.00114116 0 0.00114126 3.3 0.0011411799999999999 3.3 0.00114128 0 0.0011412 0 0.0011413 3.3 0.0011412199999999999 3.3 0.00114132 0 0.00114124 0 0.00114134 3.3 0.0011412599999999998 3.3 0.00114136 0 0.00114128 0 0.00114138 3.3 0.0011412999999999998 3.3 0.0011413999999999999 0 0.00114132 0 0.00114142 3.3 0.00114134 3.3 0.00114144 0 0.00114136 0 0.00114146 3.3 0.00114138 3.3 0.00114148 0 0.0011413999999999999 0 0.0011415 3.3 0.00114142 3.3 0.00114152 0 0.0011414399999999999 0 0.00114154 3.3 0.00114146 3.3 0.00114156 0 0.0011414799999999998 0 0.00114158 3.3 0.0011415 3.3 0.0011416 0 0.0011415199999999998 0 0.0011416199999999999 3.3 0.00114154 3.3 0.00114164 0 0.00114156 0 0.00114166 3.3 0.00114158 3.3 0.00114168 0 0.0011416 0 0.0011417 3.3 0.0011416199999999999 3.3 0.00114172 0 0.00114164 0 0.00114174 3.3 0.0011416599999999999 3.3 0.00114176 0 0.00114168 0 0.00114178 3.3 0.0011416999999999998 3.3 0.0011417999999999999 0 0.00114172 0 0.00114182 3.3 0.0011417399999999998 3.3 0.0011418399999999999 0 0.00114176 0 0.00114186 3.3 0.00114178 3.3 0.00114188 0 0.0011417999999999999 0 0.0011419 3.3 0.00114182 3.3 0.00114192 0 0.0011418399999999999 0 0.00114194 3.3 0.00114186 3.3 0.00114196 0 0.0011418799999999998 0 0.00114198 3.3 0.0011419 3.3 0.001142 0 0.0011419199999999998 0 0.0011420199999999999 3.3 0.00114194 3.3 0.00114204 0 0.00114196 0 0.00114206 3.3 0.00114198 3.3 0.00114208 0 0.001142 0 0.0011421 3.3 0.0011420199999999999 3.3 0.00114212 0 0.00114204 0 0.00114214 3.3 0.0011420599999999999 3.3 0.00114216 0 0.00114208 0 0.00114218 3.3 0.0011420999999999998 3.3 0.0011422 0 0.00114212 0 0.00114222 3.3 0.0011421399999999998 3.3 0.0011422399999999999 0 0.00114216 0 0.00114226 3.3 0.00114218 3.3 0.00114228 0 0.0011422 0 0.0011423 3.3 0.00114222 3.3 0.00114232 0 0.0011422399999999999 0 0.00114234 3.3 0.00114226 3.3 0.00114236 0 0.0011422799999999999 0 0.00114238 3.3 0.0011423 3.3 0.0011424 0 0.0011423199999999998 0 0.00114242 3.3 0.00114234 3.3 0.00114244 0 0.0011423599999999998 0 0.0011424599999999999 3.3 0.00114238 3.3 0.00114248 0 0.0011424 0 0.0011425 3.3 0.00114242 3.3 0.00114252 0 0.00114244 0 0.00114254 3.3 0.0011424599999999999 3.3 0.00114256 0 0.00114248 0 0.00114258 3.3 0.0011424999999999999 3.3 0.0011426 0 0.00114252 0 0.00114262 3.3 0.0011425399999999998 3.3 0.0011426399999999999 0 0.00114256 0 0.00114266 3.3 0.00114258 3.3 0.00114268 0 0.0011426 0 0.0011427 3.3 0.00114262 3.3 0.00114272 0 0.0011426399999999999 0 0.00114274 3.3 0.00114266 3.3 0.00114276 0 0.0011426799999999999 0 0.00114278 3.3 0.0011427 3.3 0.0011428 0 0.0011427199999999998 0 0.00114282 3.3 0.00114274 3.3 0.00114284 0 0.0011427599999999998 0 0.0011428599999999999 3.3 0.00114278 3.3 0.00114288 0 0.0011428 0 0.0011429 3.3 0.00114282 3.3 0.00114292 0 0.00114284 0 0.00114294 3.3 0.0011428599999999999 3.3 0.00114296 0 0.00114288 0 0.00114298 3.3 0.0011428999999999999 3.3 0.001143 0 0.00114292 0 0.00114302 3.3 0.0011429399999999998 3.3 0.00114304 0 0.00114296 0 0.00114306 3.3 0.0011429799999999998 3.3 0.0011430799999999999 0 0.001143 0 0.0011431 3.3 0.00114302 3.3 0.00114312 0 0.00114304 0 0.00114314 3.3 0.00114306 3.3 0.00114316 0 0.0011430799999999999 0 0.00114318 3.3 0.0011431 3.3 0.0011432 0 0.0011431199999999999 0 0.00114322 3.3 0.00114314 3.3 0.00114324 0 0.0011431599999999998 0 0.00114326 3.3 0.00114318 3.3 0.00114328 0 0.0011431999999999998 0 0.0011432999999999999 3.3 0.00114322 3.3 0.00114332 0 0.00114324 0 0.00114334 3.3 0.00114326 3.3 0.00114336 0 0.00114328 0 0.00114338 3.3 0.0011432999999999999 3.3 0.0011434 0 0.00114332 0 0.00114342 3.3 0.0011433399999999999 3.3 0.00114344 0 0.00114336 0 0.00114346 3.3 0.0011433799999999998 3.3 0.0011434799999999999 0 0.0011434 0 0.0011435 3.3 0.00114342 3.3 0.00114352 0 0.00114344 0 0.00114354 3.3 0.00114346 3.3 0.00114356 0 0.0011434799999999999 0 0.00114358 3.3 0.0011435 3.3 0.0011436 0 0.0011435199999999999 0 0.00114362 3.3 0.00114354 3.3 0.00114364 0 0.0011435599999999998 0 0.00114366 3.3 0.00114358 3.3 0.00114368 0 0.0011435999999999998 0 0.0011436999999999999 3.3 0.00114362 3.3 0.00114372 0 0.00114364 0 0.00114374 3.3 0.00114366 3.3 0.00114376 0 0.00114368 0 0.00114378 3.3 0.0011436999999999999 3.3 0.0011438 0 0.00114372 0 0.00114382 3.3 0.0011437399999999999 3.3 0.00114384 0 0.00114376 0 0.00114386 3.3 0.0011437799999999998 3.3 0.00114388 0 0.0011438 0 0.0011439 3.3 0.0011438199999999998 3.3 0.0011439199999999999 0 0.00114384 0 0.00114394 3.3 0.00114386 3.3 0.00114396 0 0.00114388 0 0.00114398 3.3 0.0011439 3.3 0.001144 0 0.0011439199999999999 0 0.00114402 3.3 0.00114394 3.3 0.00114404 0 0.0011439599999999999 0 0.00114406 3.3 0.00114398 3.3 0.00114408 0 0.0011439999999999998 0 0.0011440999999999999 3.3 0.00114402 3.3 0.00114412 0 0.0011440399999999998 0 0.0011441399999999999 3.3 0.00114406 3.3 0.00114416 0 0.00114408 0 0.00114418 3.3 0.0011440999999999999 3.3 0.0011442 0 0.00114412 0 0.00114422 3.3 0.0011441399999999999 3.3 0.00114424 0 0.00114416 0 0.00114426 3.3 0.0011441799999999998 3.3 0.00114428 0 0.0011442 0 0.0011443 3.3 0.0011442199999999998 3.3 0.0011443199999999999 0 0.00114424 0 0.00114434 3.3 0.00114426 3.3 0.00114436 0 0.00114428 0 0.00114438 3.3 0.0011443 3.3 0.0011444 0 0.0011443199999999999 0 0.00114442 3.3 0.00114434 3.3 0.00114444 0 0.0011443599999999999 0 0.00114446 3.3 0.00114438 3.3 0.00114448 0 0.0011443999999999998 0 0.0011445 3.3 0.00114442 3.3 0.00114452 0 0.0011444399999999998 0 0.0011445399999999999 3.3 0.00114446 3.3 0.00114456 0 0.00114448 0 0.00114458 3.3 0.0011445 3.3 0.0011446 0 0.00114452 0 0.00114462 3.3 0.0011445399999999999 3.3 0.00114464 0 0.00114456 0 0.00114466 3.3 0.0011445799999999999 3.3 0.00114468 0 0.0011446 0 0.0011447 3.3 0.0011446199999999998 3.3 0.00114472 0 0.00114464 0 0.00114474 3.3 0.0011446599999999998 3.3 0.0011447599999999999 0 0.00114468 0 0.00114478 3.3 0.0011447 3.3 0.0011448 0 0.00114472 0 0.00114482 3.3 0.00114474 3.3 0.00114484 0 0.0011447599999999999 0 0.00114486 3.3 0.00114478 3.3 0.00114488 0 0.0011447999999999999 0 0.0011449 3.3 0.00114482 3.3 0.00114492 0 0.0011448399999999998 0 0.0011449399999999999 3.3 0.00114486 3.3 0.00114496 0 0.0011448799999999998 0 0.0011449799999999999 3.3 0.0011449 3.3 0.001145 0 0.00114492 0 0.00114502 3.3 0.0011449399999999999 3.3 0.00114504 0 0.00114496 0 0.00114506 3.3 0.0011449799999999999 3.3 0.00114508 0 0.001145 0 0.0011451 3.3 0.0011450199999999998 3.3 0.00114512 0 0.00114504 0 0.00114514 3.3 0.0011450599999999998 3.3 0.0011451599999999999 0 0.00114508 0 0.00114518 3.3 0.0011451 3.3 0.0011452 0 0.00114512 0 0.00114522 3.3 0.00114514 3.3 0.00114524 0 0.0011451599999999999 0 0.00114526 3.3 0.00114518 3.3 0.00114528 0 0.0011451999999999999 0 0.0011453 3.3 0.00114522 3.3 0.00114532 0 0.0011452399999999998 0 0.00114534 3.3 0.00114526 3.3 0.00114536 0 0.0011452799999999998 0 0.0011453799999999999 3.3 0.0011453 3.3 0.0011454 0 0.00114532 0 0.00114542 3.3 0.00114534 3.3 0.00114544 0 0.00114536 0 0.00114546 3.3 0.0011453799999999999 3.3 0.00114548 0 0.0011454 0 0.0011455 3.3 0.0011454199999999999 3.3 0.00114552 0 0.00114544 0 0.00114554 3.3 0.0011454599999999998 3.3 0.00114556 0 0.00114548 0 0.00114558 3.3 0.0011454999999999998 3.3 0.0011455999999999999 0 0.00114552 0 0.00114562 3.3 0.00114554 3.3 0.00114564 0 0.00114556 0 0.00114566 3.3 0.00114558 3.3 0.00114568 0 0.0011455999999999999 0 0.0011457 3.3 0.00114562 3.3 0.00114572 0 0.0011456399999999999 0 0.00114574 3.3 0.00114566 3.3 0.00114576 0 0.0011456799999999998 0 0.0011457799999999999 3.3 0.0011457 3.3 0.0011458 0 0.00114572 0 0.00114582 3.3 0.00114574 3.3 0.00114584 0 0.00114576 0 0.00114586 3.3 0.0011457799999999999 3.3 0.00114588 0 0.0011458 0 0.0011459 3.3 0.0011458199999999999 3.3 0.00114592 0 0.00114584 0 0.00114594 3.3 0.0011458599999999998 3.3 0.00114596 0 0.00114588 0 0.00114598 3.3 0.0011458999999999998 3.3 0.0011459999999999999 0 0.00114592 0 0.00114602 3.3 0.00114594 3.3 0.00114604 0 0.00114596 0 0.00114606 3.3 0.00114598 3.3 0.00114608 0 0.0011459999999999999 0 0.0011461 3.3 0.00114602 3.3 0.00114612 0 0.0011460399999999999 0 0.00114614 3.3 0.00114606 3.3 0.00114616 0 0.0011460799999999998 0 0.00114618 3.3 0.0011461 3.3 0.0011462 0 0.0011461199999999998 0 0.0011462199999999999 3.3 0.00114614 3.3 0.00114624 0 0.00114616 0 0.00114626 3.3 0.00114618 3.3 0.00114628 0 0.0011462 0 0.0011463 3.3 0.0011462199999999999 3.3 0.00114632 0 0.00114624 0 0.00114634 3.3 0.0011462599999999999 3.3 0.00114636 0 0.00114628 0 0.00114638 3.3 0.0011462999999999998 3.3 0.0011464 0 0.00114632 0 0.00114642 3.3 0.0011463399999999998 3.3 0.0011464399999999999 0 0.00114636 0 0.00114646 3.3 0.00114638 3.3 0.00114648 0 0.0011464 0 0.0011465 3.3 0.00114642 3.3 0.00114652 0 0.0011464399999999999 0 0.00114654 3.3 0.00114646 3.3 0.00114656 0 0.0011464799999999999 0 0.00114658 3.3 0.0011465 3.3 0.0011466 0 0.0011465199999999998 0 0.0011466199999999999 3.3 0.00114654 3.3 0.00114664 0 0.00114656 0 0.00114666 3.3 0.00114658 3.3 0.00114668 0 0.0011466 0 0.0011467 3.3 0.0011466199999999999 3.3 0.00114672 0 0.00114664 0 0.00114674 3.3 0.0011466599999999999 3.3 0.00114676 0 0.00114668 0 0.00114678 3.3 0.0011466999999999998 3.3 0.0011468 0 0.00114672 0 0.00114682 3.3 0.0011467399999999998 3.3 0.0011468399999999999 0 0.00114676 0 0.00114686 3.3 0.00114678 3.3 0.00114688 0 0.0011468 0 0.0011469 3.3 0.00114682 3.3 0.00114692 0 0.0011468399999999999 0 0.00114694 3.3 0.00114686 3.3 0.00114696 0 0.0011468799999999999 0 0.00114698 3.3 0.0011469 3.3 0.001147 0 0.0011469199999999998 0 0.00114702 3.3 0.00114694 3.3 0.00114704 0 0.0011469599999999998 0 0.0011470599999999999 3.3 0.00114698 3.3 0.00114708 0 0.001147 0 0.0011471 3.3 0.00114702 3.3 0.00114712 0 0.00114704 0 0.00114714 3.3 0.0011470599999999999 3.3 0.00114716 0 0.00114708 0 0.00114718 3.3 0.0011470999999999999 3.3 0.0011472 0 0.00114712 0 0.00114722 3.3 0.0011471399999999998 3.3 0.00114724 0 0.00114716 0 0.00114726 3.3 0.0011471799999999998 3.3 0.0011472799999999999 0 0.0011472 0 0.0011473 3.3 0.00114722 3.3 0.00114732 0 0.00114724 0 0.00114734 3.3 0.00114726 3.3 0.00114736 0 0.0011472799999999999 0 0.00114738 3.3 0.0011473 3.3 0.0011474 0 0.0011473199999999999 0 0.00114742 3.3 0.00114734 3.3 0.00114744 0 0.0011473599999999998 0 0.0011474599999999999 3.3 0.00114738 3.3 0.00114748 0 0.0011474 0 0.0011475 3.3 0.00114742 3.3 0.00114752 0 0.00114744 0 0.00114754 3.3 0.0011474599999999999 3.3 0.00114756 0 0.00114748 0 0.00114758 3.3 0.0011474999999999999 3.3 0.0011476 0 0.00114752 0 0.00114762 3.3 0.0011475399999999998 3.3 0.00114764 0 0.00114756 0 0.00114766 3.3 0.0011475799999999998 3.3 0.0011476799999999999 0 0.0011476 0 0.0011477 3.3 0.00114762 3.3 0.00114772 0 0.00114764 0 0.00114774 3.3 0.00114766 3.3 0.00114776 0 0.0011476799999999999 0 0.00114778 3.3 0.0011477 3.3 0.0011478 0 0.0011477199999999999 0 0.00114782 3.3 0.00114774 3.3 0.00114784 0 0.0011477599999999998 0 0.00114786 3.3 0.00114778 3.3 0.00114788 0 0.0011477999999999998 0 0.0011478999999999999 3.3 0.00114782 3.3 0.00114792 0 0.00114784 0 0.00114794 3.3 0.00114786 3.3 0.00114796 0 0.00114788 0 0.00114798 3.3 0.0011478999999999999 3.3 0.001148 0 0.00114792 0 0.00114802 3.3 0.0011479399999999999 3.3 0.00114804 0 0.00114796 0 0.00114806 3.3 0.0011479799999999998 3.3 0.0011480799999999999 0 0.001148 0 0.0011481 3.3 0.0011480199999999998 3.3 0.0011481199999999999 0 0.00114804 0 0.00114814 3.3 0.00114806 3.3 0.00114816 0 0.0011480799999999999 0 0.00114818 3.3 0.0011481 3.3 0.0011482 0 0.0011481199999999999 0 0.00114822 3.3 0.00114814 3.3 0.00114824 0 0.0011481599999999998 0 0.00114826 3.3 0.00114818 3.3 0.00114828 0 0.0011481999999999998 0 0.0011482999999999999 3.3 0.00114822 3.3 0.00114832 0 0.00114824 0 0.00114834 3.3 0.00114826 3.3 0.00114836 0 0.00114828 0 0.00114838 3.3 0.0011482999999999999 3.3 0.0011484 0 0.00114832 0 0.00114842 3.3 0.0011483399999999999 3.3 0.00114844 0 0.00114836 0 0.00114846 3.3 0.0011483799999999998 3.3 0.00114848 0 0.0011484 0 0.0011485 3.3 0.0011484199999999998 3.3 0.0011485199999999999 0 0.00114844 0 0.00114854 3.3 0.00114846 3.3 0.00114856 0 0.00114848 0 0.00114858 3.3 0.0011485 3.3 0.0011486 0 0.0011485199999999999 0 0.00114862 3.3 0.00114854 3.3 0.00114864 0 0.0011485599999999999 0 0.00114866 3.3 0.00114858 3.3 0.00114868 0 0.0011485999999999998 0 0.0011487 3.3 0.00114862 3.3 0.00114872 0 0.0011486399999999998 0 0.0011487399999999999 3.3 0.00114866 3.3 0.00114876 0 0.00114868 0 0.00114878 3.3 0.0011487 3.3 0.0011488 0 0.00114872 0 0.00114882 3.3 0.0011487399999999999 3.3 0.00114884 0 0.00114876 0 0.00114886 3.3 0.0011487799999999999 3.3 0.00114888 0 0.0011488 0 0.0011489 3.3 0.0011488199999999998 3.3 0.0011489199999999999 0 0.00114884 0 0.00114894 3.3 0.0011488599999999998 3.3 0.0011489599999999999 0 0.00114888 0 0.00114898 3.3 0.0011489 3.3 0.001149 0 0.0011489199999999999 0 0.00114902 3.3 0.00114894 3.3 0.00114904 0 0.0011489599999999999 0 0.00114906 3.3 0.00114898 3.3 0.00114908 0 0.0011489999999999998 0 0.0011491 3.3 0.00114902 3.3 0.00114912 0 0.0011490399999999998 0 0.0011491399999999999 3.3 0.00114906 3.3 0.00114916 0 0.00114908 0 0.00114918 3.3 0.0011491 3.3 0.0011492 0 0.00114912 0 0.00114922 3.3 0.0011491399999999999 3.3 0.00114924 0 0.00114916 0 0.00114926 3.3 0.0011491799999999999 3.3 0.00114928 0 0.0011492 0 0.0011493 3.3 0.0011492199999999998 3.3 0.00114932 0 0.00114924 0 0.00114934 3.3 0.0011492599999999998 3.3 0.0011493599999999999 0 0.00114928 0 0.00114938 3.3 0.0011493 3.3 0.0011494 0 0.00114932 0 0.00114942 3.3 0.00114934 3.3 0.00114944 0 0.0011493599999999999 0 0.00114946 3.3 0.00114938 3.3 0.00114948 0 0.0011493999999999999 0 0.0011495 3.3 0.00114942 3.3 0.00114952 0 0.0011494399999999998 0 0.00114954 3.3 0.00114946 3.3 0.00114956 0 0.0011494799999999998 0 0.0011495799999999999 3.3 0.0011495 3.3 0.0011496 0 0.00114952 0 0.00114962 3.3 0.00114954 3.3 0.00114964 0 0.00114956 0 0.00114966 3.3 0.0011495799999999999 3.3 0.00114968 0 0.0011496 0 0.0011497 3.3 0.0011496199999999999 3.3 0.00114972 0 0.00114964 0 0.00114974 3.3 0.0011496599999999998 3.3 0.0011497599999999999 0 0.00114968 0 0.00114978 3.3 0.0011497 3.3 0.0011498 0 0.00114972 0 0.00114982 3.3 0.00114974 3.3 0.00114984 0 0.0011497599999999999 0 0.00114986 3.3 0.00114978 3.3 0.00114988 0 0.0011497999999999999 0 0.0011499 3.3 0.00114982 3.3 0.00114992 0 0.0011498399999999998 0 0.00114994 3.3 0.00114986 3.3 0.00114996 0 0.0011498799999999998 0 0.0011499799999999999 3.3 0.0011499 3.3 0.00115 0 0.00114992 0 0.00115002 3.3 0.00114994 3.3 0.00115004 0 0.00114996 0 0.00115006 3.3 0.0011499799999999999 3.3 0.00115008 0 0.00115 0 0.0011501 3.3 0.0011500199999999999 3.3 0.00115012 0 0.00115004 0 0.00115014 3.3 0.0011500599999999998 3.3 0.00115016 0 0.00115008 0 0.00115018 3.3 0.0011500999999999998 3.3 0.0011501999999999999 0 0.00115012 0 0.00115022 3.3 0.00115014 3.3 0.00115024 0 0.00115016 0 0.00115026 3.3 0.00115018 3.3 0.00115028 0 0.0011501999999999999 0 0.0011503 3.3 0.00115022 3.3 0.00115032 0 0.0011502399999999999 0 0.00115034 3.3 0.00115026 3.3 0.00115036 0 0.0011502799999999998 0 0.00115038 3.3 0.0011503 3.3 0.0011504 0 0.0011503199999999998 0 0.0011504199999999999 3.3 0.00115034 3.3 0.00115044 0 0.00115036 0 0.00115046 3.3 0.00115038 3.3 0.00115048 0 0.0011504 0 0.0011505 3.3 0.0011504199999999999 3.3 0.00115052 0 0.00115044 0 0.00115054 3.3 0.0011504599999999999 3.3 0.00115056 0 0.00115048 0 0.00115058 3.3 0.0011504999999999998 3.3 0.0011505999999999999 0 0.00115052 0 0.00115062 3.3 0.00115054 3.3 0.00115064 0 0.00115056 0 0.00115066 3.3 0.00115058 3.3 0.00115068 0 0.0011505999999999999 0 0.0011507 3.3 0.00115062 3.3 0.00115072 0 0.0011506399999999999 0 0.00115074 3.3 0.00115066 3.3 0.00115076 0 0.0011506799999999998 0 0.00115078 3.3 0.0011507 3.3 0.0011508 0 0.0011507199999999998 0 0.0011508199999999999 3.3 0.00115074 3.3 0.00115084 0 0.00115076 0 0.00115086 3.3 0.00115078 3.3 0.00115088 0 0.0011508 0 0.0011509 3.3 0.0011508199999999999 3.3 0.00115092 0 0.00115084 0 0.00115094 3.3 0.0011508599999999999 3.3 0.00115096 0 0.00115088 0 0.00115098 3.3 0.0011508999999999998 3.3 0.001151 0 0.00115092 0 0.00115102 3.3 0.0011509399999999998 3.3 0.0011510399999999999 0 0.00115096 0 0.00115106 3.3 0.00115098 3.3 0.00115108 0 0.001151 0 0.0011511 3.3 0.00115102 3.3 0.00115112 0 0.0011510399999999999 0 0.00115114 3.3 0.00115106 3.3 0.00115116 0 0.0011510799999999999 0 0.00115118 3.3 0.0011511 3.3 0.0011512 0 0.0011511199999999998 0 0.0011512199999999999 3.3 0.00115114 3.3 0.00115124 0 0.0011511599999999998 0 0.0011512599999999999 3.3 0.00115118 3.3 0.00115128 0 0.0011512 0 0.0011513 3.3 0.0011512199999999999 3.3 0.00115132 0 0.00115124 0 0.00115134 3.3 0.0011512599999999999 3.3 0.00115136 0 0.00115128 0 0.00115138 3.3 0.0011512999999999998 3.3 0.0011514 0 0.00115132 0 0.00115142 3.3 0.0011513399999999998 3.3 0.0011514399999999999 0 0.00115136 0 0.00115146 3.3 0.00115138 3.3 0.00115148 0 0.0011514 0 0.0011515 3.3 0.00115142 3.3 0.00115152 0 0.0011514399999999999 0 0.00115154 3.3 0.00115146 3.3 0.00115156 0 0.0011514799999999999 0 0.00115158 3.3 0.0011515 3.3 0.0011516 0 0.0011515199999999998 0 0.00115162 3.3 0.00115154 3.3 0.00115164 0 0.0011515599999999998 0 0.0011516599999999999 3.3 0.00115158 3.3 0.00115168 0 0.0011516 0 0.0011517 3.3 0.00115162 3.3 0.00115172 0 0.00115164 0 0.00115174 3.3 0.0011516599999999999 3.3 0.00115176 0 0.00115168 0 0.00115178 3.3 0.0011516999999999999 3.3 0.0011518 0 0.00115172 0 0.00115182 3.3 0.0011517399999999998 3.3 0.00115184 0 0.00115176 0 0.00115186 3.3 0.0011517799999999998 3.3 0.0011518799999999999 0 0.0011518 0 0.0011519 3.3 0.00115182 3.3 0.00115192 0 0.00115184 0 0.00115194 3.3 0.00115186 3.3 0.00115196 0 0.0011518799999999999 0 0.00115198 3.3 0.0011519 3.3 0.001152 0 0.0011519199999999999 0 0.00115202 3.3 0.00115194 3.3 0.00115204 0 0.0011519599999999998 0 0.0011520599999999999 3.3 0.00115198 3.3 0.00115208 0 0.0011519999999999998 0 0.0011520999999999999 3.3 0.00115202 3.3 0.00115212 0 0.00115204 0 0.00115214 3.3 0.0011520599999999999 3.3 0.00115216 0 0.00115208 0 0.00115218 3.3 0.0011520999999999999 3.3 0.0011522 0 0.00115212 0 0.00115222 3.3 0.0011521399999999998 3.3 0.00115224 0 0.00115216 0 0.00115226 3.3 0.0011521799999999998 3.3 0.0011522799999999999 0 0.0011522 0 0.0011523 3.3 0.00115222 3.3 0.00115232 0 0.00115224 0 0.00115234 3.3 0.00115226 3.3 0.00115236 0 0.0011522799999999999 0 0.00115238 3.3 0.0011523 3.3 0.0011524 0 0.0011523199999999999 0 0.00115242 3.3 0.00115234 3.3 0.00115244 0 0.0011523599999999998 0 0.00115246 3.3 0.00115238 3.3 0.00115248 0 0.0011523999999999998 0 0.0011524999999999999 3.3 0.00115242 3.3 0.00115252 0 0.00115244 0 0.00115254 3.3 0.00115246 3.3 0.00115256 0 0.00115248 0 0.00115258 3.3 0.0011524999999999999 3.3 0.0011526 0 0.00115252 0 0.00115262 3.3 0.0011525399999999999 3.3 0.00115264 0 0.00115256 0 0.00115266 3.3 0.0011525799999999998 3.3 0.00115268 0 0.0011526 0 0.0011527 3.3 0.0011526199999999998 3.3 0.0011527199999999999 0 0.00115264 0 0.00115274 3.3 0.00115266 3.3 0.00115276 0 0.00115268 0 0.00115278 3.3 0.0011527 3.3 0.0011528 0 0.0011527199999999999 0 0.00115282 3.3 0.00115274 3.3 0.00115284 0 0.0011527599999999999 0 0.00115286 3.3 0.00115278 3.3 0.00115288 0 0.0011527999999999998 0 0.0011528999999999999 3.3 0.00115282 3.3 0.00115292 0 0.00115284 0 0.00115294 3.3 0.00115286 3.3 0.00115296 0 0.00115288 0 0.00115298 3.3 0.0011528999999999999 3.3 0.001153 0 0.00115292 0 0.00115302 3.3 0.0011529399999999999 3.3 0.00115304 0 0.00115296 0 0.00115306 3.3 0.0011529799999999998 3.3 0.00115308 0 0.001153 0 0.0011531 3.3 0.0011530199999999998 3.3 0.0011531199999999999 0 0.00115304 0 0.00115314 3.3 0.00115306 3.3 0.00115316 0 0.00115308 0 0.00115318 3.3 0.0011531 3.3 0.0011532 0 0.0011531199999999999 0 0.00115322 3.3 0.00115314 3.3 0.00115324 0 0.0011531599999999999 0 0.00115326 3.3 0.00115318 3.3 0.00115328 0 0.0011531999999999998 0 0.0011533 3.3 0.00115322 3.3 0.00115332 0 0.0011532399999999998 0 0.0011533399999999999 3.3 0.00115326 3.3 0.00115336 0 0.00115328 0 0.00115338 3.3 0.0011533 3.3 0.0011534 0 0.00115332 0 0.00115342 3.3 0.0011533399999999999 3.3 0.00115344 0 0.00115336 0 0.00115346 3.3 0.0011533799999999999 3.3 0.00115348 0 0.0011534 0 0.0011535 3.3 0.0011534199999999998 3.3 0.00115352 0 0.00115344 0 0.00115354 3.3 0.0011534599999999998 3.3 0.0011535599999999999 0 0.00115348 0 0.00115358 3.3 0.0011535 3.3 0.0011536 0 0.00115352 0 0.00115362 3.3 0.00115354 3.3 0.00115364 0 0.0011535599999999999 0 0.00115366 3.3 0.00115358 3.3 0.00115368 0 0.0011535999999999999 0 0.0011537 3.3 0.00115362 3.3 0.00115372 0 0.0011536399999999998 0 0.0011537399999999999 3.3 0.00115366 3.3 0.00115376 0 0.00115368 0 0.00115378 3.3 0.0011537 3.3 0.0011538 0 0.00115372 0 0.00115382 3.3 0.0011537399999999999 3.3 0.00115384 0 0.00115376 0 0.00115386 3.3 0.0011537799999999999 3.3 0.00115388 0 0.0011538 0 0.0011539 3.3 0.0011538199999999998 3.3 0.00115392 0 0.00115384 0 0.00115394 3.3 0.0011538599999999998 3.3 0.0011539599999999999 0 0.00115388 0 0.00115398 3.3 0.0011539 3.3 0.001154 0 0.00115392 0 0.00115402 3.3 0.00115394 3.3 0.00115404 0 0.0011539599999999999 0 0.00115406 3.3 0.00115398 3.3 0.00115408 0 0.0011539999999999999 0 0.0011541 3.3 0.00115402 3.3 0.00115412 0 0.0011540399999999998 0 0.00115414 3.3 0.00115406 3.3 0.00115416 0 0.0011540799999999998 0 0.0011541799999999999 3.3 0.0011541 3.3 0.0011542 0 0.00115412 0 0.00115422 3.3 0.00115414 3.3 0.00115424 0 0.00115416 0 0.00115426 3.3 0.0011541799999999999 3.3 0.00115428 0 0.0011542 0 0.0011543 3.3 0.0011542199999999999 3.3 0.00115432 0 0.00115424 0 0.00115434 3.3 0.0011542599999999998 3.3 0.0011543599999999999 0 0.00115428 0 0.00115438 3.3 0.0011542999999999998 3.3 0.0011543999999999999 0 0.00115432 0 0.00115442 3.3 0.00115434 3.3 0.00115444 0 0.0011543599999999999 0 0.00115446 3.3 0.00115438 3.3 0.00115448 0 0.0011543999999999999 0 0.0011545 3.3 0.00115442 3.3 0.00115452 0 0.0011544399999999998 0 0.00115454 3.3 0.00115446 3.3 0.00115456 0 0.0011544799999999998 0 0.0011545799999999999 3.3 0.0011545 3.3 0.0011546 0 0.00115452 0 0.00115462 3.3 0.00115454 3.3 0.00115464 0 0.00115456 0 0.00115466 3.3 0.0011545799999999999 3.3 0.00115468 0 0.0011546 0 0.0011547 3.3 0.0011546199999999999 3.3 0.00115472 0 0.00115464 0 0.00115474 3.3 0.0011546599999999998 3.3 0.00115476 0 0.00115468 0 0.00115478 3.3 0.0011546999999999998 3.3 0.0011547999999999999 0 0.00115472 0 0.00115482 3.3 0.00115474 3.3 0.00115484 0 0.00115476 0 0.00115486 3.3 0.00115478 3.3 0.00115488 0 0.0011547999999999999 0 0.0011549 3.3 0.00115482 3.3 0.00115492 0 0.0011548399999999999 0 0.00115494 3.3 0.00115486 3.3 0.00115496 0 0.0011548799999999998 0 0.00115498 3.3 0.0011549 3.3 0.001155 0 0.0011549199999999998 0 0.0011550199999999999 3.3 0.00115494 3.3 0.00115504 0 0.00115496 0 0.00115506 3.3 0.00115498 3.3 0.00115508 0 0.001155 0 0.0011551 3.3 0.0011550199999999999 3.3 0.00115512 0 0.00115504 0 0.00115514 3.3 0.0011550599999999999 3.3 0.00115516 0 0.00115508 0 0.00115518 3.3 0.0011550999999999998 3.3 0.0011551999999999999 0 0.00115512 0 0.00115522 3.3 0.0011551399999999998 3.3 0.0011552399999999999 0 0.00115516 0 0.00115526 3.3 0.00115518 3.3 0.00115528 0 0.0011551999999999999 0 0.0011553 3.3 0.00115522 3.3 0.00115532 0 0.0011552399999999999 0 0.00115534 3.3 0.00115526 3.3 0.00115536 0 0.0011552799999999998 0 0.00115538 3.3 0.0011553 3.3 0.0011554 0 0.0011553199999999998 0 0.0011554199999999999 3.3 0.00115534 3.3 0.00115544 0 0.00115536 0 0.00115546 3.3 0.00115538 3.3 0.00115548 0 0.0011554 0 0.0011555 3.3 0.0011554199999999999 3.3 0.00115552 0 0.00115544 0 0.00115554 3.3 0.0011554599999999999 3.3 0.00115556 0 0.00115548 0 0.00115558 3.3 0.0011554999999999998 3.3 0.0011556 0 0.00115552 0 0.00115562 3.3 0.0011555399999999998 3.3 0.0011556399999999999 0 0.00115556 0 0.00115566 3.3 0.00115558 3.3 0.00115568 0 0.0011556 0 0.0011557 3.3 0.00115562 3.3 0.00115572 0 0.0011556399999999999 0 0.00115574 3.3 0.00115566 3.3 0.00115576 0 0.0011556799999999999 0 0.00115578 3.3 0.0011557 3.3 0.0011558 0 0.0011557199999999998 0 0.00115582 3.3 0.00115574 3.3 0.00115584 0 0.0011557599999999998 0 0.0011558599999999999 3.3 0.00115578 3.3 0.00115588 0 0.0011558 0 0.0011559 3.3 0.00115582 3.3 0.00115592 0 0.00115584 0 0.00115594 3.3 0.0011558599999999999 3.3 0.00115596 0 0.00115588 0 0.00115598 3.3 0.0011558999999999999 3.3 0.001156 0 0.00115592 0 0.00115602 3.3 0.0011559399999999998 3.3 0.0011560399999999999 0 0.00115596 0 0.00115606 3.3 0.00115598 3.3 0.00115608 0 0.001156 0 0.0011561 3.3 0.00115602 3.3 0.00115612 0 0.0011560399999999999 0 0.00115614 3.3 0.00115606 3.3 0.00115616 0 0.0011560799999999999 0 0.00115618 3.3 0.0011561 3.3 0.0011562 0 0.0011561199999999998 0 0.00115622 3.3 0.00115614 3.3 0.00115624 0 0.0011561599999999998 0 0.0011562599999999999 3.3 0.00115618 3.3 0.00115628 0 0.0011562 0 0.0011563 3.3 0.00115622 3.3 0.00115632 0 0.00115624 0 0.00115634 3.3 0.0011562599999999999 3.3 0.00115636 0 0.00115628 0 0.00115638 3.3 0.0011562999999999999 3.3 0.0011564 0 0.00115632 0 0.00115642 3.3 0.0011563399999999998 3.3 0.00115644 0 0.00115636 0 0.00115646 3.3 0.0011563799999999998 3.3 0.0011564799999999999 0 0.0011564 0 0.0011565 3.3 0.00115642 3.3 0.00115652 0 0.00115644 0 0.00115654 3.3 0.00115646 3.3 0.00115656 0 0.0011564799999999999 0 0.00115658 3.3 0.0011565 3.3 0.0011566 0 0.0011565199999999999 0 0.00115662 3.3 0.00115654 3.3 0.00115664 0 0.0011565599999999998 0 0.00115666 3.3 0.00115658 3.3 0.00115668 0 0.0011565999999999998 0 0.0011566999999999999 3.3 0.00115662 3.3 0.00115672 0 0.00115664 0 0.00115674 3.3 0.00115666 3.3 0.00115676 0 0.00115668 0 0.00115678 3.3 0.0011566999999999999 3.3 0.0011568 0 0.00115672 0 0.00115682 3.3 0.0011567399999999999 3.3 0.00115684 0 0.00115676 0 0.00115686 3.3 0.0011567799999999998 3.3 0.0011568799999999999 0 0.0011568 0 0.0011569 3.3 0.00115682 3.3 0.00115692 0 0.00115684 0 0.00115694 3.3 0.00115686 3.3 0.00115696 0 0.0011568799999999999 0 0.00115698 3.3 0.0011569 3.3 0.001157 0 0.0011569199999999999 0 0.00115702 3.3 0.00115694 3.3 0.00115704 0 0.0011569599999999998 0 0.00115706 3.3 0.00115698 3.3 0.00115708 0 0.0011569999999999998 0 0.0011570999999999999 3.3 0.00115702 3.3 0.00115712 0 0.00115704 0 0.00115714 3.3 0.00115706 3.3 0.00115716 0 0.00115708 0 0.00115718 3.3 0.0011570999999999999 3.3 0.0011572 0 0.00115712 0 0.00115722 3.3 0.0011571399999999999 3.3 0.00115724 0 0.00115716 0 0.00115726 3.3 0.0011571799999999998 3.3 0.00115728 0 0.0011572 0 0.0011573 3.3 0.0011572199999999998 3.3 0.0011573199999999999 0 0.00115724 0 0.00115734 3.3 0.00115726 3.3 0.00115736 0 0.00115728 0 0.00115738 3.3 0.0011573 3.3 0.0011574 0 0.0011573199999999999 0 0.00115742 3.3 0.00115734 3.3 0.00115744 0 0.0011573599999999999 0 0.00115746 3.3 0.00115738 3.3 0.00115748 0 0.0011573999999999998 0 0.0011575 3.3 0.00115742 3.3 0.00115752 0 0.0011574399999999998 0 0.0011575399999999999 3.3 0.00115746 3.3 0.00115756 0 0.00115748 0 0.00115758 3.3 0.0011575 3.3 0.0011576 0 0.00115752 0 0.00115762 3.3 0.0011575399999999999 3.3 0.00115764 0 0.00115756 0 0.00115766 3.3 0.0011575799999999999 3.3 0.00115768 0 0.0011576 0 0.0011577 3.3 0.0011576199999999998 3.3 0.0011577199999999999 0 0.00115764 0 0.00115774 3.3 0.00115766 3.3 0.00115776 0 0.00115768 0 0.00115778 3.3 0.0011577 3.3 0.0011578 0 0.0011577199999999999 0 0.00115782 3.3 0.00115774 3.3 0.00115784 0 0.0011577599999999999 0 0.00115786 3.3 0.00115778 3.3 0.00115788 0 0.0011577999999999998 0 0.0011579 3.3 0.00115782 3.3 0.00115792 0 0.0011578399999999998 0 0.0011579399999999999 3.3 0.00115786 3.3 0.00115796 0 0.00115788 0 0.00115798 3.3 0.0011579 3.3 0.001158 0 0.00115792 0 0.00115802 3.3 0.0011579399999999999 3.3 0.00115804 0 0.00115796 0 0.00115806 3.3 0.0011579799999999999 3.3 0.00115808 0 0.001158 0 0.0011581 3.3 0.0011580199999999998 3.3 0.00115812 0 0.00115804 0 0.00115814 3.3 0.0011580599999999998 3.3 0.0011581599999999999 0 0.00115808 0 0.00115818 3.3 0.0011581 3.3 0.0011582 0 0.00115812 0 0.00115822 3.3 0.00115814 3.3 0.00115824 0 0.0011581599999999999 0 0.00115826 3.3 0.00115818 3.3 0.00115828 0 0.0011581999999999999 0 0.0011583 3.3 0.00115822 3.3 0.00115832 0 0.0011582399999999998 0 0.0011583399999999999 3.3 0.00115826 3.3 0.00115836 0 0.0011582799999999998 0 0.0011583799999999999 3.3 0.0011583 3.3 0.0011584 0 0.00115832 0 0.00115842 3.3 0.0011583399999999999 3.3 0.00115844 0 0.00115836 0 0.00115846 3.3 0.0011583799999999999 3.3 0.00115848 0 0.0011584 0 0.0011585 3.3 0.0011584199999999998 3.3 0.00115852 0 0.00115844 0 0.00115854 3.3 0.0011584599999999998 3.3 0.0011585599999999999 0 0.00115848 0 0.00115858 3.3 0.0011585 3.3 0.0011586 0 0.00115852 0 0.00115862 3.3 0.00115854 3.3 0.00115864 0 0.0011585599999999999 0 0.00115866 3.3 0.00115858 3.3 0.00115868 0 0.0011585999999999999 0 0.0011587 3.3 0.00115862 3.3 0.00115872 0 0.0011586399999999998 0 0.00115874 3.3 0.00115866 3.3 0.00115876 0 0.0011586799999999998 0 0.0011587799999999999 3.3 0.0011587 3.3 0.0011588 0 0.00115872 0 0.00115882 3.3 0.00115874 3.3 0.00115884 0 0.00115876 0 0.00115886 3.3 0.0011587799999999999 3.3 0.00115888 0 0.0011588 0 0.0011589 3.3 0.0011588199999999999 3.3 0.00115892 0 0.00115884 0 0.00115894 3.3 0.0011588599999999998 3.3 0.00115896 0 0.00115888 0 0.00115898 3.3 0.0011588999999999998 3.3 0.0011589999999999999 0 0.00115892 0 0.00115902 3.3 0.00115894 3.3 0.00115904 0 0.00115896 0 0.00115906 3.3 0.00115898 3.3 0.00115908 0 0.0011589999999999999 0 0.0011591 3.3 0.00115902 3.3 0.00115912 0 0.0011590399999999999 0 0.00115914 3.3 0.00115906 3.3 0.00115916 0 0.0011590799999999998 0 0.0011591799999999999 3.3 0.0011591 3.3 0.0011592 0 0.0011591199999999998 0 0.0011592199999999999 3.3 0.00115914 3.3 0.00115924 0 0.00115916 0 0.00115926 3.3 0.0011591799999999999 3.3 0.00115928 0 0.0011592 0 0.0011593 3.3 0.0011592199999999999 3.3 0.00115932 0 0.00115924 0 0.00115934 3.3 0.0011592599999999998 3.3 0.00115936 0 0.00115928 0 0.00115938 3.3 0.0011592999999999998 3.3 0.0011593999999999999 0 0.00115932 0 0.00115942 3.3 0.00115934 3.3 0.00115944 0 0.00115936 0 0.00115946 3.3 0.00115938 3.3 0.00115948 0 0.0011593999999999999 0 0.0011595 3.3 0.00115942 3.3 0.00115952 0 0.0011594399999999999 0 0.00115954 3.3 0.00115946 3.3 0.00115956 0 0.0011594799999999998 0 0.00115958 3.3 0.0011595 3.3 0.0011596 0 0.0011595199999999998 0 0.0011596199999999999 3.3 0.00115954 3.3 0.00115964 0 0.00115956 0 0.00115966 3.3 0.00115958 3.3 0.00115968 0 0.0011596 0 0.0011597 3.3 0.0011596199999999999 3.3 0.00115972 0 0.00115964 0 0.00115974 3.3 0.0011596599999999999 3.3 0.00115976 0 0.00115968 0 0.00115978 3.3 0.0011596999999999998 3.3 0.0011598 0 0.00115972 0 0.00115982 3.3 0.0011597399999999998 3.3 0.0011598399999999999 0 0.00115976 0 0.00115986 3.3 0.00115978 3.3 0.00115988 0 0.0011598 0 0.0011599 3.3 0.00115982 3.3 0.00115992 0 0.0011598399999999999 0 0.00115994 3.3 0.00115986 3.3 0.00115996 0 0.0011598799999999999 0 0.00115998 3.3 0.0011599 3.3 0.00116 0 0.0011599199999999998 0 0.0011600199999999999 3.3 0.00115994 3.3 0.00116004 0 0.00115996 0 0.00116006 3.3 0.00115998 3.3 0.00116008 0 0.00116 0 0.0011601 3.3 0.0011600199999999999 3.3 0.00116012 0 0.00116004 0 0.00116014 3.3 0.0011600599999999999 3.3 0.00116016 0 0.00116008 0 0.00116018 3.3 0.0011600999999999998 3.3 0.0011602 0 0.00116012 0 0.00116022 3.3 0.0011601399999999998 3.3 0.0011602399999999999 0 0.00116016 0 0.00116026 3.3 0.00116018 3.3 0.00116028 0 0.0011602 0 0.0011603 3.3 0.00116022 3.3 0.00116032 0 0.0011602399999999999 0 0.00116034 3.3 0.00116026 3.3 0.00116036 0 0.0011602799999999999 0 0.00116038 3.3 0.0011603 3.3 0.0011604 0 0.0011603199999999998 0 0.00116042 3.3 0.00116034 3.3 0.00116044 0 0.0011603599999999998 0 0.0011604599999999999 3.3 0.00116038 3.3 0.00116048 0 0.0011604 0 0.0011605 3.3 0.00116042 3.3 0.00116052 0 0.00116044 0 0.00116054 3.3 0.0011604599999999999 3.3 0.00116056 0 0.00116048 0 0.00116058 3.3 0.0011604999999999999 3.3 0.0011606 0 0.00116052 0 0.00116062 3.3 0.0011605399999999998 3.3 0.00116064 0 0.00116056 0 0.00116066 3.3 0.0011605799999999998 3.3 0.0011606799999999999 0 0.0011606 0 0.0011607 3.3 0.00116062 3.3 0.00116072 0 0.00116064 0 0.00116074 3.3 0.00116066 3.3 0.00116076 0 0.0011606799999999999 0 0.00116078 3.3 0.0011607 3.3 0.0011608 0 0.0011607199999999999 0 0.00116082 3.3 0.00116074 3.3 0.00116084 0 0.0011607599999999998 0 0.0011608599999999999 3.3 0.00116078 3.3 0.00116088 0 0.0011608 0 0.0011609 3.3 0.00116082 3.3 0.00116092 0 0.00116084 0 0.00116094 3.3 0.0011608599999999999 3.3 0.00116096 0 0.00116088 0 0.00116098 3.3 0.0011608999999999999 3.3 0.001161 0 0.00116092 0 0.00116102 3.3 0.0011609399999999998 3.3 0.00116104 0 0.00116096 0 0.00116106 3.3 0.0011609799999999998 3.3 0.0011610799999999999 0 0.001161 0 0.0011611 3.3 0.00116102 3.3 0.00116112 0 0.00116104 0 0.00116114 3.3 0.00116106 3.3 0.00116116 0 0.0011610799999999999 0 0.00116118 3.3 0.0011611 3.3 0.0011612 0 0.0011611199999999999 0 0.00116122 3.3 0.00116114 3.3 0.00116124 0 0.0011611599999999998 0 0.00116126 3.3 0.00116118 3.3 0.00116128 0 0.0011611999999999998 0 0.0011612999999999999 3.3 0.00116122 3.3 0.00116132 0 0.00116124 0 0.00116134 3.3 0.00116126 3.3 0.00116136 0 0.00116128 0 0.00116138 3.3 0.0011612999999999999 3.3 0.0011614 0 0.00116132 0 0.00116142 3.3 0.0011613399999999999 3.3 0.00116144 0 0.00116136 0 0.00116146 3.3 0.0011613799999999998 3.3 0.0011614799999999999 0 0.0011614 0 0.0011615 3.3 0.0011614199999999998 3.3 0.0011615199999999999 0 0.00116144 0 0.00116154 3.3 0.00116146 3.3 0.00116156 0 0.0011614799999999999 0 0.00116158 3.3 0.0011615 3.3 0.0011616 0 0.0011615199999999999 0 0.00116162 3.3 0.00116154 3.3 0.00116164 0 0.0011615599999999998 0 0.00116166 3.3 0.00116158 3.3 0.00116168 0 0.0011615999999999998 0 0.0011616999999999999 3.3 0.00116162 3.3 0.00116172 0 0.00116164 0 0.00116174 3.3 0.00116166 3.3 0.00116176 0 0.00116168 0 0.00116178 3.3 0.0011616999999999999 3.3 0.0011618 0 0.00116172 0 0.00116182 3.3 0.0011617399999999999 3.3 0.00116184 0 0.00116176 0 0.00116186 3.3 0.0011617799999999998 3.3 0.00116188 0 0.0011618 0 0.0011619 3.3 0.0011618199999999998 3.3 0.0011619199999999999 0 0.00116184 0 0.00116194 3.3 0.00116186 3.3 0.00116196 0 0.00116188 0 0.00116198 3.3 0.0011619 3.3 0.001162 0 0.0011619199999999999 0 0.00116202 3.3 0.00116194 3.3 0.00116204 0 0.0011619599999999999 0 0.00116206 3.3 0.00116198 3.3 0.00116208 0 0.0011619999999999998 0 0.0011621 3.3 0.00116202 3.3 0.00116212 0 0.0011620399999999998 0 0.0011621399999999999 3.3 0.00116206 3.3 0.00116216 0 0.00116208 0 0.00116218 3.3 0.0011621 3.3 0.0011622 0 0.00116212 0 0.00116222 3.3 0.0011621399999999999 3.3 0.00116224 0 0.00116216 0 0.00116226 3.3 0.0011621799999999999 3.3 0.00116228 0 0.0011622 0 0.0011623 3.3 0.0011622199999999998 3.3 0.0011623199999999999 0 0.00116224 0 0.00116234 3.3 0.0011622599999999998 3.3 0.0011623599999999999 0 0.00116228 0 0.00116238 3.3 0.0011623 3.3 0.0011624 0 0.0011623199999999999 0 0.00116242 3.3 0.00116234 3.3 0.00116244 0 0.0011623599999999999 0 0.00116246 3.3 0.00116238 3.3 0.00116248 0 0.0011623999999999998 0 0.0011625 3.3 0.00116242 3.3 0.00116252 0 0.0011624399999999998 0 0.0011625399999999999 3.3 0.00116246 3.3 0.00116256 0 0.00116248 0 0.00116258 3.3 0.0011625 3.3 0.0011626 0 0.00116252 0 0.00116262 3.3 0.0011625399999999999 3.3 0.00116264 0 0.00116256 0 0.00116266 3.3 0.0011625799999999999 3.3 0.00116268 0 0.0011626 0 0.0011627 3.3 0.0011626199999999998 3.3 0.00116272 0 0.00116264 0 0.00116274 3.3 0.0011626599999999998 3.3 0.0011627599999999999 0 0.00116268 0 0.00116278 3.3 0.0011627 3.3 0.0011628 0 0.00116272 0 0.00116282 3.3 0.00116274 3.3 0.00116284 0 0.0011627599999999999 0 0.00116286 3.3 0.00116278 3.3 0.00116288 0 0.0011627999999999999 0 0.0011629 3.3 0.00116282 3.3 0.00116292 0 0.0011628399999999998 0 0.00116294 3.3 0.00116286 3.3 0.00116296 0 0.0011628799999999998 0 0.0011629799999999999 3.3 0.0011629 3.3 0.001163 0 0.00116292 0 0.00116302 3.3 0.00116294 3.3 0.00116304 0 0.00116296 0 0.00116306 3.3 0.0011629799999999999 3.3 0.00116308 0 0.001163 0 0.0011631 3.3 0.0011630199999999999 3.3 0.00116312 0 0.00116304 0 0.00116314 3.3 0.0011630599999999998 3.3 0.0011631599999999999 0 0.00116308 0 0.00116318 3.3 0.0011631 3.3 0.0011632 0 0.00116312 0 0.00116322 3.3 0.00116314 3.3 0.00116324 0 0.0011631599999999999 0 0.00116326 3.3 0.00116318 3.3 0.00116328 0 0.0011631999999999999 0 0.0011633 3.3 0.00116322 3.3 0.00116332 0 0.0011632399999999998 0 0.00116334 3.3 0.00116326 3.3 0.00116336 0 0.0011632799999999998 0 0.0011633799999999999 3.3 0.0011633 3.3 0.0011634 0 0.00116332 0 0.00116342 3.3 0.00116334 3.3 0.00116344 0 0.00116336 0 0.00116346 3.3 0.0011633799999999999 3.3 0.00116348 0 0.0011634 0 0.0011635 3.3 0.0011634199999999999 3.3 0.00116352 0 0.00116344 0 0.00116354 3.3 0.0011634599999999998 3.3 0.00116356 0 0.00116348 0 0.00116358 3.3 0.0011634999999999998 3.3 0.0011635999999999999 0 0.00116352 0 0.00116362 3.3 0.00116354 3.3 0.00116364 0 0.00116356 0 0.00116366 3.3 0.00116358 3.3 0.00116368 0 0.0011635999999999999 0 0.0011637 3.3 0.00116362 3.3 0.00116372 0 0.0011636399999999999 0 0.00116374 3.3 0.00116366 3.3 0.00116376 0 0.0011636799999999998 0 0.00116378 3.3 0.0011637 3.3 0.0011638 0 0.0011637199999999998 0 0.0011638199999999999 3.3 0.00116374 3.3 0.00116384 0 0.00116376 0 0.00116386 3.3 0.00116378 3.3 0.00116388 0 0.0011638 0 0.0011639 3.3 0.0011638199999999999 3.3 0.00116392 0 0.00116384 0 0.00116394 3.3 0.0011638599999999999 3.3 0.00116396 0 0.00116388 0 0.00116398 3.3 0.0011638999999999998 3.3 0.0011639999999999999 0 0.00116392 0 0.00116402 3.3 0.00116394 3.3 0.00116404 0 0.00116396 0 0.00116406 3.3 0.00116398 3.3 0.00116408 0 0.0011639999999999999 0 0.0011641 3.3 0.00116402 3.3 0.00116412 0 0.0011640399999999999 0 0.00116414 3.3 0.00116406 3.3 0.00116416 0 0.0011640799999999998 0 0.00116418 3.3 0.0011641 3.3 0.0011642 0 0.0011641199999999998 0 0.0011642199999999999 3.3 0.00116414 3.3 0.00116424 0 0.00116416 0 0.00116426 3.3 0.00116418 3.3 0.00116428 0 0.0011642 0 0.0011643 3.3 0.0011642199999999999 3.3 0.00116432 0 0.00116424 0 0.00116434 3.3 0.0011642599999999999 3.3 0.00116436 0 0.00116428 0 0.00116438 3.3 0.0011642999999999998 3.3 0.0011644 0 0.00116432 0 0.00116442 3.3 0.0011643399999999998 3.3 0.0011644399999999999 0 0.00116436 0 0.00116446 3.3 0.00116438 3.3 0.00116448 0 0.0011644 0 0.0011645 3.3 0.00116442 3.3 0.00116452 0 0.0011644399999999999 0 0.00116454 3.3 0.00116446 3.3 0.00116456 0 0.0011644799999999999 0 0.00116458 3.3 0.0011645 3.3 0.0011646 0 0.0011645199999999998 0 0.0011646199999999999 3.3 0.00116454 3.3 0.00116464 0 0.0011645599999999998 0 0.0011646599999999999 3.3 0.00116458 3.3 0.00116468 0 0.0011646 0 0.0011647 3.3 0.0011646199999999999 3.3 0.00116472 0 0.00116464 0 0.00116474 3.3 0.0011646599999999999 3.3 0.00116476 0 0.00116468 0 0.00116478 3.3 0.0011646999999999998 3.3 0.0011648 0 0.00116472 0 0.00116482 3.3 0.0011647399999999998 3.3 0.0011648399999999999 0 0.00116476 0 0.00116486 3.3 0.00116478 3.3 0.00116488 0 0.0011648 0 0.0011649 3.3 0.00116482 3.3 0.00116492 0 0.0011648399999999999 0 0.00116494 3.3 0.00116486 3.3 0.00116496 0 0.0011648799999999999 0 0.00116498 3.3 0.0011649 3.3 0.001165 0 0.0011649199999999998 0 0.00116502 3.3 0.00116494 3.3 0.00116504 0 0.0011649599999999998 0 0.0011650599999999999 3.3 0.00116498 3.3 0.00116508 0 0.001165 0 0.0011651 3.3 0.00116502 3.3 0.00116512 0 0.00116504 0 0.00116514 3.3 0.0011650599999999999 3.3 0.00116516 0 0.00116508 0 0.00116518 3.3 0.0011650999999999999 3.3 0.0011652 0 0.00116512 0 0.00116522 3.3 0.0011651399999999998 3.3 0.00116524 0 0.00116516 0 0.00116526 3.3 0.0011651799999999998 3.3 0.0011652799999999999 0 0.0011652 0 0.0011653 3.3 0.00116522 3.3 0.00116532 0 0.00116524 0 0.00116534 3.3 0.00116526 3.3 0.00116536 0 0.0011652799999999999 0 0.00116538 3.3 0.0011653 3.3 0.0011654 0 0.0011653199999999999 0 0.00116542 3.3 0.00116534 3.3 0.00116544 0 0.0011653599999999998 0 0.0011654599999999999 3.3 0.00116538 3.3 0.00116548 0 0.0011653999999999998 0 0.0011654999999999999 3.3 0.00116542 3.3 0.00116552 0 0.00116544 0 0.00116554 3.3 0.0011654599999999999 3.3 0.00116556 0 0.00116548 0 0.00116558 3.3 0.0011654999999999999 3.3 0.0011656 0 0.00116552 0 0.00116562 3.3 0.0011655399999999998 3.3 0.00116564 0 0.00116556 0 0.00116566 3.3 0.0011655799999999998 3.3 0.0011656799999999999 0 0.0011656 0 0.0011657 3.3 0.00116562 3.3 0.00116572 0 0.00116564 0 0.00116574 3.3 0.00116566 3.3 0.00116576 0 0.0011656799999999999 0 0.00116578 3.3 0.0011657 3.3 0.0011658 0 0.0011657199999999999 0 0.00116582 3.3 0.00116574 3.3 0.00116584 0 0.0011657599999999998 0 0.00116586 3.3 0.00116578 3.3 0.00116588 0 0.0011657999999999998 0 0.0011658999999999999 3.3 0.00116582 3.3 0.00116592 0 0.00116584 0 0.00116594 3.3 0.00116586 3.3 0.00116596 0 0.00116588 0 0.00116598 3.3 0.0011658999999999999 3.3 0.001166 0 0.00116592 0 0.00116602 3.3 0.0011659399999999999 3.3 0.00116604 0 0.00116596 0 0.00116606 3.3 0.0011659799999999998 3.3 0.00116608 0 0.001166 0 0.0011661 3.3 0.0011660199999999998 3.3 0.0011661199999999999 0 0.00116604 0 0.00116614 3.3 0.00116606 3.3 0.00116616 0 0.00116608 0 0.00116618 3.3 0.0011661 3.3 0.0011662 0 0.0011661199999999999 0 0.00116622 3.3 0.00116614 3.3 0.00116624 0 0.0011661599999999999 0 0.00116626 3.3 0.00116618 3.3 0.00116628 0 0.0011661999999999998 0 0.0011662999999999999 3.3 0.00116622 3.3 0.00116632 0 0.0011662399999999998 0 0.0011663399999999999 3.3 0.00116626 3.3 0.00116636 0 0.00116628 0 0.00116638 3.3 0.0011662999999999999 3.3 0.0011664 0 0.00116632 0 0.00116642 3.3 0.0011663399999999999 3.3 0.00116644 0 0.00116636 0 0.00116646 3.3 0.0011663799999999998 3.3 0.00116648 0 0.0011664 0 0.0011665 3.3 0.0011664199999999998 3.3 0.0011665199999999999 0 0.00116644 0 0.00116654 3.3 0.00116646 3.3 0.00116656 0 0.00116648 0 0.00116658 3.3 0.0011665 3.3 0.0011666 0 0.0011665199999999999 0 0.00116662 3.3 0.00116654 3.3 0.00116664 0 0.0011665599999999999 0 0.00116666 3.3 0.00116658 3.3 0.00116668 0 0.0011665999999999998 0 0.0011667 3.3 0.00116662 3.3 0.00116672 0 0.0011666399999999998 0 0.0011667399999999999 3.3 0.00116666 3.3 0.00116676 0 0.00116668 0 0.00116678 3.3 0.0011667 3.3 0.0011668 0 0.00116672 0 0.00116682 3.3 0.0011667399999999999 3.3 0.00116684 0 0.00116676 0 0.00116686 3.3 0.0011667799999999999 3.3 0.00116688 0 0.0011668 0 0.0011669 3.3 0.0011668199999999998 3.3 0.00116692 0 0.00116684 0 0.00116694 3.3 0.0011668599999999998 3.3 0.0011669599999999999 0 0.00116688 0 0.00116698 3.3 0.0011669 3.3 0.001167 0 0.00116692 0 0.00116702 3.3 0.00116694 3.3 0.00116704 0 0.0011669599999999999 0 0.00116706 3.3 0.00116698 3.3 0.00116708 0 0.0011669999999999999 0 0.0011671 3.3 0.00116702 3.3 0.00116712 0 0.0011670399999999998 0 0.0011671399999999999 3.3 0.00116706 3.3 0.00116716 0 0.00116708 0 0.00116718 3.3 0.0011671 3.3 0.0011672 0 0.00116712 0 0.00116722 3.3 0.0011671399999999999 3.3 0.00116724 0 0.00116716 0 0.00116726 3.3 0.0011671799999999999 3.3 0.00116728 0 0.0011672 0 0.0011673 3.3 0.0011672199999999998 3.3 0.00116732 0 0.00116724 0 0.00116734 3.3 0.0011672599999999998 3.3 0.0011673599999999999 0 0.00116728 0 0.00116738 3.3 0.0011673 3.3 0.0011674 0 0.00116732 0 0.00116742 3.3 0.00116734 3.3 0.00116744 0 0.0011673599999999999 0 0.00116746 3.3 0.00116738 3.3 0.00116748 0 0.0011673999999999999 0 0.0011675 3.3 0.00116742 3.3 0.00116752 0 0.0011674399999999998 0 0.00116754 3.3 0.00116746 3.3 0.00116756 0 0.0011674799999999998 0 0.0011675799999999999 3.3 0.0011675 3.3 0.0011676 0 0.00116752 0 0.00116762 3.3 0.00116754 3.3 0.00116764 0 0.00116756 0 0.00116766 3.3 0.0011675799999999999 3.3 0.00116768 0 0.0011676 0 0.0011677 3.3 0.0011676199999999999 3.3 0.00116772 0 0.00116764 0 0.00116774 3.3 0.0011676599999999998 3.3 0.00116776 0 0.00116768 0 0.00116778 3.3 0.0011676999999999998 3.3 0.0011677999999999999 0 0.00116772 0 0.00116782 3.3 0.00116774 3.3 0.00116784 0 0.00116776 0 0.00116786 3.3 0.00116778 3.3 0.00116788 0 0.0011677999999999999 0 0.0011679 3.3 0.00116782 3.3 0.00116792 0 0.0011678399999999999 0 0.00116794 3.3 0.00116786 3.3 0.00116796 0 0.0011678799999999998 0 0.0011679799999999999 3.3 0.0011679 3.3 0.001168 0 0.00116792 0 0.00116802 3.3 0.00116794 3.3 0.00116804 0 0.00116796 0 0.00116806 3.3 0.0011679799999999999 3.3 0.00116808 0 0.001168 0 0.0011681 3.3 0.0011680199999999999 3.3 0.00116812 0 0.00116804 0 0.00116814 3.3 0.0011680599999999998 3.3 0.00116816 0 0.00116808 0 0.00116818 3.3 0.0011680999999999998 3.3 0.0011681999999999999 0 0.00116812 0 0.00116822 3.3 0.00116814 3.3 0.00116824 0 0.00116816 0 0.00116826 3.3 0.00116818 3.3 0.00116828 0 0.0011681999999999999 0 0.0011683 3.3 0.00116822 3.3 0.00116832 0 0.0011682399999999999 0 0.00116834 3.3 0.00116826 3.3 0.00116836 0 0.0011682799999999998 0 0.00116838 3.3 0.0011683 3.3 0.0011684 0 0.0011683199999999998 0 0.0011684199999999999 3.3 0.00116834 3.3 0.00116844 0 0.00116836 0 0.00116846 3.3 0.00116838 3.3 0.00116848 0 0.0011684 0 0.0011685 3.3 0.0011684199999999999 3.3 0.00116852 0 0.00116844 0 0.00116854 3.3 0.0011684599999999999 3.3 0.00116856 0 0.00116848 0 0.00116858 3.3 0.0011684999999999998 3.3 0.0011685999999999999 0 0.00116852 0 0.00116862 3.3 0.0011685399999999998 3.3 0.0011686399999999999 0 0.00116856 0 0.00116866 3.3 0.00116858 3.3 0.00116868 0 0.0011685999999999999 0 0.0011687 3.3 0.00116862 3.3 0.00116872 0 0.0011686399999999999 0 0.00116874 3.3 0.00116866 3.3 0.00116876 0 0.0011686799999999998 0 0.00116878 3.3 0.0011687 3.3 0.0011688 0 0.0011687199999999998 0 0.0011688199999999999 3.3 0.00116874 3.3 0.00116884 0 0.00116876 0 0.00116886 3.3 0.00116878 3.3 0.00116888 0 0.0011688 0 0.0011689 3.3 0.0011688199999999999 3.3 0.00116892 0 0.00116884 0 0.00116894 3.3 0.0011688599999999999 3.3 0.00116896 0 0.00116888 0 0.00116898 3.3 0.0011688999999999998 3.3 0.001169 0 0.00116892 0 0.00116902 3.3 0.0011689399999999998 3.3 0.0011690399999999999 0 0.00116896 0 0.00116906 3.3 0.00116898 3.3 0.00116908 0 0.001169 0 0.0011691 3.3 0.00116902 3.3 0.00116912 0 0.0011690399999999999 0 0.00116914 3.3 0.00116906 3.3 0.00116916 0 0.0011690799999999999 0 0.00116918 3.3 0.0011691 3.3 0.0011692 0 0.0011691199999999998 0 0.00116922 3.3 0.00116914 3.3 0.00116924 0 0.0011691599999999998 0 0.0011692599999999999 3.3 0.00116918 3.3 0.00116928 0 0.0011692 0 0.0011693 3.3 0.00116922 3.3 0.00116932 0 0.00116924 0 0.00116934 3.3 0.0011692599999999999 3.3 0.00116936 0 0.00116928 0 0.00116938 3.3 0.0011692999999999999 3.3 0.0011694 0 0.00116932 0 0.00116942 3.3 0.0011693399999999998 3.3 0.0011694399999999999 0 0.00116936 0 0.00116946 3.3 0.0011693799999999998 3.3 0.0011694799999999999 0 0.0011694 0 0.0011695 3.3 0.00116942 3.3 0.00116952 0 0.0011694399999999999 0 0.00116954 3.3 0.00116946 3.3 0.00116956 0 0.0011694799999999999 0 0.00116958 3.3 0.0011695 3.3 0.0011696 0 0.0011695199999999998 0 0.00116962 3.3 0.00116954 3.3 0.00116964 0 0.0011695599999999998 0 0.0011696599999999999 3.3 0.00116958 3.3 0.00116968 0 0.0011696 0 0.0011697 3.3 0.00116962 3.3 0.00116972 0 0.00116964 0 0.00116974 3.3 0.0011696599999999999 3.3 0.00116976 0 0.00116968 0 0.00116978 3.3 0.0011696999999999999 3.3 0.0011698 0 0.00116972 0 0.00116982 3.3 0.0011697399999999998 3.3 0.00116984 0 0.00116976 0 0.00116986 3.3 0.0011697799999999998 3.3 0.0011698799999999999 0 0.0011698 0 0.0011699 3.3 0.00116982 3.3 0.00116992 0 0.00116984 0 0.00116994 3.3 0.00116986 3.3 0.00116996 0 0.0011698799999999999 0 0.00116998 3.3 0.0011699 3.3 0.00117 0 0.0011699199999999999 0 0.00117002 3.3 0.00116994 3.3 0.00117004 0 0.0011699599999999998 0 0.00117006 3.3 0.00116998 3.3 0.00117008 0 0.0011699999999999998 0 0.0011700999999999999 3.3 0.00117002 3.3 0.00117012 0 0.00117004 0 0.00117014 3.3 0.00117006 3.3 0.00117016 0 0.00117008 0 0.00117018 3.3 0.0011700999999999999 3.3 0.0011702 0 0.00117012 0 0.00117022 3.3 0.0011701399999999999 3.3 0.00117024 0 0.00117016 0 0.00117026 3.3 0.0011701799999999998 3.3 0.0011702799999999999 0 0.0011702 0 0.0011703 3.3 0.00117022 3.3 0.00117032 0 0.00117024 0 0.00117034 3.3 0.00117026 3.3 0.00117036 0 0.0011702799999999999 0 0.00117038 3.3 0.0011703 3.3 0.0011704 0 0.0011703199999999999 0 0.00117042 3.3 0.00117034 3.3 0.00117044 0 0.0011703599999999998 0 0.00117046 3.3 0.00117038 3.3 0.00117048 0 0.0011703999999999998 0 0.0011704999999999999 3.3 0.00117042 3.3 0.00117052 0 0.00117044 0 0.00117054 3.3 0.00117046 3.3 0.00117056 0 0.00117048 0 0.00117058 3.3 0.0011704999999999999 3.3 0.0011706 0 0.00117052 0 0.00117062 3.3 0.0011705399999999999 3.3 0.00117064 0 0.00117056 0 0.00117066 3.3 0.0011705799999999998 3.3 0.00117068 0 0.0011706 0 0.0011707 3.3 0.0011706199999999998 3.3 0.0011707199999999999 0 0.00117064 0 0.00117074 3.3 0.00117066 3.3 0.00117076 0 0.00117068 0 0.00117078 3.3 0.0011707 3.3 0.0011708 0 0.0011707199999999999 0 0.00117082 3.3 0.00117074 3.3 0.00117084 0 0.0011707599999999999 0 0.00117086 3.3 0.00117078 3.3 0.00117088 0 0.0011707999999999998 0 0.0011709 3.3 0.00117082 3.3 0.00117092 0 0.0011708399999999998 0 0.0011709399999999999 3.3 0.00117086 3.3 0.00117096 0 0.00117088 0 0.00117098 3.3 0.0011709 3.3 0.001171 0 0.00117092 0 0.00117102 3.3 0.0011709399999999999 3.3 0.00117104 0 0.00117096 0 0.00117106 3.3 0.0011709799999999999 3.3 0.00117108 0 0.001171 0 0.0011711 3.3 0.0011710199999999998 3.3 0.0011711199999999999 0 0.00117104 0 0.00117114 3.3 0.00117106 3.3 0.00117116 0 0.00117108 0 0.00117118 3.3 0.0011711 3.3 0.0011712 0 0.0011711199999999999 0 0.00117122 3.3 0.00117114 3.3 0.00117124 0 0.0011711599999999999 0 0.00117126 3.3 0.00117118 3.3 0.00117128 0 0.0011711999999999998 0 0.0011713 3.3 0.00117122 3.3 0.00117132 0 0.0011712399999999998 0 0.0011713399999999999 3.3 0.00117126 3.3 0.00117136 0 0.00117128 0 0.00117138 3.3 0.0011713 3.3 0.0011714 0 0.00117132 0 0.00117142 3.3 0.0011713399999999999 3.3 0.00117144 0 0.00117136 0 0.00117146 3.3 0.0011713799999999999 3.3 0.00117148 0 0.0011714 0 0.0011715 3.3 0.0011714199999999998 3.3 0.00117152 0 0.00117144 0 0.00117154 3.3 0.0011714599999999998 3.3 0.0011715599999999999 0 0.00117148 0 0.00117158 3.3 0.0011715 3.3 0.0011716 0 0.00117152 0 0.00117162 3.3 0.00117154 3.3 0.00117164 0 0.0011715599999999999 0 0.00117166 3.3 0.00117158 3.3 0.00117168 0 0.0011715999999999999 0 0.0011717 3.3 0.00117162 3.3 0.00117172 0 0.0011716399999999998 0 0.0011717399999999999 3.3 0.00117166 3.3 0.00117176 0 0.0011716799999999998 0 0.0011717799999999999 3.3 0.0011717 3.3 0.0011718 0 0.00117172 0 0.00117182 3.3 0.0011717399999999999 3.3 0.00117184 0 0.00117176 0 0.00117186 3.3 0.0011717799999999999 3.3 0.00117188 0 0.0011718 0 0.0011719 3.3 0.0011718199999999998 3.3 0.00117192 0 0.00117184 0 0.00117194 3.3 0.0011718599999999998 3.3 0.0011719599999999999 0 0.00117188 0 0.00117198 3.3 0.0011719 3.3 0.001172 0 0.00117192 0 0.00117202 3.3 0.00117194 3.3 0.00117204 0 0.0011719599999999999 0 0.00117206 3.3 0.00117198 3.3 0.00117208 0 0.0011719999999999999 0 0.0011721 3.3 0.00117202 3.3 0.00117212 0 0.0011720399999999998 0 0.00117214 3.3 0.00117206 3.3 0.00117216 0 0.0011720799999999998 0 0.0011721799999999999 3.3 0.0011721 3.3 0.0011722 0 0.00117212 0 0.00117222 3.3 0.00117214 3.3 0.00117224 0 0.00117216 0 0.00117226 3.3 0.0011721799999999999 3.3 0.00117228 0 0.0011722 0 0.0011723 3.3 0.0011722199999999999 3.3 0.00117232 0 0.00117224 0 0.00117234 3.3 0.0011722599999999998 3.3 0.00117236 0 0.00117228 0 0.00117238 3.3 0.0011722999999999998 3.3 0.0011723999999999999 0 0.00117232 0 0.00117242 3.3 0.00117234 3.3 0.00117244 0 0.00117236 0 0.00117246 3.3 0.00117238 3.3 0.00117248 0 0.0011723999999999999 0 0.0011725 3.3 0.00117242 3.3 0.00117252 0 0.0011724399999999999 0 0.00117254 3.3 0.00117246 3.3 0.00117256 0 0.0011724799999999998 0 0.0011725799999999999 3.3 0.0011725 3.3 0.0011726 0 0.0011725199999999998 0 0.0011726199999999999 3.3 0.00117254 3.3 0.00117264 0 0.00117256 0 0.00117266 3.3 0.0011725799999999999 3.3 0.00117268 0 0.0011726 0 0.0011727 3.3 0.0011726199999999999 3.3 0.00117272 0 0.00117264 0 0.00117274 3.3 0.0011726599999999998 3.3 0.00117276 0 0.00117268 0 0.00117278 3.3 0.0011726999999999998 3.3 0.0011727999999999999 0 0.00117272 0 0.00117282 3.3 0.00117274 3.3 0.00117284 0 0.00117276 0 0.00117286 3.3 0.00117278 3.3 0.00117288 0 0.0011727999999999999 0 0.0011729 3.3 0.00117282 3.3 0.00117292 0 0.0011728399999999999 0 0.00117294 3.3 0.00117286 3.3 0.00117296 0 0.0011728799999999998 0 0.00117298 3.3 0.0011729 3.3 0.001173 0 0.0011729199999999998 0 0.0011730199999999999 3.3 0.00117294 3.3 0.00117304 0 0.00117296 0 0.00117306 3.3 0.00117298 3.3 0.00117308 0 0.001173 0 0.0011731 3.3 0.0011730199999999999 3.3 0.00117312 0 0.00117304 0 0.00117314 3.3 0.0011730599999999999 3.3 0.00117316 0 0.00117308 0 0.00117318 3.3 0.0011730999999999998 3.3 0.0011732 0 0.00117312 0 0.00117322 3.3 0.0011731399999999998 3.3 0.0011732399999999999 0 0.00117316 0 0.00117326 3.3 0.00117318 3.3 0.00117328 0 0.0011732 0 0.0011733 3.3 0.00117322 3.3 0.00117332 0 0.0011732399999999999 0 0.00117334 3.3 0.00117326 3.3 0.00117336 0 0.0011732799999999999 0 0.00117338 3.3 0.0011733 3.3 0.0011734 0 0.0011733199999999998 0 0.0011734199999999999 3.3 0.00117334 3.3 0.00117344 0 0.00117336 0 0.00117346 3.3 0.00117338 3.3 0.00117348 0 0.0011734 0 0.0011735 3.3 0.0011734199999999999 3.3 0.00117352 0 0.00117344 0 0.00117354 3.3 0.0011734599999999999 3.3 0.00117356 0 0.00117348 0 0.00117358 3.3 0.0011734999999999998 3.3 0.0011736 0 0.00117352 0 0.00117362 3.3 0.0011735399999999998 3.3 0.0011736399999999999 0 0.00117356 0 0.00117366 3.3 0.00117358 3.3 0.00117368 0 0.0011736 0 0.0011737 3.3 0.00117362 3.3 0.00117372 0 0.0011736399999999999 0 0.00117374 3.3 0.00117366 3.3 0.00117376 0 0.0011736799999999999 0 0.00117378 3.3 0.0011737 3.3 0.0011738 0 0.0011737199999999998 0 0.00117382 3.3 0.00117374 3.3 0.00117384 0 0.0011737599999999998 0 0.0011738599999999999 3.3 0.00117378 3.3 0.00117388 0 0.0011738 0 0.0011739 3.3 0.00117382 3.3 0.00117392 0 0.00117384 0 0.00117394 3.3 0.0011738599999999999 3.3 0.00117396 0 0.00117388 0 0.00117398 3.3 0.0011738999999999999 3.3 0.001174 0 0.00117392 0 0.00117402 3.3 0.0011739399999999998 3.3 0.00117404 0 0.00117396 0 0.00117406 3.3 0.0011739799999999998 3.3 0.0011740799999999999 0 0.001174 0 0.0011741 3.3 0.00117402 3.3 0.00117412 0 0.00117404 0 0.00117414 3.3 0.00117406 3.3 0.00117416 0 0.0011740799999999999 0 0.00117418 3.3 0.0011741 3.3 0.0011742 0 0.0011741199999999999 0 0.00117422 3.3 0.00117414 3.3 0.00117424 0 0.0011741599999999998 0 0.0011742599999999999 3.3 0.00117418 3.3 0.00117428 0 0.0011742 0 0.0011743 3.3 0.00117422 3.3 0.00117432 0 0.00117424 0 0.00117434 3.3 0.0011742599999999999 3.3 0.00117436 0 0.00117428 0 0.00117438 3.3 0.0011742999999999999 3.3 0.0011744 0 0.00117432 0 0.00117442 3.3 0.0011743399999999998 3.3 0.00117444 0 0.00117436 0 0.00117446 3.3 0.0011743799999999998 3.3 0.0011744799999999999 0 0.0011744 0 0.0011745 3.3 0.00117442 3.3 0.00117452 0 0.00117444 0 0.00117454 3.3 0.00117446 3.3 0.00117456 0 0.0011744799999999999 0 0.00117458 3.3 0.0011745 3.3 0.0011746 0 0.0011745199999999999 0 0.00117462 3.3 0.00117454 3.3 0.00117464 0 0.0011745599999999998 0 0.00117466 3.3 0.00117458 3.3 0.00117468 0 0.0011745999999999998 0 0.0011746999999999999 3.3 0.00117462 3.3 0.00117472 0 0.00117464 0 0.00117474 3.3 0.00117466 3.3 0.00117476 0 0.00117468 0 0.00117478 3.3 0.0011746999999999999 3.3 0.0011748 0 0.00117472 0 0.00117482 3.3 0.0011747399999999999 3.3 0.00117484 0 0.00117476 0 0.00117486 3.3 0.0011747799999999998 3.3 0.0011748799999999999 0 0.0011748 0 0.0011749 3.3 0.0011748199999999998 3.3 0.0011749199999999999 0 0.00117484 0 0.00117494 3.3 0.00117486 3.3 0.00117496 0 0.0011748799999999999 0 0.00117498 3.3 0.0011749 3.3 0.001175 0 0.0011749199999999999 0 0.00117502 3.3 0.00117494 3.3 0.00117504 0 0.0011749599999999999 0 0.00117506 3.3 0.00117498 3.3 0.00117508 0 0.0011749999999999998 0 0.0011750999999999999 3.3 0.00117502 3.3 0.00117512 0 0.00117504 0 0.00117514 3.3 0.00117506 3.3 0.00117516 0 0.00117508 0 0.00117518 3.3 0.0011750999999999999 3.3 0.0011752 0 0.00117512 0 0.00117522 3.3 0.0011751399999999999 3.3 0.00117524 0 0.00117516 0 0.00117526 3.3 0.0011751799999999998 3.3 0.00117528 0 0.0011752 0 0.0011753 3.3 0.0011752199999999998 3.3 0.0011753199999999999 0 0.00117524 0 0.00117534 3.3 0.00117526 3.3 0.00117536 0 0.00117528 0 0.00117538 3.3 0.0011753 3.3 0.0011754 0 0.0011753199999999999 0 0.00117542 3.3 0.00117534 3.3 0.00117544 0 0.0011753599999999999 0 0.00117546 3.3 0.00117538 3.3 0.00117548 0 0.0011753999999999998 0 0.0011755 3.3 0.00117542 3.3 0.00117552 0 0.0011754399999999998 0 0.0011755399999999999 3.3 0.00117546 3.3 0.00117556 0 0.00117548 0 0.00117558 3.3 0.0011755 3.3 0.0011756 0 0.00117552 0 0.00117562 3.3 0.0011755399999999999 3.3 0.00117564 0 0.00117556 0 0.00117566 3.3 0.0011755799999999999 3.3 0.00117568 0 0.0011756 0 0.0011757 3.3 0.0011756199999999998 3.3 0.0011757199999999999 0 0.00117564 0 0.00117574 3.3 0.0011756599999999998 3.3 0.0011757599999999999 0 0.00117568 0 0.00117578 3.3 0.0011757 3.3 0.0011758 0 0.0011757199999999999 0 0.00117582 3.3 0.00117574 3.3 0.00117584 0 0.0011757599999999999 0 0.00117586 3.3 0.00117578 3.3 0.00117588 0 0.0011757999999999998 0 0.0011759 3.3 0.00117582 3.3 0.00117592 0 0.0011758399999999998 0 0.0011759399999999999 3.3 0.00117586 3.3 0.00117596 0 0.00117588 0 0.00117598 3.3 0.0011759 3.3 0.001176 0 0.00117592 0 0.00117602 3.3 0.0011759399999999999 3.3 0.00117604 0 0.00117596 0 0.00117606 3.3 0.0011759799999999999 3.3 0.00117608 0 0.001176 0 0.0011761 3.3 0.0011760199999999998 3.3 0.00117612 0 0.00117604 0 0.00117614 3.3 0.0011760599999999998 3.3 0.0011761599999999999 0 0.00117608 0 0.00117618 3.3 0.0011761 3.3 0.0011762 0 0.00117612 0 0.00117622 3.3 0.00117614 3.3 0.00117624 0 0.0011761599999999999 0 0.00117626 3.3 0.00117618 3.3 0.00117628 0 0.0011761999999999999 0 0.0011763 3.3 0.00117622 3.3 0.00117632 0 0.0011762399999999998 0 0.00117634 3.3 0.00117626 3.3 0.00117636 0 0.0011762799999999998 0 0.0011763799999999999 3.3 0.0011763 3.3 0.0011764 0 0.00117632 0 0.00117642 3.3 0.00117634 3.3 0.00117644 0 0.00117636 0 0.00117646 3.3 0.0011763799999999999 3.3 0.00117648 0 0.0011764 0 0.0011765 3.3 0.0011764199999999999 3.3 0.00117652 0 0.00117644 0 0.00117654 3.3 0.0011764599999999998 3.3 0.0011765599999999999 0 0.00117648 0 0.00117658 3.3 0.0011764999999999998 3.3 0.0011765999999999999 0 0.00117652 0 0.00117662 3.3 0.00117654 3.3 0.00117664 0 0.0011765599999999999 0 0.00117666 3.3 0.00117658 3.3 0.00117668 0 0.0011765999999999999 0 0.0011767 3.3 0.00117662 3.3 0.00117672 0 0.0011766399999999998 0 0.00117674 3.3 0.00117666 3.3 0.00117676 0 0.0011766799999999998 0 0.0011767799999999999 3.3 0.0011767 3.3 0.0011768 0 0.00117672 0 0.00117682 3.3 0.00117674 3.3 0.00117684 0 0.00117676 0 0.00117686 3.3 0.0011767799999999999 3.3 0.00117688 0 0.0011768 0 0.0011769 3.3 0.0011768199999999999 3.3 0.00117692 0 0.00117684 0 0.00117694 3.3 0.0011768599999999998 3.3 0.00117696 0 0.00117688 0 0.00117698 3.3 0.0011768999999999998 3.3 0.0011769999999999999 0 0.00117692 0 0.00117702 3.3 0.00117694 3.3 0.00117704 0 0.00117696 0 0.00117706 3.3 0.00117698 3.3 0.00117708 0 0.0011769999999999999 0 0.0011771 3.3 0.00117702 3.3 0.00117712 0 0.0011770399999999999 0 0.00117714 3.3 0.00117706 3.3 0.00117716 0 0.0011770799999999998 0 0.00117718 3.3 0.0011771 3.3 0.0011772 0 0.0011771199999999998 0 0.0011772199999999999 3.3 0.00117714 3.3 0.00117724 0 0.00117716 0 0.00117726 3.3 0.00117718 3.3 0.00117728 0 0.0011772 0 0.0011773 3.3 0.0011772199999999999 3.3 0.00117732 0 0.00117724 0 0.00117734 3.3 0.0011772599999999999 3.3 0.00117736 0 0.00117728 0 0.00117738 3.3 0.0011772999999999998 3.3 0.0011773999999999999 0 0.00117732 0 0.00117742 3.3 0.00117734 3.3 0.00117744 0 0.00117736 0 0.00117746 3.3 0.00117738 3.3 0.00117748 0 0.0011773999999999999 0 0.0011775 3.3 0.00117742 3.3 0.00117752 0 0.0011774399999999999 0 0.00117754 3.3 0.00117746 3.3 0.00117756 0 0.0011774799999999998 0 0.00117758 3.3 0.0011775 3.3 0.0011776 0 0.0011775199999999998 0 0.0011776199999999999 3.3 0.00117754 3.3 0.00117764 0 0.00117756 0 0.00117766 3.3 0.00117758 3.3 0.00117768 0 0.0011776 0 0.0011777 3.3 0.0011776199999999999 3.3 0.00117772 0 0.00117764 0 0.00117774 3.3 0.0011776599999999999 3.3 0.00117776 0 0.00117768 0 0.00117778 3.3 0.0011776999999999998 3.3 0.0011778 0 0.00117772 0 0.00117782 3.3 0.0011777399999999998 3.3 0.0011778399999999999 0 0.00117776 0 0.00117786 3.3 0.00117778 3.3 0.00117788 0 0.0011778 0 0.0011779 3.3 0.00117782 3.3 0.00117792 0 0.0011778399999999999 0 0.00117794 3.3 0.00117786 3.3 0.00117796 0 0.0011778799999999999 0 0.00117798 3.3 0.0011779 3.3 0.001178 0 0.0011779199999999998 0 0.00117802 3.3 0.00117794 3.3 0.00117804 0 0.0011779599999999998 0 0.0011780599999999999 3.3 0.00117798 3.3 0.00117808 0 0.001178 0 0.0011781 3.3 0.00117802 3.3 0.00117812 0 0.00117804 0 0.00117814 3.3 0.0011780599999999999 3.3 0.00117816 0 0.00117808 0 0.00117818 3.3 0.0011780999999999999 3.3 0.0011782 0 0.00117812 0 0.00117822 3.3 0.0011781399999999998 3.3 0.0011782399999999999 0 0.00117816 0 0.00117826 3.3 0.00117818 3.3 0.00117828 0 0.0011782 0 0.0011783 3.3 0.00117822 3.3 0.00117832 0 0.0011782399999999999 0 0.00117834 3.3 0.00117826 3.3 0.00117836 0 0.0011782799999999999 0 0.00117838 3.3 0.0011783 3.3 0.0011784 0 0.0011783199999999998 0 0.00117842 3.3 0.00117834 3.3 0.00117844 0 0.0011783599999999998 0 0.0011784599999999999 3.3 0.00117838 3.3 0.00117848 0 0.0011784 0 0.0011785 3.3 0.00117842 3.3 0.00117852 0 0.00117844 0 0.00117854 3.3 0.0011784599999999999 3.3 0.00117856 0 0.00117848 0 0.00117858 3.3 0.0011784999999999999 3.3 0.0011786 0 0.00117852 0 0.00117862 3.3 0.0011785399999999998 3.3 0.00117864 0 0.00117856 0 0.00117866 3.3 0.0011785799999999998 3.3 0.0011786799999999999 0 0.0011786 0 0.0011787 3.3 0.00117862 3.3 0.00117872 0 0.00117864 0 0.00117874 3.3 0.00117866 3.3 0.00117876 0 0.0011786799999999999 0 0.00117878 3.3 0.0011787 3.3 0.0011788 0 0.0011787199999999999 0 0.00117882 3.3 0.00117874 3.3 0.00117884 0 0.0011787599999999998 0 0.0011788599999999999 3.3 0.00117878 3.3 0.00117888 0 0.0011787999999999998 0 0.0011788999999999999 3.3 0.00117882 3.3 0.00117892 0 0.00117884 0 0.00117894 3.3 0.0011788599999999999 3.3 0.00117896 0 0.00117888 0 0.00117898 3.3 0.0011788999999999999 3.3 0.001179 0 0.00117892 0 0.00117902 3.3 0.0011789399999999998 3.3 0.00117904 0 0.00117896 0 0.00117906 3.3 0.0011789799999999998 3.3 0.0011790799999999999 0 0.001179 0 0.0011791 3.3 0.00117902 3.3 0.00117912 0 0.00117904 0 0.00117914 3.3 0.00117906 3.3 0.00117916 0 0.0011790799999999999 0 0.00117918 3.3 0.0011791 3.3 0.0011792 0 0.0011791199999999999 0 0.00117922 3.3 0.00117914 3.3 0.00117924 0 0.0011791599999999998 0 0.00117926 3.3 0.00117918 3.3 0.00117928 0 0.0011791999999999998 0 0.0011792999999999999 3.3 0.00117922 3.3 0.00117932 0 0.00117924 0 0.00117934 3.3 0.00117926 3.3 0.00117936 0 0.00117928 0 0.00117938 3.3 0.0011792999999999999 3.3 0.0011794 0 0.00117932 0 0.00117942 3.3 0.0011793399999999999 3.3 0.00117944 0 0.00117936 0 0.00117946 3.3 0.0011793799999999998 3.3 0.00117948 0 0.0011794 0 0.0011795 3.3 0.0011794199999999998 3.3 0.0011795199999999999 0 0.00117944 0 0.00117954 3.3 0.00117946 3.3 0.00117956 0 0.00117948 0 0.00117958 3.3 0.0011795 3.3 0.0011796 0 0.0011795199999999999 0 0.00117962 3.3 0.00117954 3.3 0.00117964 0 0.0011795599999999999 0 0.00117966 3.3 0.00117958 3.3 0.00117968 0 0.0011795999999999998 0 0.0011796999999999999 3.3 0.00117962 3.3 0.00117972 0 0.0011796399999999998 0 0.0011797399999999999 3.3 0.00117966 3.3 0.00117976 0 0.00117968 0 0.00117978 3.3 0.0011796999999999999 3.3 0.0011798 0 0.00117972 0 0.00117982 3.3 0.0011797399999999999 3.3 0.00117984 0 0.00117976 0 0.00117986 3.3 0.0011797799999999998 3.3 0.00117988 0 0.0011798 0 0.0011799 3.3 0.0011798199999999998 3.3 0.0011799199999999999 0 0.00117984 0 0.00117994 3.3 0.00117986 3.3 0.00117996 0 0.00117988 0 0.00117998 3.3 0.0011799 3.3 0.00118 0 0.0011799199999999999 0 0.00118002 3.3 0.00117994 3.3 0.00118004 0 0.0011799599999999999 0 0.00118006 3.3 0.00117998 3.3 0.00118008 0 0.0011799999999999998 0 0.0011801 3.3 0.00118002 3.3 0.00118012 0 0.0011800399999999998 0 0.0011801399999999999 3.3 0.00118006 3.3 0.00118016 0 0.00118008 0 0.00118018 3.3 0.0011801 3.3 0.0011802 0 0.00118012 0 0.00118022 3.3 0.0011801399999999999 3.3 0.00118024 0 0.00118016 0 0.00118026 3.3 0.0011801799999999999 3.3 0.00118028 0 0.0011802 0 0.0011803 3.3 0.0011802199999999998 3.3 0.00118032 0 0.00118024 0 0.00118034 3.3 0.0011802599999999998 3.3 0.0011803599999999999 0 0.00118028 0 0.00118038 3.3 0.0011803 3.3 0.0011804 0 0.00118032 0 0.00118042 3.3 0.00118034 3.3 0.00118044 0 0.0011803599999999999 0 0.00118046 3.3 0.00118038 3.3 0.00118048 0 0.0011803999999999999 0 0.0011805 3.3 0.00118042 3.3 0.00118052 0 0.0011804399999999998 0 0.0011805399999999999 3.3 0.00118046 3.3 0.00118056 0 0.00118048 0 0.00118058 3.3 0.0011805 3.3 0.0011806 0 0.00118052 0 0.00118062 3.3 0.0011805399999999999 3.3 0.00118064 0 0.00118056 0 0.00118066 3.3 0.0011805799999999999 3.3 0.00118068 0 0.0011806 0 0.0011807 3.3 0.0011806199999999998 3.3 0.00118072 0 0.00118064 0 0.00118074 3.3 0.0011806599999999998 3.3 0.0011807599999999999 0 0.00118068 0 0.00118078 3.3 0.0011807 3.3 0.0011808 0 0.00118072 0 0.00118082 3.3 0.00118074 3.3 0.00118084 0 0.0011807599999999999 0 0.00118086 3.3 0.00118078 3.3 0.00118088 0 0.0011807999999999999 0 0.0011809 3.3 0.00118082 3.3 0.00118092 0 0.0011808399999999998 0 0.00118094 3.3 0.00118086 3.3 0.00118096 0 0.0011808799999999998 0 0.0011809799999999999 3.3 0.0011809 3.3 0.001181 0 0.00118092 0 0.00118102 3.3 0.00118094 3.3 0.00118104 0 0.00118096 0 0.00118106 3.3 0.0011809799999999999 3.3 0.00118108 0 0.001181 0 0.0011811 3.3 0.0011810199999999999 3.3 0.00118112 0 0.00118104 0 0.00118114 3.3 0.0011810599999999998 3.3 0.00118116 0 0.00118108 0 0.00118118 3.3 0.0011810999999999998 3.3 0.0011811999999999999 0 0.00118112 0 0.00118122 3.3 0.00118114 3.3 0.00118124 0 0.00118116 0 0.00118126 3.3 0.00118118 3.3 0.00118128 0 0.0011811999999999999 0 0.0011813 3.3 0.00118122 3.3 0.00118132 0 0.0011812399999999999 0 0.00118134 3.3 0.00118126 3.3 0.00118136 0 0.0011812799999999998 0 0.0011813799999999999 3.3 0.0011813 3.3 0.0011814 0 0.00118132 0 0.00118142 3.3 0.00118134 3.3 0.00118144 0 0.00118136 0 0.00118146 3.3 0.0011813799999999999 3.3 0.00118148 0 0.0011814 0 0.0011815 3.3 0.0011814199999999999 3.3 0.00118152 0 0.00118144 0 0.00118154 3.3 0.0011814599999999998 3.3 0.00118156 0 0.00118148 0 0.00118158 3.3 0.0011814999999999998 3.3 0.0011815999999999999 0 0.00118152 0 0.00118162 3.3 0.00118154 3.3 0.00118164 0 0.00118156 0 0.00118166 3.3 0.00118158 3.3 0.00118168 0 0.0011815999999999999 0 0.0011817 3.3 0.00118162 3.3 0.00118172 0 0.0011816399999999999 0 0.00118174 3.3 0.00118166 3.3 0.00118176 0 0.0011816799999999998 0 0.00118178 3.3 0.0011817 3.3 0.0011818 0 0.0011817199999999998 0 0.0011818199999999999 3.3 0.00118174 3.3 0.00118184 0 0.00118176 0 0.00118186 3.3 0.00118178 3.3 0.00118188 0 0.0011818 0 0.0011819 3.3 0.0011818199999999999 3.3 0.00118192 0 0.00118184 0 0.00118194 3.3 0.0011818599999999999 3.3 0.00118196 0 0.00118188 0 0.00118198 3.3 0.0011818999999999998 3.3 0.0011819999999999999 0 0.00118192 0 0.00118202 3.3 0.0011819399999999998 3.3 0.0011820399999999999 0 0.00118196 0 0.00118206 3.3 0.00118198 3.3 0.00118208 0 0.0011819999999999999 0 0.0011821 3.3 0.00118202 3.3 0.00118212 0 0.0011820399999999999 0 0.00118214 3.3 0.00118206 3.3 0.00118216 0 0.0011820799999999998 0 0.00118218 3.3 0.0011821 3.3 0.0011822 0 0.0011821199999999998 0 0.0011822199999999999 3.3 0.00118214 3.3 0.00118224 0 0.00118216 0 0.00118226 3.3 0.00118218 3.3 0.00118228 0 0.0011822 0 0.0011823 3.3 0.0011822199999999999 3.3 0.00118232 0 0.00118224 0 0.00118234 3.3 0.0011822599999999999 3.3 0.00118236 0 0.00118228 0 0.00118238 3.3 0.0011822999999999998 3.3 0.0011824 0 0.00118232 0 0.00118242 3.3 0.0011823399999999998 3.3 0.0011824399999999999 0 0.00118236 0 0.00118246 3.3 0.00118238 3.3 0.00118248 0 0.0011824 0 0.0011825 3.3 0.00118242 3.3 0.00118252 0 0.0011824399999999999 0 0.00118254 3.3 0.00118246 3.3 0.00118256 0 0.0011824799999999999 0 0.00118258 3.3 0.0011825 3.3 0.0011826 0 0.0011825199999999998 0 0.00118262 3.3 0.00118254 3.3 0.00118264 0 0.0011825599999999998 0 0.0011826599999999999 3.3 0.00118258 3.3 0.00118268 0 0.0011826 0 0.0011827 3.3 0.00118262 3.3 0.00118272 0 0.00118264 0 0.00118274 3.3 0.0011826599999999999 3.3 0.00118276 0 0.00118268 0 0.00118278 3.3 0.0011826999999999999 3.3 0.0011828 0 0.00118272 0 0.00118282 3.3 0.0011827399999999998 3.3 0.0011828399999999999 0 0.00118276 0 0.00118286 3.3 0.0011827799999999998 3.3 0.0011828799999999999 0 0.0011828 0 0.0011829 3.3 0.00118282 3.3 0.00118292 0 0.0011828399999999999 0 0.00118294 3.3 0.00118286 3.3 0.00118296 0 0.0011828799999999999 0 0.00118298 3.3 0.0011829 3.3 0.001183 0 0.0011829199999999998 0 0.00118302 3.3 0.00118294 3.3 0.00118304 0 0.0011829599999999998 0 0.0011830599999999999 3.3 0.00118298 3.3 0.00118308 0 0.001183 0 0.0011831 3.3 0.00118302 3.3 0.00118312 0 0.00118304 0 0.00118314 3.3 0.0011830599999999999 3.3 0.00118316 0 0.00118308 0 0.00118318 3.3 0.0011830999999999999 3.3 0.0011832 0 0.00118312 0 0.00118322 3.3 0.0011831399999999998 3.3 0.00118324 0 0.00118316 0 0.00118326 3.3 0.0011831799999999998 3.3 0.0011832799999999999 0 0.0011832 0 0.0011833 3.3 0.00118322 3.3 0.00118332 0 0.00118324 0 0.00118334 3.3 0.00118326 3.3 0.00118336 0 0.0011832799999999999 0 0.00118338 3.3 0.0011833 3.3 0.0011834 0 0.0011833199999999999 0 0.00118342 3.3 0.00118334 3.3 0.00118344 0 0.0011833599999999998 0 0.00118346 3.3 0.00118338 3.3 0.00118348 0 0.0011833999999999998 0 0.0011834999999999999 3.3 0.00118342 3.3 0.00118352 0 0.00118344 0 0.00118354 3.3 0.00118346 3.3 0.00118356 0 0.00118348 0 0.00118358 3.3 0.0011834999999999999 3.3 0.0011836 0 0.00118352 0 0.00118362 3.3 0.0011835399999999999 3.3 0.00118364 0 0.00118356 0 0.00118366 3.3 0.0011835799999999998 3.3 0.0011836799999999999 0 0.0011836 0 0.0011837 3.3 0.0011836199999999998 3.3 0.0011837199999999999 0 0.00118364 0 0.00118374 3.3 0.00118366 3.3 0.00118376 0 0.0011836799999999999 0 0.00118378 3.3 0.0011837 3.3 0.0011838 0 0.0011837199999999999 0 0.00118382 3.3 0.00118374 3.3 0.00118384 0 0.0011837599999999998 0 0.00118386 3.3 0.00118378 3.3 0.00118388 0 0.0011837999999999998 0 0.0011838999999999999 3.3 0.00118382 3.3 0.00118392 0 0.00118384 0 0.00118394 3.3 0.00118386 3.3 0.00118396 0 0.00118388 0 0.00118398 3.3 0.0011838999999999999 3.3 0.001184 0 0.00118392 0 0.00118402 3.3 0.0011839399999999999 3.3 0.00118404 0 0.00118396 0 0.00118406 3.3 0.0011839799999999998 3.3 0.00118408 0 0.001184 0 0.0011841 3.3 0.0011840199999999998 3.3 0.0011841199999999999 0 0.00118404 0 0.00118414 3.3 0.00118406 3.3 0.00118416 0 0.00118408 0 0.00118418 3.3 0.0011841 3.3 0.0011842 0 0.0011841199999999999 0 0.00118422 3.3 0.00118414 3.3 0.00118424 0 0.0011841599999999999 0 0.00118426 3.3 0.00118418 3.3 0.00118428 0 0.0011841999999999998 0 0.0011843 3.3 0.00118422 3.3 0.00118432 0 0.0011842399999999998 0 0.0011843399999999999 3.3 0.00118426 3.3 0.00118436 0 0.00118428 0 0.00118438 3.3 0.0011843 3.3 0.0011844 0 0.00118432 0 0.00118442 3.3 0.0011843399999999999 3.3 0.00118444 0 0.00118436 0 0.00118446 3.3 0.0011843799999999999 3.3 0.00118448 0 0.0011844 0 0.0011845 3.3 0.0011844199999999998 3.3 0.0011845199999999999 0 0.00118444 0 0.00118454 3.3 0.00118446 3.3 0.00118456 0 0.00118448 0 0.00118458 3.3 0.0011845 3.3 0.0011846 0 0.0011845199999999999 0 0.00118462 3.3 0.00118454 3.3 0.00118464 0 0.0011845599999999999 0 0.00118466 3.3 0.00118458 3.3 0.00118468 0 0.0011845999999999998 0 0.0011847 3.3 0.00118462 3.3 0.00118472 0 0.0011846399999999998 0 0.0011847399999999999 3.3 0.00118466 3.3 0.00118476 0 0.00118468 0 0.00118478 3.3 0.0011847 3.3 0.0011848 0 0.00118472 0 0.00118482 3.3 0.0011847399999999999 3.3 0.00118484 0 0.00118476 0 0.00118486 3.3 0.0011847799999999999 3.3 0.00118488 0 0.0011848 0 0.0011849 3.3 0.0011848199999999998 3.3 0.00118492 0 0.00118484 0 0.00118494 3.3 0.0011848599999999998 3.3 0.0011849599999999999 0 0.00118488 0 0.00118498 3.3 0.0011849 3.3 0.001185 0 0.00118492 0 0.00118502 3.3 0.00118494 3.3 0.00118504 0 0.0011849599999999999 0 0.00118506 3.3 0.00118498 3.3 0.00118508 0 0.0011849999999999999 0 0.0011851 3.3 0.00118502 3.3 0.00118512 0 0.0011850399999999998 0 0.0011851399999999999 3.3 0.00118506 3.3 0.00118516 0 0.0011850799999999998 0 0.0011851799999999999 3.3 0.0011851 3.3 0.0011852 0 0.00118512 0 0.00118522 3.3 0.0011851399999999999 3.3 0.00118524 0 0.00118516 0 0.00118526 3.3 0.0011851799999999999 3.3 0.00118528 0 0.0011852 0 0.0011853 3.3 0.0011852199999999999 3.3 0.00118532 0 0.00118524 0 0.00118534 3.3 0.0011852599999999998 3.3 0.0011853599999999999 0 0.00118528 0 0.00118538 3.3 0.0011853 3.3 0.0011854 0 0.00118532 0 0.00118542 3.3 0.00118534 3.3 0.00118544 0 0.0011853599999999999 0 0.00118546 3.3 0.00118538 3.3 0.00118548 0 0.0011853999999999999 0 0.0011855 3.3 0.00118542 3.3 0.00118552 0 0.0011854399999999998 0 0.00118554 3.3 0.00118546 3.3 0.00118556 0 0.0011854799999999998 0 0.0011855799999999999 3.3 0.0011855 3.3 0.0011856 0 0.00118552 0 0.00118562 3.3 0.00118554 3.3 0.00118564 0 0.00118556 0 0.00118566 3.3 0.0011855799999999999 3.3 0.00118568 0 0.0011856 0 0.0011857 3.3 0.0011856199999999999 3.3 0.00118572 0 0.00118564 0 0.00118574 3.3 0.0011856599999999998 3.3 0.00118576 0 0.00118568 0 0.00118578 3.3 0.0011856999999999998 3.3 0.0011857999999999999 0 0.00118572 0 0.00118582 3.3 0.00118574 3.3 0.00118584 0 0.00118576 0 0.00118586 3.3 0.00118578 3.3 0.00118588 0 0.0011857999999999999 0 0.0011859 3.3 0.00118582 3.3 0.00118592 0 0.0011858399999999999 0 0.00118594 3.3 0.00118586 3.3 0.00118596 0 0.0011858799999999998 0 0.0011859799999999999 3.3 0.0011859 3.3 0.001186 0 0.0011859199999999998 0 0.0011860199999999999 3.3 0.00118594 3.3 0.00118604 0 0.00118596 0 0.00118606 3.3 0.0011859799999999999 3.3 0.00118608 0 0.001186 0 0.0011861 3.3 0.0011860199999999999 3.3 0.00118612 0 0.00118604 0 0.00118614 3.3 0.0011860599999999998 3.3 0.00118616 0 0.00118608 0 0.00118618 3.3 0.0011860999999999998 3.3 0.0011861999999999999 0 0.00118612 0 0.00118622 3.3 0.00118614 3.3 0.00118624 0 0.00118616 0 0.00118626 3.3 0.00118618 3.3 0.00118628 0 0.0011861999999999999 0 0.0011863 3.3 0.00118622 3.3 0.00118632 0 0.0011862399999999999 0 0.00118634 3.3 0.00118626 3.3 0.00118636 0 0.0011862799999999998 0 0.00118638 3.3 0.0011863 3.3 0.0011864 0 0.0011863199999999998 0 0.0011864199999999999 3.3 0.00118634 3.3 0.00118644 0 0.00118636 0 0.00118646 3.3 0.00118638 3.3 0.00118648 0 0.0011864 0 0.0011865 3.3 0.0011864199999999999 3.3 0.00118652 0 0.00118644 0 0.00118654 3.3 0.0011864599999999999 3.3 0.00118656 0 0.00118648 0 0.00118658 3.3 0.0011864999999999998 3.3 0.0011866 0 0.00118652 0 0.00118662 3.3 0.0011865399999999998 3.3 0.0011866399999999999 0 0.00118656 0 0.00118666 3.3 0.00118658 3.3 0.00118668 0 0.0011866 0 0.0011867 3.3 0.00118662 3.3 0.00118672 0 0.0011866399999999999 0 0.00118674 3.3 0.00118666 3.3 0.00118676 0 0.0011866799999999999 0 0.00118678 3.3 0.0011867 3.3 0.0011868 0 0.0011867199999999998 0 0.0011868199999999999 3.3 0.00118674 3.3 0.00118684 0 0.0011867599999999998 0 0.0011868599999999999 3.3 0.00118678 3.3 0.00118688 0 0.0011868 0 0.0011869 3.3 0.0011868199999999999 3.3 0.00118692 0 0.00118684 0 0.00118694 3.3 0.0011868599999999999 3.3 0.00118696 0 0.00118688 0 0.00118698 3.3 0.0011868999999999998 3.3 0.001187 0 0.00118692 0 0.00118702 3.3 0.0011869399999999998 3.3 0.0011870399999999999 0 0.00118696 0 0.00118706 3.3 0.00118698 3.3 0.00118708 0 0.001187 0 0.0011871 3.3 0.00118702 3.3 0.00118712 0 0.0011870399999999999 0 0.00118714 3.3 0.00118706 3.3 0.00118716 0 0.0011870799999999999 0 0.00118718 3.3 0.0011871 3.3 0.0011872 0 0.0011871199999999998 0 0.00118722 3.3 0.00118714 3.3 0.00118724 0 0.0011871599999999998 0 0.0011872599999999999 3.3 0.00118718 3.3 0.00118728 0 0.0011872 0 0.0011873 3.3 0.00118722 3.3 0.00118732 0 0.00118724 0 0.00118734 3.3 0.0011872599999999999 3.3 0.00118736 0 0.00118728 0 0.00118738 3.3 0.0011872999999999999 3.3 0.0011874 0 0.00118732 0 0.00118742 3.3 0.0011873399999999998 3.3 0.00118744 0 0.00118736 0 0.00118746 3.3 0.0011873799999999998 3.3 0.0011874799999999999 0 0.0011874 0 0.0011875 3.3 0.00118742 3.3 0.00118752 0 0.00118744 0 0.00118754 3.3 0.00118746 3.3 0.00118756 0 0.0011874799999999999 0 0.00118758 3.3 0.0011875 3.3 0.0011876 0 0.0011875199999999999 0 0.00118762 3.3 0.00118754 3.3 0.00118764 0 0.0011875599999999998 0 0.0011876599999999999 3.3 0.00118758 3.3 0.00118768 0 0.0011876 0 0.0011877 3.3 0.00118762 3.3 0.00118772 0 0.00118764 0 0.00118774 3.3 0.0011876599999999999 3.3 0.00118776 0 0.00118768 0 0.00118778 3.3 0.0011876999999999999 3.3 0.0011878 0 0.00118772 0 0.00118782 3.3 0.0011877399999999998 3.3 0.00118784 0 0.00118776 0 0.00118786 3.3 0.0011877799999999998 3.3 0.0011878799999999999 0 0.0011878 0 0.0011879 3.3 0.00118782 3.3 0.00118792 0 0.00118784 0 0.00118794 3.3 0.00118786 3.3 0.00118796 0 0.0011878799999999999 0 0.00118798 3.3 0.0011879 3.3 0.001188 0 0.0011879199999999999 0 0.00118802 3.3 0.00118794 3.3 0.00118804 0 0.0011879599999999998 0 0.00118806 3.3 0.00118798 3.3 0.00118808 0 0.0011879999999999998 0 0.0011880999999999999 3.3 0.00118802 3.3 0.00118812 0 0.00118804 0 0.00118814 3.3 0.00118806 3.3 0.00118816 0 0.00118808 0 0.00118818 3.3 0.0011880999999999999 3.3 0.0011882 0 0.00118812 0 0.00118822 3.3 0.0011881399999999999 3.3 0.00118824 0 0.00118816 0 0.00118826 3.3 0.0011881799999999998 3.3 0.00118828 0 0.0011882 0 0.0011883 3.3 0.0011882199999999998 3.3 0.0011883199999999999 0 0.00118824 0 0.00118834 3.3 0.00118826 3.3 0.00118836 0 0.00118828 0 0.00118838 3.3 0.0011883 3.3 0.0011884 0 0.0011883199999999999 0 0.00118842 3.3 0.00118834 3.3 0.00118844 0 0.0011883599999999999 0 0.00118846 3.3 0.00118838 3.3 0.00118848 0 0.0011883999999999998 0 0.0011884999999999999 3.3 0.00118842 3.3 0.00118852 0 0.00118844 0 0.00118854 3.3 0.00118846 3.3 0.00118856 0 0.00118848 0 0.00118858 3.3 0.0011884999999999999 3.3 0.0011886 0 0.00118852 0 0.00118862 3.3 0.0011885399999999999 3.3 0.00118864 0 0.00118856 0 0.00118866 3.3 0.0011885799999999998 3.3 0.00118868 0 0.0011886 0 0.0011887 3.3 0.0011886199999999998 3.3 0.0011887199999999999 0 0.00118864 0 0.00118874 3.3 0.00118866 3.3 0.00118876 0 0.00118868 0 0.00118878 3.3 0.0011887 3.3 0.0011888 0 0.0011887199999999999 0 0.00118882 3.3 0.00118874 3.3 0.00118884 0 0.0011887599999999999 0 0.00118886 3.3 0.00118878 3.3 0.00118888 0 0.0011887999999999998 0 0.0011889 3.3 0.00118882 3.3 0.00118892 0 0.0011888399999999998 0 0.0011889399999999999 3.3 0.00118886 3.3 0.00118896 0 0.00118888 0 0.00118898 3.3 0.0011889 3.3 0.001189 0 0.00118892 0 0.00118902 3.3 0.0011889399999999999 3.3 0.00118904 0 0.00118896 0 0.00118906 3.3 0.0011889799999999999 3.3 0.00118908 0 0.001189 0 0.0011891 3.3 0.0011890199999999998 3.3 0.0011891199999999999 0 0.00118904 0 0.00118914 3.3 0.0011890599999999998 3.3 0.0011891599999999999 0 0.00118908 0 0.00118918 3.3 0.0011891 3.3 0.0011892 0 0.0011891199999999999 0 0.00118922 3.3 0.00118914 3.3 0.00118924 0 0.0011891599999999999 0 0.00118926 3.3 0.00118918 3.3 0.00118928 0 0.0011891999999999998 0 0.0011893 3.3 0.00118922 3.3 0.00118932 0 0.0011892399999999998 0 0.0011893399999999999 3.3 0.00118926 3.3 0.00118936 0 0.00118928 0 0.00118938 3.3 0.0011893 3.3 0.0011894 0 0.00118932 0 0.00118942 3.3 0.0011893399999999999 3.3 0.00118944 0 0.00118936 0 0.00118946 3.3 0.0011893799999999999 3.3 0.00118948 0 0.0011894 0 0.0011895 3.3 0.0011894199999999998 3.3 0.00118952 0 0.00118944 0 0.00118954 3.3 0.0011894599999999998 3.3 0.0011895599999999999 0 0.00118948 0 0.00118958 3.3 0.0011895 3.3 0.0011896 0 0.00118952 0 0.00118962 3.3 0.00118954 3.3 0.00118964 0 0.0011895599999999999 0 0.00118966 3.3 0.00118958 3.3 0.00118968 0 0.0011895999999999999 0 0.0011897 3.3 0.00118962 3.3 0.00118972 0 0.0011896399999999998 0 0.00118974 3.3 0.00118966 3.3 0.00118976 0 0.0011896799999999998 0 0.0011897799999999999 3.3 0.0011897 3.3 0.0011898 0 0.00118972 0 0.00118982 3.3 0.00118974 3.3 0.00118984 0 0.00118976 0 0.00118986 3.3 0.0011897799999999999 3.3 0.00118988 0 0.0011898 0 0.0011899 3.3 0.0011898199999999999 3.3 0.00118992 0 0.00118984 0 0.00118994 3.3 0.0011898599999999998 3.3 0.0011899599999999999 0 0.00118988 0 0.00118998 3.3 0.0011898999999999998 3.3 0.0011899999999999999 0 0.00118992 0 0.00119002 3.3 0.00118994 3.3 0.00119004 0 0.0011899599999999999 0 0.00119006 3.3 0.00118998 3.3 0.00119008 0 0.0011899999999999999 0 0.0011901 3.3 0.00119002 3.3 0.00119012 0 0.0011900399999999998 0 0.00119014 3.3 0.00119006 3.3 0.00119016 0 0.0011900799999999998 0 0.0011901799999999999 3.3 0.0011901 3.3 0.0011902 0 0.00119012 0 0.00119022 3.3 0.00119014 3.3 0.00119024 0 0.00119016 0 0.00119026 3.3 0.0011901799999999999 3.3 0.00119028 0 0.0011902 0 0.0011903 3.3 0.0011902199999999999 3.3 0.00119032 0 0.00119024 0 0.00119034 3.3 0.0011902599999999998 3.3 0.00119036 0 0.00119028 0 0.00119038 3.3 0.0011902999999999998 3.3 0.0011903999999999999 0 0.00119032 0 0.00119042 3.3 0.00119034 3.3 0.00119044 0 0.00119036 0 0.00119046 3.3 0.00119038 3.3 0.00119048 0 0.0011903999999999999 0 0.0011905 3.3 0.00119042 3.3 0.00119052 0 0.0011904399999999999 0 0.00119054 3.3 0.00119046 3.3 0.00119056 0 0.0011904799999999998 0 0.00119058 3.3 0.0011905 3.3 0.0011906 0 0.0011905199999999998 0 0.0011906199999999999 3.3 0.00119054 3.3 0.00119064 0 0.00119056 0 0.00119066 3.3 0.00119058 3.3 0.00119068 0 0.0011906 0 0.0011907 3.3 0.0011906199999999999 3.3 0.00119072 0 0.00119064 0 0.00119074 3.3 0.0011906599999999999 3.3 0.00119076 0 0.00119068 0 0.00119078 3.3 0.0011906999999999998 3.3 0.0011907999999999999 0 0.00119072 0 0.00119082 3.3 0.00119074 3.3 0.00119084 0 0.00119076 0 0.00119086 3.3 0.00119078 3.3 0.00119088 0 0.0011907999999999999 0 0.0011909 3.3 0.00119082 3.3 0.00119092 0 0.0011908399999999999 0 0.00119094 3.3 0.00119086 3.3 0.00119096 0 0.0011908799999999998 0 0.00119098 3.3 0.0011909 3.3 0.001191 0 0.0011909199999999998 0 0.0011910199999999999 3.3 0.00119094 3.3 0.00119104 0 0.00119096 0 0.00119106 3.3 0.00119098 3.3 0.00119108 0 0.001191 0 0.0011911 3.3 0.0011910199999999999 3.3 0.00119112 0 0.00119104 0 0.00119114 3.3 0.0011910599999999999 3.3 0.00119116 0 0.00119108 0 0.00119118 3.3 0.0011910999999999998 3.3 0.0011912 0 0.00119112 0 0.00119122 3.3 0.0011911399999999998 3.3 0.0011912399999999999 0 0.00119116 0 0.00119126 3.3 0.00119118 3.3 0.00119128 0 0.0011912 0 0.0011913 3.3 0.00119122 3.3 0.00119132 0 0.0011912399999999999 0 0.00119134 3.3 0.00119126 3.3 0.00119136 0 0.0011912799999999999 0 0.00119138 3.3 0.0011913 3.3 0.0011914 0 0.0011913199999999998 0 0.00119142 3.3 0.00119134 3.3 0.00119144 0 0.0011913599999999998 0 0.0011914599999999999 3.3 0.00119138 3.3 0.00119148 0 0.0011914 0 0.0011915 3.3 0.00119142 3.3 0.00119152 0 0.00119144 0 0.00119154 3.3 0.0011914599999999999 3.3 0.00119156 0 0.00119148 0 0.00119158 3.3 0.0011914999999999999 3.3 0.0011916 0 0.00119152 0 0.00119162 3.3 0.0011915399999999998 3.3 0.0011916399999999999 0 0.00119156 0 0.00119166 3.3 0.00119158 3.3 0.00119168 0 0.0011916 0 0.0011917 3.3 0.00119162 3.3 0.00119172 0 0.0011916399999999999 0 0.00119174 3.3 0.00119166 3.3 0.00119176 0 0.0011916799999999999 0 0.00119178 3.3 0.0011917 3.3 0.0011918 0 0.0011917199999999998 0 0.00119182 3.3 0.00119174 3.3 0.00119184 0 0.0011917599999999998 0 0.0011918599999999999 3.3 0.00119178 3.3 0.00119188 0 0.0011918 0 0.0011919 3.3 0.00119182 3.3 0.00119192 0 0.00119184 0 0.00119194 3.3 0.0011918599999999999 3.3 0.00119196 0 0.00119188 0 0.00119198 3.3 0.0011918999999999999 3.3 0.001192 0 0.00119192 0 0.00119202 3.3 0.0011919399999999998 3.3 0.00119204 0 0.00119196 0 0.00119206 3.3 0.0011919799999999998 3.3 0.0011920799999999999 0 0.001192 0 0.0011921 3.3 0.00119202 3.3 0.00119212 0 0.00119204 0 0.00119214 3.3 0.00119206 3.3 0.00119216 0 0.0011920799999999999 0 0.00119218 3.3 0.0011921 3.3 0.0011922 0 0.0011921199999999999 0 0.00119222 3.3 0.00119214 3.3 0.00119224 0 0.0011921599999999998 0 0.0011922599999999999 3.3 0.00119218 3.3 0.00119228 0 0.0011921999999999998 0 0.0011922999999999999 3.3 0.00119222 3.3 0.00119232 0 0.00119224 0 0.00119234 3.3 0.0011922599999999999 3.3 0.00119236 0 0.00119228 0 0.00119238 3.3 0.0011922999999999999 3.3 0.0011924 0 0.00119232 0 0.00119242 3.3 0.0011923399999999998 3.3 0.00119244 0 0.00119236 0 0.00119246 3.3 0.0011923799999999998 3.3 0.0011924799999999999 0 0.0011924 0 0.0011925 3.3 0.00119242 3.3 0.00119252 0 0.00119244 0 0.00119254 3.3 0.00119246 3.3 0.00119256 0 0.0011924799999999999 0 0.00119258 3.3 0.0011925 3.3 0.0011926 0 0.0011925199999999999 0 0.00119262 3.3 0.00119254 3.3 0.00119264 0 0.0011925599999999998 0 0.00119266 3.3 0.00119258 3.3 0.00119268 0 0.0011925999999999998 0 0.0011926999999999999 3.3 0.00119262 3.3 0.00119272 0 0.00119264 0 0.00119274 3.3 0.00119266 3.3 0.00119276 0 0.00119268 0 0.00119278 3.3 0.0011926999999999999 3.3 0.0011928 0 0.00119272 0 0.00119282 3.3 0.0011927399999999999 3.3 0.00119284 0 0.00119276 0 0.00119286 3.3 0.0011927799999999998 3.3 0.00119288 0 0.0011928 0 0.0011929 3.3 0.0011928199999999998 3.3 0.0011929199999999999 0 0.00119284 0 0.00119294 3.3 0.00119286 3.3 0.00119296 0 0.00119288 0 0.00119298 3.3 0.0011929 3.3 0.001193 0 0.0011929199999999999 0 0.00119302 3.3 0.00119294 3.3 0.00119304 0 0.0011929599999999999 0 0.00119306 3.3 0.00119298 3.3 0.00119308 0 0.0011929999999999998 0 0.0011930999999999999 3.3 0.00119302 3.3 0.00119312 0 0.0011930399999999998 0 0.0011931399999999999 3.3 0.00119306 3.3 0.00119316 0 0.00119308 0 0.00119318 3.3 0.0011930999999999999 3.3 0.0011932 0 0.00119312 0 0.00119322 3.3 0.0011931399999999999 3.3 0.00119324 0 0.00119316 0 0.00119326 3.3 0.0011931799999999998 3.3 0.00119328 0 0.0011932 0 0.0011933 3.3 0.0011932199999999998 3.3 0.0011933199999999999 0 0.00119324 0 0.00119334 3.3 0.00119326 3.3 0.00119336 0 0.00119328 0 0.00119338 3.3 0.0011933 3.3 0.0011934 0 0.0011933199999999999 0 0.00119342 3.3 0.00119334 3.3 0.00119344 0 0.0011933599999999999 0 0.00119346 3.3 0.00119338 3.3 0.00119348 0 0.0011933999999999998 0 0.0011935 3.3 0.00119342 3.3 0.00119352 0 0.0011934399999999998 0 0.0011935399999999999 3.3 0.00119346 3.3 0.00119356 0 0.00119348 0 0.00119358 3.3 0.0011935 3.3 0.0011936 0 0.00119352 0 0.00119362 3.3 0.0011935399999999999 3.3 0.00119364 0 0.00119356 0 0.00119366 3.3 0.0011935799999999999 3.3 0.00119368 0 0.0011936 0 0.0011937 3.3 0.0011936199999999998 3.3 0.00119372 0 0.00119364 0 0.00119374 3.3 0.0011936599999999998 3.3 0.0011937599999999999 0 0.00119368 0 0.00119378 3.3 0.0011937 3.3 0.0011938 0 0.00119372 0 0.00119382 3.3 0.00119374 3.3 0.00119384 0 0.0011937599999999999 0 0.00119386 3.3 0.00119378 3.3 0.00119388 0 0.0011937999999999999 0 0.0011939 3.3 0.00119382 3.3 0.00119392 0 0.0011938399999999998 0 0.0011939399999999999 3.3 0.00119386 3.3 0.00119396 0 0.0011938799999999998 0 0.0011939799999999999 3.3 0.0011939 3.3 0.001194 0 0.00119392 0 0.00119402 3.3 0.0011939399999999999 3.3 0.00119404 0 0.00119396 0 0.00119406 3.3 0.0011939799999999999 3.3 0.00119408 0 0.001194 0 0.0011941 3.3 0.0011940199999999998 3.3 0.00119412 0 0.00119404 0 0.00119414 3.3 0.0011940599999999998 3.3 0.0011941599999999999 0 0.00119408 0 0.00119418 3.3 0.0011941 3.3 0.0011942 0 0.00119412 0 0.00119422 3.3 0.00119414 3.3 0.00119424 0 0.0011941599999999999 0 0.00119426 3.3 0.00119418 3.3 0.00119428 0 0.0011941999999999999 0 0.0011943 3.3 0.00119422 3.3 0.00119432 0 0.0011942399999999998 0 0.00119434 3.3 0.00119426 3.3 0.00119436 0 0.0011942799999999998 0 0.0011943799999999999 3.3 0.0011943 3.3 0.0011944 0 0.00119432 0 0.00119442 3.3 0.00119434 3.3 0.00119444 0 0.00119436 0 0.00119446 3.3 0.0011943799999999999 3.3 0.00119448 0 0.0011944 0 0.0011945 3.3 0.0011944199999999999 3.3 0.00119452 0 0.00119444 0 0.00119454 3.3 0.0011944599999999998 3.3 0.00119456 0 0.00119448 0 0.00119458 3.3 0.0011944999999999998 3.3 0.0011945999999999999 0 0.00119452 0 0.00119462 3.3 0.00119454 3.3 0.00119464 0 0.00119456 0 0.00119466 3.3 0.00119458 3.3 0.00119468 0 0.0011945999999999999 0 0.0011947 3.3 0.00119462 3.3 0.00119472 0 0.0011946399999999999 0 0.00119474 3.3 0.00119466 3.3 0.00119476 0 0.0011946799999999998 0 0.0011947799999999999 3.3 0.0011947 3.3 0.0011948 0 0.00119472 0 0.00119482 3.3 0.00119474 3.3 0.00119484 0 0.00119476 0 0.00119486 3.3 0.0011947799999999999 3.3 0.00119488 0 0.0011948 0 0.0011949 3.3 0.0011948199999999999 3.3 0.00119492 0 0.00119484 0 0.00119494 3.3 0.0011948599999999998 3.3 0.00119496 0 0.00119488 0 0.00119498 3.3 0.0011948999999999998 3.3 0.0011949999999999999 0 0.00119492 0 0.00119502 3.3 0.00119494 3.3 0.00119504 0 0.00119496 0 0.00119506 3.3 0.00119498 3.3 0.00119508 0 0.0011949999999999999 0 0.0011951 3.3 0.00119502 3.3 0.00119512 0 0.0011950399999999999 0 0.00119514 3.3 0.00119506 3.3 0.00119516 0 0.0011950799999999998 0 0.00119518 3.3 0.0011951 3.3 0.0011952 0 0.0011951199999999998 0 0.0011952199999999999 3.3 0.00119514 3.3 0.00119524 0 0.00119516 0 0.00119526 3.3 0.00119518 3.3 0.00119528 0 0.0011952 0 0.0011953 3.3 0.0011952199999999999 3.3 0.00119532 0 0.00119524 0 0.00119534 3.3 0.0011952599999999999 3.3 0.00119536 0 0.00119528 0 0.00119538 3.3 0.0011952999999999998 3.3 0.0011953999999999999 0 0.00119532 0 0.00119542 3.3 0.0011953399999999998 3.3 0.0011954399999999999 0 0.00119536 0 0.00119546 3.3 0.00119538 3.3 0.00119548 0 0.0011953999999999999 0 0.0011955 3.3 0.00119542 3.3 0.00119552 0 0.0011954399999999999 0 0.00119554 3.3 0.00119546 3.3 0.00119556 0 0.0011954799999999999 0 0.00119558 3.3 0.0011955 3.3 0.0011956 0 0.0011955199999999998 0 0.0011956199999999999 3.3 0.00119554 3.3 0.00119564 0 0.00119556 0 0.00119566 3.3 0.00119558 3.3 0.00119568 0 0.0011956 0 0.0011957 3.3 0.0011956199999999999 3.3 0.00119572 0 0.00119564 0 0.00119574 3.3 0.0011956599999999999 3.3 0.00119576 0 0.00119568 0 0.00119578 3.3 0.0011956999999999998 3.3 0.0011958 0 0.00119572 0 0.00119582 3.3 0.0011957399999999998 3.3 0.0011958399999999999 0 0.00119576 0 0.00119586 3.3 0.00119578 3.3 0.00119588 0 0.0011958 0 0.0011959 3.3 0.00119582 3.3 0.00119592 0 0.0011958399999999999 0 0.00119594 3.3 0.00119586 3.3 0.00119596 0 0.0011958799999999999 0 0.00119598 3.3 0.0011959 3.3 0.001196 0 0.0011959199999999998 0 0.00119602 3.3 0.00119594 3.3 0.00119604 0 0.0011959599999999998 0 0.0011960599999999999 3.3 0.00119598 3.3 0.00119608 0 0.001196 0 0.0011961 3.3 0.00119602 3.3 0.00119612 0 0.00119604 0 0.00119614 3.3 0.0011960599999999999 3.3 0.00119616 0 0.00119608 0 0.00119618 3.3 0.0011960999999999999 3.3 0.0011962 0 0.00119612 0 0.00119622 3.3 0.0011961399999999998 3.3 0.0011962399999999999 0 0.00119616 0 0.00119626 3.3 0.0011961799999999998 3.3 0.0011962799999999999 0 0.0011962 0 0.0011963 3.3 0.00119622 3.3 0.00119632 0 0.0011962399999999999 0 0.00119634 3.3 0.00119626 3.3 0.00119636 0 0.0011962799999999999 0 0.00119638 3.3 0.0011963 3.3 0.0011964 0 0.0011963199999999998 0 0.00119642 3.3 0.00119634 3.3 0.00119644 0 0.0011963599999999998 0 0.0011964599999999999 3.3 0.00119638 3.3 0.00119648 0 0.0011964 0 0.0011965 3.3 0.00119642 3.3 0.00119652 0 0.00119644 0 0.00119654 3.3 0.0011964599999999999 3.3 0.00119656 0 0.00119648 0 0.00119658 3.3 0.0011964999999999999 3.3 0.0011966 0 0.00119652 0 0.00119662 3.3 0.0011965399999999998 3.3 0.00119664 0 0.00119656 0 0.00119666 3.3 0.0011965799999999998 3.3 0.0011966799999999999 0 0.0011966 0 0.0011967 3.3 0.00119662 3.3 0.00119672 0 0.00119664 0 0.00119674 3.3 0.00119666 3.3 0.00119676 0 0.0011966799999999999 0 0.00119678 3.3 0.0011967 3.3 0.0011968 0 0.0011967199999999999 0 0.00119682 3.3 0.00119674 3.3 0.00119684 0 0.0011967599999999998 0 0.00119686 3.3 0.00119678 3.3 0.00119688 0 0.0011967999999999998 0 0.0011968999999999999 3.3 0.00119682 3.3 0.00119692 0 0.00119684 0 0.00119694 3.3 0.00119686 3.3 0.00119696 0 0.00119688 0 0.00119698 3.3 0.0011968999999999999 3.3 0.001197 0 0.00119692 0 0.00119702 3.3 0.0011969399999999999 3.3 0.00119704 0 0.00119696 0 0.00119706 3.3 0.0011969799999999998 3.3 0.0011970799999999999 0 0.001197 0 0.0011971 3.3 0.0011970199999999998 3.3 0.0011971199999999999 0 0.00119704 0 0.00119714 3.3 0.00119706 3.3 0.00119716 0 0.0011970799999999999 0 0.00119718 3.3 0.0011971 3.3 0.0011972 0 0.0011971199999999999 0 0.00119722 3.3 0.00119714 3.3 0.00119724 0 0.0011971599999999998 0 0.00119726 3.3 0.00119718 3.3 0.00119728 0 0.0011971999999999998 0 0.0011972999999999999 3.3 0.00119722 3.3 0.00119732 0 0.00119724 0 0.00119734 3.3 0.00119726 3.3 0.00119736 0 0.00119728 0 0.00119738 3.3 0.0011972999999999999 3.3 0.0011974 0 0.00119732 0 0.00119742 3.3 0.0011973399999999999 3.3 0.00119744 0 0.00119736 0 0.00119746 3.3 0.0011973799999999998 3.3 0.00119748 0 0.0011974 0 0.0011975 3.3 0.0011974199999999998 3.3 0.0011975199999999999 0 0.00119744 0 0.00119754 3.3 0.00119746 3.3 0.00119756 0 0.00119748 0 0.00119758 3.3 0.0011975 3.3 0.0011976 0 0.0011975199999999999 0 0.00119762 3.3 0.00119754 3.3 0.00119764 0 0.0011975599999999999 0 0.00119766 3.3 0.00119758 3.3 0.00119768 0 0.0011975999999999998 0 0.0011977 3.3 0.00119762 3.3 0.00119772 0 0.0011976399999999998 0 0.0011977399999999999 3.3 0.00119766 3.3 0.00119776 0 0.00119768 0 0.00119778 3.3 0.0011977 3.3 0.0011978 0 0.00119772 0 0.00119782 3.3 0.0011977399999999999 3.3 0.00119784 0 0.00119776 0 0.00119786 3.3 0.0011977799999999999 3.3 0.00119788 0 0.0011978 0 0.0011979 3.3 0.0011978199999999998 3.3 0.0011979199999999999 0 0.00119784 0 0.00119794 3.3 0.00119786 3.3 0.00119796 0 0.00119788 0 0.00119798 3.3 0.0011979 3.3 0.001198 0 0.0011979199999999999 0 0.00119802 3.3 0.00119794 3.3 0.00119804 0 0.0011979599999999999 0 0.00119806 3.3 0.00119798 3.3 0.00119808 0 0.0011979999999999998 0 0.0011981 3.3 0.00119802 3.3 0.00119812 0 0.0011980399999999998 0 0.0011981399999999999 3.3 0.00119806 3.3 0.00119816 0 0.00119808 0 0.00119818 3.3 0.0011981 3.3 0.0011982 0 0.00119812 0 0.00119822 3.3 0.0011981399999999999 3.3 0.00119824 0 0.00119816 0 0.00119826 3.3 0.0011981799999999999 3.3 0.00119828 0 0.0011982 0 0.0011983 3.3 0.0011982199999999998 3.3 0.00119832 0 0.00119824 0 0.00119834 3.3 0.0011982599999999998 3.3 0.0011983599999999999 0 0.00119828 0 0.00119838 3.3 0.0011983 3.3 0.0011984 0 0.00119832 0 0.00119842 3.3 0.00119834 3.3 0.00119844 0 0.0011983599999999999 0 0.00119846 3.3 0.00119838 3.3 0.00119848 0 0.0011983999999999999 0 0.0011985 3.3 0.00119842 3.3 0.00119852 0 0.0011984399999999998 0 0.00119854 3.3 0.00119846 3.3 0.00119856 0 0.0011984799999999998 0 0.0011985799999999999 3.3 0.0011985 3.3 0.0011986 0 0.00119852 0 0.00119862 3.3 0.00119854 3.3 0.00119864 0 0.00119856 0 0.00119866 3.3 0.0011985799999999999 3.3 0.00119868 0 0.0011986 0 0.0011987 3.3 0.0011986199999999999 3.3 0.00119872 0 0.00119864 0 0.00119874 3.3 0.0011986599999999998 3.3 0.0011987599999999999 0 0.00119868 0 0.00119878 3.3 0.0011987 3.3 0.0011988 0 0.00119872 0 0.00119882 3.3 0.00119874 3.3 0.00119884 0 0.0011987599999999999 0 0.00119886 3.3 0.00119878 3.3 0.00119888 0 0.0011987999999999999 0 0.0011989 3.3 0.00119882 3.3 0.00119892 0 0.0011988399999999998 0 0.00119894 3.3 0.00119886 3.3 0.00119896 0 0.0011988799999999998 0 0.0011989799999999999 3.3 0.0011989 3.3 0.001199 0 0.00119892 0 0.00119902 3.3 0.00119894 3.3 0.00119904 0 0.00119896 0 0.00119906 3.3 0.0011989799999999999 3.3 0.00119908 0 0.001199 0 0.0011991 3.3 0.0011990199999999999 3.3 0.00119912 0 0.00119904 0 0.00119914 3.3 0.0011990599999999998 3.3 0.00119916 0 0.00119908 0 0.00119918 3.3 0.0011990999999999998 3.3 0.0011991999999999999 0 0.00119912 0 0.00119922 3.3 0.00119914 3.3 0.00119924 0 0.00119916 0 0.00119926 3.3 0.00119918 3.3 0.00119928 0 0.0011991999999999999 0 0.0011993 3.3 0.00119922 3.3 0.00119932 0 0.0011992399999999999 0 0.00119934 3.3 0.00119926 3.3 0.00119936 0 0.0011992799999999998 0 0.0011993799999999999 3.3 0.0011993 3.3 0.0011994 0 0.0011993199999999998 0 0.0011994199999999999 3.3 0.00119934 3.3 0.00119944 0 0.00119936 0 0.00119946 3.3 0.0011993799999999999 3.3 0.00119948 0 0.0011994 0 0.0011995 3.3 0.0011994199999999999 3.3 0.00119952 0 0.00119944 0 0.00119954 3.3 0.0011994599999999998 3.3 0.00119956 0 0.00119948 0 0.00119958 3.3 0.0011994999999999998 3.3 0.0011995999999999999 0 0.00119952 0 0.00119962 3.3 0.00119954 3.3 0.00119964 0 0.00119956 0 0.00119966 3.3 0.00119958 3.3 0.00119968 0 0.0011995999999999999 0 0.0011997 3.3 0.00119962 3.3 0.00119972 0 0.0011996399999999999 0 0.00119974 3.3 0.00119966 3.3 0.00119976 0 0.0011996799999999998 0 0.00119978 3.3 0.0011997 3.3 0.0011998 0 0.0011997199999999998 0 0.0011998199999999999 3.3 0.00119974 3.3 0.00119984 0 0.00119976 0 0.00119986 3.3 0.00119978 3.3 0.00119988 0 0.0011998 0 0.0011999 3.3 0.0011998199999999999 3.3 0.00119992 0 0.00119984 0 0.00119994 3.3 0.0011998599999999999 3.3 0.00119996 0 0.00119988 0 0.00119998 3.3 0.0011998999999999998 3.3 0.0012 0 0.00119992 0 0.00120002 3.3 0.0011999399999999998 3.3 0.0012000399999999999 0 0.00119996 0 0.00120006 3.3 0.00119998 3.3 0.00120008 0 0.0012 0 0.0012001 3.3 0.00120002 3.3 0.00120012 0 0.0012000399999999999 0 0.00120014 3.3 0.00120006 3.3 0.00120016 0 0.0012000799999999999 0 0.00120018 3.3 0.0012001 3.3 0.0012002 0 0.0012001199999999998 0 0.0012002199999999999 3.3 0.00120014 3.3 0.00120024 0 0.0012001599999999998 0 0.0012002599999999999 3.3 0.00120018 3.3 0.00120028 0 0.0012002 0 0.0012003 3.3 0.0012002199999999999 3.3 0.00120032 0 0.00120024 0 0.00120034 3.3 0.0012002599999999999 3.3 0.00120036 0 0.00120028 0 0.00120038 3.3 0.0012002999999999998 3.3 0.0012004 0 0.00120032 0 0.00120042 3.3 0.0012003399999999998 3.3 0.0012004399999999999 0 0.00120036 0 0.00120046 3.3 0.00120038 3.3 0.00120048 0 0.0012004 0 0.0012005 3.3 0.00120042 3.3 0.00120052 0 0.0012004399999999999 0 0.00120054 3.3 0.00120046 3.3 0.00120056 0 0.0012004799999999999 0 0.00120058 3.3 0.0012005 3.3 0.0012006 0 0.0012005199999999998 0 0.00120062 3.3 0.00120054 3.3 0.00120064 0 0.0012005599999999998 0 0.0012006599999999999 3.3 0.00120058 3.3 0.00120068 0 0.0012006 0 0.0012007 3.3 0.00120062 3.3 0.00120072 0 0.00120064 0 0.00120074 3.3 0.0012006599999999999 3.3 0.00120076 0 0.00120068 0 0.00120078 3.3 0.0012006999999999999 3.3 0.0012008 0 0.00120072 0 0.00120082 3.3 0.0012007399999999998 3.3 0.00120084 0 0.00120076 0 0.00120086 3.3 0.0012007799999999998 3.3 0.0012008799999999999 0 0.0012008 0 0.0012009 3.3 0.00120082 3.3 0.00120092 0 0.00120084 0 0.00120094 3.3 0.00120086 3.3 0.00120096 0 0.0012008799999999999 0 0.00120098 3.3 0.0012009 3.3 0.001201 0 0.0012009199999999999 0 0.00120102 3.3 0.00120094 3.3 0.00120104 0 0.0012009599999999998 0 0.0012010599999999999 3.3 0.00120098 3.3 0.00120108 0 0.001201 0 0.0012011 3.3 0.00120102 3.3 0.00120112 0 0.00120104 0 0.00120114 3.3 0.0012010599999999999 3.3 0.00120116 0 0.00120108 0 0.00120118 3.3 0.0012010999999999999 3.3 0.0012012 0 0.00120112 0 0.00120122 3.3 0.0012011399999999998 3.3 0.00120124 0 0.00120116 0 0.00120126 3.3 0.0012011799999999998 3.3 0.0012012799999999999 0 0.0012012 0 0.0012013 3.3 0.00120122 3.3 0.00120132 0 0.00120124 0 0.00120134 3.3 0.00120126 3.3 0.00120136 0 0.0012012799999999999 0 0.00120138 3.3 0.0012013 3.3 0.0012014 0 0.0012013199999999999 0 0.00120142 3.3 0.00120134 3.3 0.00120144 0 0.0012013599999999998 0 0.00120146 3.3 0.00120138 3.3 0.00120148 0 0.0012013999999999998 0 0.0012014999999999999 3.3 0.00120142 3.3 0.00120152 0 0.00120144 0 0.00120154 3.3 0.00120146 3.3 0.00120156 0 0.00120148 0 0.00120158 3.3 0.0012014999999999999 3.3 0.0012016 0 0.00120152 0 0.00120162 3.3 0.0012015399999999999 3.3 0.00120164 0 0.00120156 0 0.00120166 3.3 0.0012015799999999998 3.3 0.00120168 0 0.0012016 0 0.0012017 3.3 0.0012016199999999998 3.3 0.0012017199999999999 0 0.00120164 0 0.00120174 3.3 0.00120166 3.3 0.00120176 0 0.00120168 0 0.00120178 3.3 0.0012017 3.3 0.0012018 0 0.0012017199999999999 0 0.00120182 3.3 0.00120174 3.3 0.00120184 0 0.0012017599999999999 0 0.00120186 3.3 0.00120178 3.3 0.00120188 0 0.0012017999999999998 0 0.0012018999999999999 3.3 0.00120182 3.3 0.00120192 0 0.00120184 0 0.00120194 3.3 0.00120186 3.3 0.00120196 0 0.00120188 0 0.00120198 3.3 0.0012018999999999999 3.3 0.001202 0 0.00120192 0 0.00120202 3.3 0.0012019399999999999 3.3 0.00120204 0 0.00120196 0 0.00120206 3.3 0.0012019799999999998 3.3 0.00120208 0 0.001202 0 0.0012021 3.3 0.0012020199999999998 3.3 0.0012021199999999999 0 0.00120204 0 0.00120214 3.3 0.00120206 3.3 0.00120216 0 0.00120208 0 0.00120218 3.3 0.0012021 3.3 0.0012022 0 0.0012021199999999999 0 0.00120222 3.3 0.00120214 3.3 0.00120224 0 0.0012021599999999999 0 0.00120226 3.3 0.00120218 3.3 0.00120228 0 0.0012021999999999998 0 0.0012023 3.3 0.00120222 3.3 0.00120232 0 0.0012022399999999998 0 0.0012023399999999999 3.3 0.00120226 3.3 0.00120236 0 0.00120228 0 0.00120238 3.3 0.0012023 3.3 0.0012024 0 0.00120232 0 0.00120242 3.3 0.0012023399999999999 3.3 0.00120244 0 0.00120236 0 0.00120246 3.3 0.0012023799999999999 3.3 0.00120248 0 0.0012024 0 0.0012025 3.3 0.0012024199999999998 3.3 0.0012025199999999999 0 0.00120244 0 0.00120254 3.3 0.0012024599999999998 3.3 0.0012025599999999999 0 0.00120248 0 0.00120258 3.3 0.0012025 3.3 0.0012026 0 0.0012025199999999999 0 0.00120262 3.3 0.00120254 3.3 0.00120264 0 0.0012025599999999999 0 0.00120266 3.3 0.00120258 3.3 0.00120268 0 0.0012025999999999998 0 0.0012027 3.3 0.00120262 3.3 0.00120272 0 0.0012026399999999998 0 0.0012027399999999999 3.3 0.00120266 3.3 0.00120276 0 0.00120268 0 0.00120278 3.3 0.0012027 3.3 0.0012028 0 0.00120272 0 0.00120282 3.3 0.0012027399999999999 3.3 0.00120284 0 0.00120276 0 0.00120286 3.3 0.0012027799999999999 3.3 0.00120288 0 0.0012028 0 0.0012029 3.3 0.0012028199999999998 3.3 0.00120292 0 0.00120284 0 0.00120294 3.3 0.0012028599999999998 3.3 0.0012029599999999999 0 0.00120288 0 0.00120298 3.3 0.0012029 3.3 0.001203 0 0.00120292 0 0.00120302 3.3 0.00120294 3.3 0.00120304 0 0.0012029599999999999 0 0.00120306 3.3 0.00120298 3.3 0.00120308 0 0.0012029999999999999 0 0.0012031 3.3 0.00120302 3.3 0.00120312 0 0.0012030399999999998 0 0.00120314 3.3 0.00120306 3.3 0.00120316 0 0.0012030799999999998 0 0.0012031799999999999 3.3 0.0012031 3.3 0.0012032 0 0.00120312 0 0.00120322 3.3 0.00120314 3.3 0.00120324 0 0.00120316 0 0.00120326 3.3 0.0012031799999999999 3.3 0.00120328 0 0.0012032 0 0.0012033 3.3 0.0012032199999999999 3.3 0.00120332 0 0.00120324 0 0.00120334 3.3 0.0012032599999999998 3.3 0.0012033599999999999 0 0.00120328 0 0.00120338 3.3 0.0012032999999999998 3.3 0.0012033999999999999 0 0.00120332 0 0.00120342 3.3 0.00120334 3.3 0.00120344 0 0.0012033599999999999 0 0.00120346 3.3 0.00120338 3.3 0.00120348 0 0.0012033999999999999 0 0.0012035 3.3 0.00120342 3.3 0.00120352 0 0.0012034399999999998 0 0.00120354 3.3 0.00120346 3.3 0.00120356 0 0.0012034799999999998 0 0.0012035799999999999 3.3 0.0012035 3.3 0.0012036 0 0.00120352 0 0.00120362 3.3 0.00120354 3.3 0.00120364 0 0.00120356 0 0.00120366 3.3 0.0012035799999999999 3.3 0.00120368 0 0.0012036 0 0.0012037 3.3 0.0012036199999999999 3.3 0.00120372 0 0.00120364 0 0.00120374 3.3 0.0012036599999999998 3.3 0.00120376 0 0.00120368 0 0.00120378 3.3 0.0012036999999999998 3.3 0.0012037999999999999 0 0.00120372 0 0.00120382 3.3 0.00120374 3.3 0.00120384 0 0.00120376 0 0.00120386 3.3 0.00120378 3.3 0.00120388 0 0.0012037999999999999 0 0.0012039 3.3 0.00120382 3.3 0.00120392 0 0.0012038399999999999 0 0.00120394 3.3 0.00120386 3.3 0.00120396 0 0.0012038799999999998 0 0.00120398 3.3 0.0012039 3.3 0.001204 0 0.0012039199999999998 0 0.0012040199999999999 3.3 0.00120394 3.3 0.00120404 0 0.00120396 0 0.00120406 3.3 0.00120398 3.3 0.00120408 0 0.001204 0 0.0012041 3.3 0.0012040199999999999 3.3 0.00120412 0 0.00120404 0 0.00120414 3.3 0.0012040599999999999 3.3 0.00120416 0 0.00120408 0 0.00120418 3.3 0.0012040999999999998 3.3 0.0012041999999999999 0 0.00120412 0 0.00120422 3.3 0.0012041399999999998 3.3 0.0012042399999999999 0 0.00120416 0 0.00120426 3.3 0.00120418 3.3 0.00120428 0 0.0012041999999999999 0 0.0012043 3.3 0.00120422 3.3 0.00120432 0 0.0012042399999999999 0 0.00120434 3.3 0.00120426 3.3 0.00120436 0 0.0012042799999999998 0 0.00120438 3.3 0.0012043 3.3 0.0012044 0 0.0012043199999999998 0 0.0012044199999999999 3.3 0.00120434 3.3 0.00120444 0 0.00120436 0 0.00120446 3.3 0.00120438 3.3 0.00120448 0 0.0012044 0 0.0012045 3.3 0.0012044199999999999 3.3 0.00120452 0 0.00120444 0 0.00120454 3.3 0.0012044599999999999 3.3 0.00120456 0 0.00120448 0 0.00120458 3.3 0.0012044999999999998 3.3 0.0012046 0 0.00120452 0 0.00120462 3.3 0.0012045399999999998 3.3 0.0012046399999999999 0 0.00120456 0 0.00120466 3.3 0.00120458 3.3 0.00120468 0 0.0012046 0 0.0012047 3.3 0.00120462 3.3 0.00120472 0 0.0012046399999999999 0 0.00120474 3.3 0.00120466 3.3 0.00120476 0 0.0012046799999999999 0 0.00120478 3.3 0.0012047 3.3 0.0012048 0 0.0012047199999999998 0 0.00120482 3.3 0.00120474 3.3 0.00120484 0 0.0012047599999999998 0 0.0012048599999999999 3.3 0.00120478 3.3 0.00120488 0 0.0012048 0 0.0012049 3.3 0.00120482 3.3 0.00120492 0 0.00120484 0 0.00120494 3.3 0.0012048599999999999 3.3 0.00120496 0 0.00120488 0 0.00120498 3.3 0.0012048999999999999 3.3 0.001205 0 0.00120492 0 0.00120502 3.3 0.0012049399999999998 3.3 0.0012050399999999999 0 0.00120496 0 0.00120506 3.3 0.00120498 3.3 0.00120508 0 0.001205 0 0.0012051 3.3 0.00120502 3.3 0.00120512 0 0.0012050399999999999 0 0.00120514 3.3 0.00120506 3.3 0.00120516 0 0.0012050799999999999 0 0.00120518 3.3 0.0012051 3.3 0.0012052 0 0.0012051199999999998 0 0.00120522 3.3 0.00120514 3.3 0.00120524 0 0.0012051599999999998 0 0.0012052599999999999 3.3 0.00120518 3.3 0.00120528 0 0.0012052 0 0.0012053 3.3 0.00120522 3.3 0.00120532 0 0.00120524 0 0.00120534 3.3 0.0012052599999999999 3.3 0.00120536 0 0.00120528 0 0.00120538 3.3 0.0012052999999999999 3.3 0.0012054 0 0.00120532 0 0.00120542 3.3 0.0012053399999999998 3.3 0.00120544 0 0.00120536 0 0.00120546 3.3 0.0012053799999999998 3.3 0.0012054799999999999 0 0.0012054 0 0.0012055 3.3 0.00120542 3.3 0.00120552 0 0.00120544 0 0.00120554 3.3 0.00120546 3.3 0.00120556 0 0.0012054799999999999 0 0.00120558 3.3 0.0012055 3.3 0.0012056 0 0.0012055199999999999 0 0.00120562 3.3 0.00120554 3.3 0.00120564 0 0.0012055599999999998 0 0.0012056599999999999 3.3 0.00120558 3.3 0.00120568 0 0.0012055999999999998 0 0.0012056999999999999 3.3 0.00120562 3.3 0.00120572 0 0.00120564 0 0.00120574 3.3 0.0012056599999999999 3.3 0.00120576 0 0.00120568 0 0.00120578 3.3 0.0012056999999999999 3.3 0.0012058 0 0.00120572 0 0.00120582 3.3 0.0012057399999999999 3.3 0.00120584 0 0.00120576 0 0.00120586 3.3 0.0012057799999999998 3.3 0.0012058799999999999 0 0.0012058 0 0.0012059 3.3 0.00120582 3.3 0.00120592 0 0.00120584 0 0.00120594 3.3 0.00120586 3.3 0.00120596 0 0.0012058799999999999 0 0.00120598 3.3 0.0012059 3.3 0.001206 0 0.0012059199999999999 0 0.00120602 3.3 0.00120594 3.3 0.00120604 0 0.0012059599999999998 0 0.00120606 3.3 0.00120598 3.3 0.00120608 0 0.0012059999999999998 0 0.0012060999999999999 3.3 0.00120602 3.3 0.00120612 0 0.00120604 0 0.00120614 3.3 0.00120606 3.3 0.00120616 0 0.00120608 0 0.00120618 3.3 0.0012060999999999999 3.3 0.0012062 0 0.00120612 0 0.00120622 3.3 0.0012061399999999999 3.3 0.00120624 0 0.00120616 0 0.00120626 3.3 0.0012061799999999998 3.3 0.00120628 0 0.0012062 0 0.0012063 3.3 0.0012062199999999998 3.3 0.0012063199999999999 0 0.00120624 0 0.00120634 3.3 0.00120626 3.3 0.00120636 0 0.00120628 0 0.00120638 3.3 0.0012063 3.3 0.0012064 0 0.0012063199999999999 0 0.00120642 3.3 0.00120634 3.3 0.00120644 0 0.0012063599999999999 0 0.00120646 3.3 0.00120638 3.3 0.00120648 0 0.0012063999999999998 0 0.0012064999999999999 3.3 0.00120642 3.3 0.00120652 0 0.0012064399999999998 0 0.0012065399999999999 3.3 0.00120646 3.3 0.00120656 0 0.00120648 0 0.00120658 3.3 0.0012064999999999999 3.3 0.0012066 0 0.00120652 0 0.00120662 3.3 0.0012065399999999999 3.3 0.00120664 0 0.00120656 0 0.00120666 3.3 0.0012065799999999998 3.3 0.00120668 0 0.0012066 0 0.0012067 3.3 0.0012066199999999998 3.3 0.0012067199999999999 0 0.00120664 0 0.00120674 3.3 0.00120666 3.3 0.00120676 0 0.00120668 0 0.00120678 3.3 0.0012067 3.3 0.0012068 0 0.0012067199999999999 0 0.00120682 3.3 0.00120674 3.3 0.00120684 0 0.0012067599999999999 0 0.00120686 3.3 0.00120678 3.3 0.00120688 0 0.0012067999999999998 0 0.0012069 3.3 0.00120682 3.3 0.00120692 0 0.0012068399999999998 0 0.0012069399999999999 3.3 0.00120686 3.3 0.00120696 0 0.00120688 0 0.00120698 3.3 0.0012069 3.3 0.001207 0 0.00120692 0 0.00120702 3.3 0.0012069399999999999 3.3 0.00120704 0 0.00120696 0 0.00120706 3.3 0.0012069799999999999 3.3 0.00120708 0 0.001207 0 0.0012071 3.3 0.0012070199999999998 3.3 0.00120712 0 0.00120704 0 0.00120714 3.3 0.0012070599999999998 3.3 0.0012071599999999999 0 0.00120708 0 0.00120718 3.3 0.0012071 3.3 0.0012072 0 0.00120712 0 0.00120722 3.3 0.00120714 3.3 0.00120724 0 0.0012071599999999999 0 0.00120726 3.3 0.00120718 3.3 0.00120728 0 0.0012071999999999999 0 0.0012073 3.3 0.00120722 3.3 0.00120732 0 0.0012072399999999998 0 0.0012073399999999999 3.3 0.00120726 3.3 0.00120736 0 0.0012072799999999998 0 0.0012073799999999999 3.3 0.0012073 3.3 0.0012074 0 0.00120732 0 0.00120742 3.3 0.0012073399999999999 3.3 0.00120744 0 0.00120736 0 0.00120746 3.3 0.0012073799999999999 3.3 0.00120748 0 0.0012074 0 0.0012075 3.3 0.0012074199999999998 3.3 0.00120752 0 0.00120744 0 0.00120754 3.3 0.0012074599999999998 3.3 0.0012075599999999999 0 0.00120748 0 0.00120758 3.3 0.0012075 3.3 0.0012076 0 0.00120752 0 0.00120762 3.3 0.00120754 3.3 0.00120764 0 0.0012075599999999999 0 0.00120766 3.3 0.00120758 3.3 0.00120768 0 0.0012075999999999999 0 0.0012077 3.3 0.00120762 3.3 0.00120772 0 0.0012076399999999998 0 0.00120774 3.3 0.00120766 3.3 0.00120776 0 0.0012076799999999998 0 0.0012077799999999999 3.3 0.0012077 3.3 0.0012078 0 0.00120772 0 0.00120782 3.3 0.00120774 3.3 0.00120784 0 0.00120776 0 0.00120786 3.3 0.0012077799999999999 3.3 0.00120788 0 0.0012078 0 0.0012079 3.3 0.0012078199999999999 3.3 0.00120792 0 0.00120784 0 0.00120794 3.3 0.0012078599999999998 3.3 0.00120796 0 0.00120788 0 0.00120798 3.3 0.0012078999999999998 3.3 0.0012079999999999999 0 0.00120792 0 0.00120802 3.3 0.00120794 3.3 0.00120804 0 0.00120796 0 0.00120806 3.3 0.00120798 3.3 0.00120808 0 0.0012079999999999999 0 0.0012081 3.3 0.00120802 3.3 0.00120812 0 0.0012080399999999999 0 0.00120814 3.3 0.00120806 3.3 0.00120816 0 0.0012080799999999998 0 0.0012081799999999999 3.3 0.0012081 3.3 0.0012082 0 0.00120812 0 0.00120822 3.3 0.00120814 3.3 0.00120824 0 0.00120816 0 0.00120826 3.3 0.0012081799999999999 3.3 0.00120828 0 0.0012082 0 0.0012083 3.3 0.0012082199999999999 3.3 0.00120832 0 0.00120824 0 0.00120834 3.3 0.0012082599999999998 3.3 0.00120836 0 0.00120828 0 0.00120838 3.3 0.0012082999999999998 3.3 0.0012083999999999999 0 0.00120832 0 0.00120842 3.3 0.00120834 3.3 0.00120844 0 0.00120836 0 0.00120846 3.3 0.00120838 3.3 0.00120848 0 0.0012083999999999999 0 0.0012085 3.3 0.00120842 3.3 0.00120852 0 0.0012084399999999999 0 0.00120854 3.3 0.00120846 3.3 0.00120856 0 0.0012084799999999998 0 0.00120858 3.3 0.0012085 3.3 0.0012086 0 0.0012085199999999998 0 0.0012086199999999999 3.3 0.00120854 3.3 0.00120864 0 0.00120856 0 0.00120866 3.3 0.00120858 3.3 0.00120868 0 0.0012086 0 0.0012087 3.3 0.0012086199999999999 3.3 0.00120872 0 0.00120864 0 0.00120874 3.3 0.0012086599999999999 3.3 0.00120876 0 0.00120868 0 0.00120878 3.3 0.0012086999999999998 3.3 0.0012088 0 0.00120872 0 0.00120882 3.3 0.0012087399999999998 3.3 0.0012088399999999999 0 0.00120876 0 0.00120886 3.3 0.00120878 3.3 0.00120888 0 0.0012088 0 0.0012089 3.3 0.00120882 3.3 0.00120892 0 0.0012088399999999999 0 0.00120894 3.3 0.00120886 3.3 0.00120896 0 0.0012088799999999999 0 0.00120898 3.3 0.0012089 3.3 0.001209 0 0.0012089199999999998 0 0.0012090199999999999 3.3 0.00120894 3.3 0.00120904 0 0.00120896 0 0.00120906 3.3 0.00120898 3.3 0.00120908 0 0.001209 0 0.0012091 3.3 0.0012090199999999999 3.3 0.00120912 0 0.00120904 0 0.00120914 3.3 0.0012090599999999999 3.3 0.00120916 0 0.00120908 0 0.00120918 3.3 0.0012090999999999998 3.3 0.0012092 0 0.00120912 0 0.00120922 3.3 0.0012091399999999998 3.3 0.0012092399999999999 0 0.00120916 0 0.00120926 3.3 0.00120918 3.3 0.00120928 0 0.0012092 0 0.0012093 3.3 0.00120922 3.3 0.00120932 0 0.0012092399999999999 0 0.00120934 3.3 0.00120926 3.3 0.00120936 0 0.0012092799999999999 0 0.00120938 3.3 0.0012093 3.3 0.0012094 0 0.0012093199999999998 0 0.00120942 3.3 0.00120934 3.3 0.00120944 0 0.0012093599999999998 0 0.0012094599999999999 3.3 0.00120938 3.3 0.00120948 0 0.0012094 0 0.0012095 3.3 0.00120942 3.3 0.00120952 0 0.00120944 0 0.00120954 3.3 0.0012094599999999999 3.3 0.00120956 0 0.00120948 0 0.00120958 3.3 0.0012094999999999999 3.3 0.0012096 0 0.00120952 0 0.00120962 3.3 0.0012095399999999998 3.3 0.0012096399999999999 0 0.00120956 0 0.00120966 3.3 0.0012095799999999998 3.3 0.0012096799999999999 0 0.0012096 0 0.0012097 3.3 0.00120962 3.3 0.00120972 0 0.0012096399999999999 0 0.00120974 3.3 0.00120966 3.3 0.00120976 0 0.0012096799999999999 0 0.00120978 3.3 0.0012097 3.3 0.0012098 0 0.0012097199999999998 0 0.00120982 3.3 0.00120974 3.3 0.00120984 0 0.0012097599999999998 0 0.0012098599999999999 3.3 0.00120978 3.3 0.00120988 0 0.0012098 0 0.0012099 3.3 0.00120982 3.3 0.00120992 0 0.00120984 0 0.00120994 3.3 0.0012098599999999999 3.3 0.00120996 0 0.00120988 0 0.00120998 3.3 0.0012098999999999999 3.3 0.00121 0 0.00120992 0 0.00121002 3.3 0.0012099399999999998 3.3 0.00121004 0 0.00120996 0 0.00121006 3.3 0.0012099799999999998 3.3 0.0012100799999999999 0 0.00121 0 0.0012101 3.3 0.00121002 3.3 0.00121012 0 0.00121004 0 0.00121014 3.3 0.00121006 3.3 0.00121016 0 0.0012100799999999999 0 0.00121018 3.3 0.0012101 3.3 0.0012102 0 0.0012101199999999999 0 0.00121022 3.3 0.00121014 3.3 0.00121024 0 0.0012101599999999998 0 0.00121026 3.3 0.00121018 3.3 0.00121028 0 0.0012101999999999998 0 0.0012102999999999999 3.3 0.00121022 3.3 0.00121032 0 0.00121024 0 0.00121034 3.3 0.00121026 3.3 0.00121036 0 0.00121028 0 0.00121038 3.3 0.0012102999999999999 3.3 0.0012104 0 0.00121032 0 0.00121042 3.3 0.0012103399999999999 3.3 0.00121044 0 0.00121036 0 0.00121046 3.3 0.0012103799999999998 3.3 0.0012104799999999999 0 0.0012104 0 0.0012105 3.3 0.0012104199999999998 3.3 0.0012105199999999999 0 0.00121044 0 0.00121054 3.3 0.00121046 3.3 0.00121056 0 0.0012104799999999999 0 0.00121058 3.3 0.0012105 3.3 0.0012106 0 0.0012105199999999999 0 0.00121062 3.3 0.00121054 3.3 0.00121064 0 0.0012105599999999998 0 0.00121066 3.3 0.00121058 3.3 0.00121068 0 0.0012105999999999998 0 0.0012106999999999999 3.3 0.00121062 3.3 0.00121072 0 0.00121064 0 0.00121074 3.3 0.00121066 3.3 0.00121076 0 0.00121068 0 0.00121078 3.3 0.0012106999999999999 3.3 0.0012108 0 0.00121072 0 0.00121082 3.3 0.0012107399999999999 3.3 0.00121084 0 0.00121076 0 0.00121086 3.3 0.0012107799999999998 3.3 0.00121088 0 0.0012108 0 0.0012109 3.3 0.0012108199999999998 3.3 0.0012109199999999999 0 0.00121084 0 0.00121094 3.3 0.00121086 3.3 0.00121096 0 0.00121088 0 0.00121098 3.3 0.0012109 3.3 0.001211 0 0.0012109199999999999 0 0.00121102 3.3 0.00121094 3.3 0.00121104 0 0.0012109599999999999 0 0.00121106 3.3 0.00121098 3.3 0.00121108 0 0.0012109999999999998 0 0.0012111 3.3 0.00121102 3.3 0.00121112 0 0.0012110399999999998 0 0.0012111399999999999 3.3 0.00121106 3.3 0.00121116 0 0.00121108 0 0.00121118 3.3 0.0012111 3.3 0.0012112 0 0.00121112 0 0.00121122 3.3 0.0012111399999999999 3.3 0.00121124 0 0.00121116 0 0.00121126 3.3 0.0012111799999999999 3.3 0.00121128 0 0.0012112 0 0.0012113 3.3 0.0012112199999999998 3.3 0.0012113199999999999 0 0.00121124 0 0.00121134 3.3 0.0012112599999999998 3.3 0.0012113599999999999 0 0.00121128 0 0.00121138 3.3 0.0012113 3.3 0.0012114 0 0.0012113199999999999 0 0.00121142 3.3 0.00121134 3.3 0.00121144 0 0.0012113599999999999 0 0.00121146 3.3 0.00121138 3.3 0.00121148 0 0.0012113999999999998 0 0.0012115 3.3 0.00121142 3.3 0.00121152 0 0.0012114399999999998 0 0.0012115399999999999 3.3 0.00121146 3.3 0.00121156 0 0.00121148 0 0.00121158 3.3 0.0012115 3.3 0.0012116 0 0.00121152 0 0.00121162 3.3 0.0012115399999999999 3.3 0.00121164 0 0.00121156 0 0.00121166 3.3 0.0012115799999999999 3.3 0.00121168 0 0.0012116 0 0.0012117 3.3 0.0012116199999999998 3.3 0.00121172 0 0.00121164 0 0.00121174 3.3 0.0012116599999999998 3.3 0.0012117599999999999 0 0.00121168 0 0.00121178 3.3 0.0012117 3.3 0.0012118 0 0.00121172 0 0.00121182 3.3 0.00121174 3.3 0.00121184 0 0.0012117599999999999 0 0.00121186 3.3 0.00121178 3.3 0.00121188 0 0.0012117999999999999 0 0.0012119 3.3 0.00121182 3.3 0.00121192 0 0.0012118399999999998 0 0.00121194 3.3 0.00121186 3.3 0.00121196 0 0.0012118799999999998 0 0.0012119799999999999 3.3 0.0012119 3.3 0.001212 0 0.00121192 0 0.00121202 3.3 0.00121194 3.3 0.00121204 0 0.00121196 0 0.00121206 3.3 0.0012119799999999999 3.3 0.00121208 0 0.001212 0 0.0012121 3.3 0.0012120199999999999 3.3 0.00121212 0 0.00121204 0 0.00121214 3.3 0.0012120599999999998 3.3 0.0012121599999999999 0 0.00121208 0 0.00121218 3.3 0.0012121 3.3 0.0012122 0 0.00121212 0 0.00121222 3.3 0.00121214 3.3 0.00121224 0 0.0012121599999999999 0 0.00121226 3.3 0.00121218 3.3 0.00121228 0 0.0012121999999999999 0 0.0012123 3.3 0.00121222 3.3 0.00121232 0 0.0012122399999999998 0 0.00121234 3.3 0.00121226 3.3 0.00121236 0 0.0012122799999999998 0 0.0012123799999999999 3.3 0.0012123 3.3 0.0012124 0 0.00121232 0 0.00121242 3.3 0.00121234 3.3 0.00121244 0 0.00121236 0 0.00121246 3.3 0.0012123799999999999 3.3 0.00121248 0 0.0012124 0 0.0012125 3.3 0.0012124199999999999 3.3 0.00121252 0 0.00121244 0 0.00121254 3.3 0.0012124599999999998 3.3 0.00121256 0 0.00121248 0 0.00121258 3.3 0.0012124999999999998 3.3 0.0012125999999999999 0 0.00121252 0 0.00121262 3.3 0.00121254 3.3 0.00121264 0 0.00121256 0 0.00121266 3.3 0.00121258 3.3 0.00121268 0 0.0012125999999999999 0 0.0012127 3.3 0.00121262 3.3 0.00121272 0 0.0012126399999999999 0 0.00121274 3.3 0.00121266 3.3 0.00121276 0 0.0012126799999999998 0 0.0012127799999999999 3.3 0.0012127 3.3 0.0012128 0 0.0012127199999999998 0 0.0012128199999999999 3.3 0.00121274 3.3 0.00121284 0 0.00121276 0 0.00121286 3.3 0.0012127799999999999 3.3 0.00121288 0 0.0012128 0 0.0012129 3.3 0.0012128199999999999 3.3 0.00121292 0 0.00121284 0 0.00121294 3.3 0.0012128599999999998 3.3 0.00121296 0 0.00121288 0 0.00121298 3.3 0.0012128999999999998 3.3 0.0012129999999999999 0 0.00121292 0 0.00121302 3.3 0.00121294 3.3 0.00121304 0 0.00121296 0 0.00121306 3.3 0.00121298 3.3 0.00121308 0 0.0012129999999999999 0 0.0012131 3.3 0.00121302 3.3 0.00121312 0 0.0012130399999999999 0 0.00121314 3.3 0.00121306 3.3 0.00121316 0 0.0012130799999999998 0 0.00121318 3.3 0.0012131 3.3 0.0012132 0 0.0012131199999999998 0 0.0012132199999999999 3.3 0.00121314 3.3 0.00121324 0 0.00121316 0 0.00121326 3.3 0.00121318 3.3 0.00121328 0 0.0012132 0 0.0012133 3.3 0.0012132199999999999 3.3 0.00121332 0 0.00121324 0 0.00121334 3.3 0.0012132599999999999 3.3 0.00121336 0 0.00121328 0 0.00121338 3.3 0.0012132999999999998 3.3 0.0012134 0 0.00121332 0 0.00121342 3.3 0.0012133399999999998 3.3 0.0012134399999999999 0 0.00121336 0 0.00121346 3.3 0.00121338 3.3 0.00121348 0 0.0012134 0 0.0012135 3.3 0.00121342 3.3 0.00121352 0 0.0012134399999999999 0 0.00121354 3.3 0.00121346 3.3 0.00121356 0 0.0012134799999999999 0 0.00121358 3.3 0.0012135 3.3 0.0012136 0 0.0012135199999999998 0 0.0012136199999999999 3.3 0.00121354 3.3 0.00121364 0 0.0012135599999999998 0 0.0012136599999999999 3.3 0.00121358 3.3 0.00121368 0 0.0012136 0 0.0012137 3.3 0.0012136199999999999 3.3 0.00121372 0 0.00121364 0 0.00121374 3.3 0.0012136599999999999 3.3 0.00121376 0 0.00121368 0 0.00121378 3.3 0.0012136999999999998 3.3 0.0012138 0 0.00121372 0 0.00121382 3.3 0.0012137399999999998 3.3 0.0012138399999999999 0 0.00121376 0 0.00121386 3.3 0.00121378 3.3 0.00121388 0 0.0012138 0 0.0012139 3.3 0.00121382 3.3 0.00121392 0 0.0012138399999999999 0 0.00121394 3.3 0.00121386 3.3 0.00121396 0 0.0012138799999999999 0 0.00121398 3.3 0.0012139 3.3 0.001214 0 0.0012139199999999998 0 0.00121402 3.3 0.00121394 3.3 0.00121404 0 0.0012139599999999998 0 0.0012140599999999999 3.3 0.00121398 3.3 0.00121408 0 0.001214 0 0.0012141 3.3 0.00121402 3.3 0.00121412 0 0.00121404 0 0.00121414 3.3 0.0012140599999999999 3.3 0.00121416 0 0.00121408 0 0.00121418 3.3 0.0012140999999999999 3.3 0.0012142 0 0.00121412 0 0.00121422 3.3 0.0012141399999999998 3.3 0.00121424 0 0.00121416 0 0.00121426 3.3 0.0012141799999999998 3.3 0.0012142799999999999 0 0.0012142 0 0.0012143 3.3 0.00121422 3.3 0.00121432 0 0.00121424 0 0.00121434 3.3 0.00121426 3.3 0.00121436 0 0.0012142799999999999 0 0.00121438 3.3 0.0012143 3.3 0.0012144 0 0.0012143199999999999 0 0.00121442 3.3 0.00121434 3.3 0.00121444 0 0.0012143599999999998 0 0.0012144599999999999 3.3 0.00121438 3.3 0.00121448 0 0.0012143999999999998 0 0.0012144999999999999 3.3 0.00121442 3.3 0.00121452 0 0.00121444 0 0.00121454 3.3 0.0012144599999999999 3.3 0.00121456 0 0.00121448 0 0.00121458 3.3 0.0012144999999999999 3.3 0.0012146 0 0.00121452 0 0.00121462 3.3 0.0012145399999999998 3.3 0.00121464 0 0.00121456 0 0.00121466 3.3 0.0012145799999999998 3.3 0.0012146799999999999 0 0.0012146 0 0.0012147 3.3 0.00121462 3.3 0.00121472 0 0.00121464 0 0.00121474 3.3 0.00121466 3.3 0.00121476 0 0.0012146799999999999 0 0.00121478 3.3 0.0012147 3.3 0.0012148 0 0.0012147199999999999 0 0.00121482 3.3 0.00121474 3.3 0.00121484 0 0.0012147599999999998 0 0.00121486 3.3 0.00121478 3.3 0.00121488 0 0.0012147999999999998 0 0.0012148999999999999 3.3 0.00121482 3.3 0.00121492 0 0.00121484 0 0.00121494 3.3 0.00121486 3.3 0.00121496 0 0.00121488 0 0.00121498 3.3 0.0012148999999999999 3.3 0.001215 0 0.00121492 0 0.00121502 3.3 0.0012149399999999999 3.3 0.00121504 0 0.00121496 0 0.00121506 3.3 0.0012149799999999998 3.3 0.00121508 0 0.001215 0 0.0012151 3.3 0.0012150199999999998 3.3 0.0012151199999999999 0 0.00121504 0 0.00121514 3.3 0.00121506 3.3 0.00121516 0 0.00121508 0 0.00121518 3.3 0.0012151 3.3 0.0012152 0 0.0012151199999999999 0 0.00121522 3.3 0.00121514 3.3 0.00121524 0 0.0012151599999999999 0 0.00121526 3.3 0.00121518 3.3 0.00121528 0 0.0012151999999999998 0 0.0012152999999999999 3.3 0.00121522 3.3 0.00121532 0 0.00121524 0 0.00121534 3.3 0.00121526 3.3 0.00121536 0 0.00121528 0 0.00121538 3.3 0.0012152999999999999 3.3 0.0012154 0 0.00121532 0 0.00121542 3.3 0.0012153399999999999 3.3 0.00121544 0 0.00121536 0 0.00121546 3.3 0.0012153799999999998 3.3 0.00121548 0 0.0012154 0 0.0012155 3.3 0.0012154199999999998 3.3 0.0012155199999999999 0 0.00121544 0 0.00121554 3.3 0.00121546 3.3 0.00121556 0 0.00121548 0 0.00121558 3.3 0.0012155 3.3 0.0012156 0 0.0012155199999999999 0 0.00121562 3.3 0.00121554 3.3 0.00121564 0 0.0012155599999999999 0 0.00121566 3.3 0.00121558 3.3 0.00121568 0 0.0012155999999999998 0 0.0012157 3.3 0.00121562 3.3 0.00121572 0 0.0012156399999999998 0 0.0012157399999999999 3.3 0.00121566 3.3 0.00121576 0 0.00121568 0 0.00121578 3.3 0.0012157 3.3 0.0012158 0 0.00121572 0 0.00121582 3.3 0.0012157399999999999 3.3 0.00121584 0 0.00121576 0 0.00121586 3.3 0.0012157799999999999 3.3 0.00121588 0 0.0012158 0 0.0012159 3.3 0.0012158199999999998 3.3 0.0012159199999999999 0 0.00121584 0 0.00121594 3.3 0.0012158599999999998 3.3 0.0012159599999999999 0 0.00121588 0 0.00121598 3.3 0.0012159 3.3 0.001216 0 0.0012159199999999999 0 0.00121602 3.3 0.00121594 3.3 0.00121604 0 0.0012159599999999999 0 0.00121606 3.3 0.00121598 3.3 0.00121608 0 0.0012159999999999999 0 0.0012161 3.3 0.00121602 3.3 0.00121612 0 0.0012160399999999998 0 0.0012161399999999999 3.3 0.00121606 3.3 0.00121616 0 0.00121608 0 0.00121618 3.3 0.0012161 3.3 0.0012162 0 0.00121612 0 0.00121622 3.3 0.0012161399999999999 3.3 0.00121624 0 0.00121616 0 0.00121626 3.3 0.0012161799999999999 3.3 0.00121628 0 0.0012162 0 0.0012163 3.3 0.0012162199999999998 3.3 0.00121632 0 0.00121624 0 0.00121634 3.3 0.0012162599999999998 3.3 0.0012163599999999999 0 0.00121628 0 0.00121638 3.3 0.0012163 3.3 0.0012164 0 0.00121632 0 0.00121642 3.3 0.00121634 3.3 0.00121644 0 0.0012163599999999999 0 0.00121646 3.3 0.00121638 3.3 0.00121648 0 0.0012163999999999999 0 0.0012165 3.3 0.00121642 3.3 0.00121652 0 0.0012164399999999998 0 0.00121654 3.3 0.00121646 3.3 0.00121656 0 0.0012164799999999998 0 0.0012165799999999999 3.3 0.0012165 3.3 0.0012166 0 0.00121652 0 0.00121662 3.3 0.00121654 3.3 0.00121664 0 0.00121656 0 0.00121666 3.3 0.0012165799999999999 3.3 0.00121668 0 0.0012166 0 0.0012167 3.3 0.0012166199999999999 3.3 0.00121672 0 0.00121664 0 0.00121674 3.3 0.0012166599999999998 3.3 0.0012167599999999999 0 0.00121668 0 0.00121678 3.3 0.0012166999999999998 3.3 0.0012167999999999999 0 0.00121672 0 0.00121682 3.3 0.00121674 3.3 0.00121684 0 0.0012167599999999999 0 0.00121686 3.3 0.00121678 3.3 0.00121688 0 0.0012167999999999999 0 0.0012169 3.3 0.00121682 3.3 0.00121692 0 0.0012168399999999998 0 0.00121694 3.3 0.00121686 3.3 0.00121696 0 0.0012168799999999998 0 0.0012169799999999999 3.3 0.0012169 3.3 0.001217 0 0.00121692 0 0.00121702 3.3 0.00121694 3.3 0.00121704 0 0.00121696 0 0.00121706 3.3 0.0012169799999999999 3.3 0.00121708 0 0.001217 0 0.0012171 3.3 0.0012170199999999999 3.3 0.00121712 0 0.00121704 0 0.00121714 3.3 0.0012170599999999998 3.3 0.00121716 0 0.00121708 0 0.00121718 3.3 0.0012170999999999998 3.3 0.0012171999999999999 0 0.00121712 0 0.00121722 3.3 0.00121714 3.3 0.00121724 0 0.00121716 0 0.00121726 3.3 0.00121718 3.3 0.00121728 0 0.0012171999999999999 0 0.0012173 3.3 0.00121722 3.3 0.00121732 0 0.0012172399999999999 0 0.00121734 3.3 0.00121726 3.3 0.00121736 0 0.0012172799999999998 0 0.00121738 3.3 0.0012173 3.3 0.0012174 0 0.0012173199999999998 0 0.0012174199999999999 3.3 0.00121734 3.3 0.00121744 0 0.00121736 0 0.00121746 3.3 0.00121738 3.3 0.00121748 0 0.0012174 0 0.0012175 3.3 0.0012174199999999999 3.3 0.00121752 0 0.00121744 0 0.00121754 3.3 0.0012174599999999999 3.3 0.00121756 0 0.00121748 0 0.00121758 3.3 0.0012174999999999998 3.3 0.0012175999999999999 0 0.00121752 0 0.00121762 3.3 0.0012175399999999998 3.3 0.0012176399999999999 0 0.00121756 0 0.00121766 3.3 0.00121758 3.3 0.00121768 0 0.0012175999999999999 0 0.0012177 3.3 0.00121762 3.3 0.00121772 0 0.0012176399999999999 0 0.00121774 3.3 0.00121766 3.3 0.00121776 0 0.0012176799999999998 0 0.00121778 3.3 0.0012177 3.3 0.0012178 0 0.0012177199999999998 0 0.0012178199999999999 3.3 0.00121774 3.3 0.00121784 0 0.00121776 0 0.00121786 3.3 0.00121778 3.3 0.00121788 0 0.0012178 0 0.0012179 3.3 0.0012178199999999999 3.3 0.00121792 0 0.00121784 0 0.00121794 3.3 0.0012178599999999999 3.3 0.00121796 0 0.00121788 0 0.00121798 3.3 0.0012178999999999998 3.3 0.001218 0 0.00121792 0 0.00121802 3.3 0.0012179399999999998 3.3 0.0012180399999999999 0 0.00121796 0 0.00121806 3.3 0.00121798 3.3 0.00121808 0 0.001218 0 0.0012181 3.3 0.00121802 3.3 0.00121812 0 0.0012180399999999999 0 0.00121814 3.3 0.00121806 3.3 0.00121816 0 0.0012180799999999999 0 0.00121818 3.3 0.0012181 3.3 0.0012182 0 0.0012181199999999998 0 0.00121822 3.3 0.00121814 3.3 0.00121824 0 0.0012181599999999998 0 0.0012182599999999999 3.3 0.00121818 3.3 0.00121828 0 0.0012182 0 0.0012183 3.3 0.00121822 3.3 0.00121832 0 0.00121824 0 0.00121834 3.3 0.0012182599999999999 3.3 0.00121836 0 0.00121828 0 0.00121838 3.3 0.0012182999999999999 3.3 0.0012184 0 0.00121832 0 0.00121842 3.3 0.0012183399999999998 3.3 0.0012184399999999999 0 0.00121836 0 0.00121846 3.3 0.00121838 3.3 0.00121848 0 0.0012184 0 0.0012185 3.3 0.00121842 3.3 0.00121852 0 0.0012184399999999999 0 0.00121854 3.3 0.00121846 3.3 0.00121856 0 0.0012184799999999999 0 0.00121858 3.3 0.0012185 3.3 0.0012186 0 0.0012185199999999998 0 0.00121862 3.3 0.00121854 3.3 0.00121864 0 0.0012185599999999998 0 0.0012186599999999999 3.3 0.00121858 3.3 0.00121868 0 0.0012186 0 0.0012187 3.3 0.00121862 3.3 0.00121872 0 0.00121864 0 0.00121874 3.3 0.0012186599999999999 3.3 0.00121876 0 0.00121868 0 0.00121878 3.3 0.0012186999999999999 3.3 0.0012188 0 0.00121872 0 0.00121882 3.3 0.0012187399999999998 3.3 0.00121884 0 0.00121876 0 0.00121886 3.3 0.0012187799999999998 3.3 0.0012188799999999999 0 0.0012188 0 0.0012189 3.3 0.00121882 3.3 0.00121892 0 0.00121884 0 0.00121894 3.3 0.00121886 3.3 0.00121896 0 0.0012188799999999999 0 0.00121898 3.3 0.0012189 3.3 0.001219 0 0.0012189199999999999 0 0.00121902 3.3 0.00121894 3.3 0.00121904 0 0.0012189599999999998 0 0.00121906 3.3 0.00121898 3.3 0.00121908 0 0.0012189999999999998 0 0.0012190999999999999 3.3 0.00121902 3.3 0.00121912 0 0.00121904 0 0.00121914 3.3 0.00121906 3.3 0.00121916 0 0.00121908 0 0.00121918 3.3 0.0012190999999999999 3.3 0.0012192 0 0.00121912 0 0.00121922 3.3 0.0012191399999999999 3.3 0.00121924 0 0.00121916 0 0.00121926 3.3 0.0012191799999999998 3.3 0.0012192799999999999 0 0.0012192 0 0.0012193 3.3 0.00121922 3.3 0.00121932 0 0.00121924 0 0.00121934 3.3 0.00121926 3.3 0.00121936 0 0.0012192799999999999 0 0.00121938 3.3 0.0012193 3.3 0.0012194 0 0.0012193199999999999 0 0.00121942 3.3 0.00121934 3.3 0.00121944 0 0.0012193599999999998 0 0.00121946 3.3 0.00121938 3.3 0.00121948 0 0.0012193999999999998 0 0.0012194999999999999 3.3 0.00121942 3.3 0.00121952 0 0.00121944 0 0.00121954 3.3 0.00121946 3.3 0.00121956 0 0.00121948 0 0.00121958 3.3 0.0012194999999999999 3.3 0.0012196 0 0.00121952 0 0.00121962 3.3 0.0012195399999999999 3.3 0.00121964 0 0.00121956 0 0.00121966 3.3 0.0012195799999999998 3.3 0.00121968 0 0.0012196 0 0.0012197 3.3 0.0012196199999999998 3.3 0.0012197199999999999 0 0.00121964 0 0.00121974 3.3 0.00121966 3.3 0.00121976 0 0.00121968 0 0.00121978 3.3 0.0012197 3.3 0.0012198 0 0.0012197199999999999 0 0.00121982 3.3 0.00121974 3.3 0.00121984 0 0.0012197599999999999 0 0.00121986 3.3 0.00121978 3.3 0.00121988 0 0.0012197999999999998 0 0.0012198999999999999 3.3 0.00121982 3.3 0.00121992 0 0.0012198399999999998 0 0.0012199399999999999 3.3 0.00121986 3.3 0.00121996 0 0.00121988 0 0.00121998 3.3 0.0012198999999999999 3.3 0.00122 0 0.00121992 0 0.00122002 3.3 0.0012199399999999999 3.3 0.00122004 0 0.00121996 0 0.00122006 3.3 0.0012199799999999998 3.3 0.00122008 0 0.00122 0 0.0012201 3.3 0.0012200199999999998 3.3 0.0012201199999999999 0 0.00122004 0 0.00122014 3.3 0.00122006 3.3 0.00122016 0 0.00122008 0 0.00122018 3.3 0.0012201 3.3 0.0012202 0 0.0012201199999999999 0 0.00122022 3.3 0.00122014 3.3 0.00122024 0 0.0012201599999999999 0 0.00122026 3.3 0.00122018 3.3 0.00122028 0 0.0012201999999999998 0 0.0012203 3.3 0.00122022 3.3 0.00122032 0 0.0012202399999999998 0 0.0012203399999999999 3.3 0.00122026 3.3 0.00122036 0 0.00122028 0 0.00122038 3.3 0.0012203 3.3 0.0012204 0 0.00122032 0 0.00122042 3.3 0.0012203399999999999 3.3 0.00122044 0 0.00122036 0 0.00122046 3.3 0.0012203799999999999 3.3 0.00122048 0 0.0012204 0 0.0012205 3.3 0.0012204199999999998 3.3 0.00122052 0 0.00122044 0 0.00122054 3.3 0.0012204599999999998 3.3 0.0012205599999999999 0 0.00122048 0 0.00122058 3.3 0.0012205 3.3 0.0012206 0 0.00122052 0 0.00122062 3.3 0.00122054 3.3 0.00122064 0 0.0012205599999999999 0 0.00122066 3.3 0.00122058 3.3 0.00122068 0 0.0012205999999999999 0 0.0012207 3.3 0.00122062 3.3 0.00122072 0 0.0012206399999999998 0 0.0012207399999999999 3.3 0.00122066 3.3 0.00122076 0 0.0012206799999999998 0 0.0012207799999999999 3.3 0.0012207 3.3 0.0012208 0 0.00122072 0 0.00122082 3.3 0.0012207399999999999 3.3 0.00122084 0 0.00122076 0 0.00122086 3.3 0.0012207799999999999 3.3 0.00122088 0 0.0012208 0 0.0012209 3.3 0.0012208199999999998 3.3 0.00122092 0 0.00122084 0 0.00122094 3.3 0.0012208599999999998 3.3 0.0012209599999999999 0 0.00122088 0 0.00122098 3.3 0.0012209 3.3 0.001221 0 0.00122092 0 0.00122102 3.3 0.00122094 3.3 0.00122104 0 0.0012209599999999999 0 0.00122106 3.3 0.00122098 3.3 0.00122108 0 0.0012209999999999999 0 0.0012211 3.3 0.00122102 3.3 0.00122112 0 0.0012210399999999998 0 0.00122114 3.3 0.00122106 3.3 0.00122116 0 0.0012210799999999998 0 0.0012211799999999999 3.3 0.0012211 3.3 0.0012212 0 0.00122112 0 0.00122122 3.3 0.00122114 3.3 0.00122124 0 0.00122116 0 0.00122126 3.3 0.0012211799999999999 3.3 0.00122128 0 0.0012212 0 0.0012213 3.3 0.0012212199999999999 3.3 0.00122132 0 0.00122124 0 0.00122134 3.3 0.0012212599999999998 3.3 0.00122136 0 0.00122128 0 0.00122138 3.3 0.0012212999999999998 3.3 0.0012213999999999999 0 0.00122132 0 0.00122142 3.3 0.00122134 3.3 0.00122144 0 0.00122136 0 0.00122146 3.3 0.00122138 3.3 0.00122148 0 0.0012213999999999999 0 0.0012215 3.3 0.00122142 3.3 0.00122152 0 0.0012214399999999999 0 0.00122154 3.3 0.00122146 3.3 0.00122156 0 0.0012214799999999998 0 0.0012215799999999999 3.3 0.0012215 3.3 0.0012216 0 0.0012215199999999998 0 0.0012216199999999999 3.3 0.00122154 3.3 0.00122164 0 0.00122156 0 0.00122166 3.3 0.0012215799999999999 3.3 0.00122168 0 0.0012216 0 0.0012217 3.3 0.0012216199999999999 3.3 0.00122172 0 0.00122164 0 0.00122174 3.3 0.0012216599999999998 3.3 0.00122176 0 0.00122168 0 0.00122178 3.3 0.0012216999999999998 3.3 0.0012217999999999999 0 0.00122172 0 0.00122182 3.3 0.00122174 3.3 0.00122184 0 0.00122176 0 0.00122186 3.3 0.00122178 3.3 0.00122188 0 0.0012217999999999999 0 0.0012219 3.3 0.00122182 3.3 0.00122192 0 0.0012218399999999999 0 0.00122194 3.3 0.00122186 3.3 0.00122196 0 0.0012218799999999998 0 0.00122198 3.3 0.0012219 3.3 0.001222 0 0.0012219199999999998 0 0.0012220199999999999 3.3 0.00122194 3.3 0.00122204 0 0.00122196 0 0.00122206 3.3 0.00122198 3.3 0.00122208 0 0.001222 0 0.0012221 3.3 0.0012220199999999999 3.3 0.00122212 0 0.00122204 0 0.00122214 3.3 0.0012220599999999999 3.3 0.00122216 0 0.00122208 0 0.00122218 3.3 0.0012220999999999998 3.3 0.0012222 0 0.00122212 0 0.00122222 3.3 0.0012221399999999998 3.3 0.0012222399999999999 0 0.00122216 0 0.00122226 3.3 0.00122218 3.3 0.00122228 0 0.0012222 0 0.0012223 3.3 0.00122222 3.3 0.00122232 0 0.0012222399999999999 0 0.00122234 3.3 0.00122226 3.3 0.00122236 0 0.0012222799999999999 0 0.00122238 3.3 0.0012223 3.3 0.0012224 0 0.0012223199999999998 0 0.0012224199999999999 3.3 0.00122234 3.3 0.00122244 0 0.00122236 0 0.00122246 3.3 0.00122238 3.3 0.00122248 0 0.0012224 0 0.0012225 3.3 0.0012224199999999999 3.3 0.00122252 0 0.00122244 0 0.00122254 3.3 0.0012224599999999999 3.3 0.00122256 0 0.00122248 0 0.00122258 3.3 0.0012224999999999998 3.3 0.0012226 0 0.00122252 0 0.00122262 3.3 0.0012225399999999998 3.3 0.0012226399999999999 0 0.00122256 0 0.00122266 3.3 0.00122258 3.3 0.00122268 0 0.0012226 0 0.0012227 3.3 0.00122262 3.3 0.00122272 0 0.0012226399999999999 0 0.00122274 3.3 0.00122266 3.3 0.00122276 0 0.0012226799999999999 0 0.00122278 3.3 0.0012227 3.3 0.0012228 0 0.0012227199999999998 0 0.00122282 3.3 0.00122274 3.3 0.00122284 0 0.0012227599999999998 0 0.0012228599999999999 3.3 0.00122278 3.3 0.00122288 0 0.0012228 0 0.0012229 3.3 0.00122282 3.3 0.00122292 0 0.00122284 0 0.00122294 3.3 0.0012228599999999999 3.3 0.00122296 0 0.00122288 0 0.00122298 3.3 0.0012228999999999999 3.3 0.001223 0 0.00122292 0 0.00122302 3.3 0.0012229399999999998 3.3 0.0012230399999999999 0 0.00122296 0 0.00122306 3.3 0.0012229799999999998 3.3 0.0012230799999999999 0 0.001223 0 0.0012231 3.3 0.00122302 3.3 0.00122312 0 0.0012230399999999999 0 0.00122314 3.3 0.00122306 3.3 0.00122316 0 0.0012230799999999999 0 0.00122318 3.3 0.0012231 3.3 0.0012232 0 0.0012231199999999998 0 0.00122322 3.3 0.00122314 3.3 0.00122324 0 0.0012231599999999998 0 0.0012232599999999999 3.3 0.00122318 3.3 0.00122328 0 0.0012232 0 0.0012233 3.3 0.00122322 3.3 0.00122332 0 0.00122324 0 0.00122334 3.3 0.0012232599999999999 3.3 0.00122336 0 0.00122328 0 0.00122338 3.3 0.0012232999999999999 3.3 0.0012234 0 0.00122332 0 0.00122342 3.3 0.0012233399999999998 3.3 0.00122344 0 0.00122336 0 0.00122346 3.3 0.0012233799999999998 3.3 0.0012234799999999999 0 0.0012234 0 0.0012235 3.3 0.00122342 3.3 0.00122352 0 0.00122344 0 0.00122354 3.3 0.00122346 3.3 0.00122356 0 0.0012234799999999999 0 0.00122358 3.3 0.0012235 3.3 0.0012236 0 0.0012235199999999999 0 0.00122362 3.3 0.00122354 3.3 0.00122364 0 0.0012235599999999998 0 0.00122366 3.3 0.00122358 3.3 0.00122368 0 0.0012235999999999998 0 0.0012236999999999999 3.3 0.00122362 3.3 0.00122372 0 0.00122364 0 0.00122374 3.3 0.00122366 3.3 0.00122376 0 0.00122368 0 0.00122378 3.3 0.0012236999999999999 3.3 0.0012238 0 0.00122372 0 0.00122382 3.3 0.0012237399999999999 3.3 0.00122384 0 0.00122376 0 0.00122386 3.3 0.0012237799999999998 3.3 0.0012238799999999999 0 0.0012238 0 0.0012239 3.3 0.0012238199999999998 3.3 0.0012239199999999999 0 0.00122384 0 0.00122394 3.3 0.00122386 3.3 0.00122396 0 0.0012238799999999999 0 0.00122398 3.3 0.0012239 3.3 0.001224 0 0.0012239199999999999 0 0.00122402 3.3 0.00122394 3.3 0.00122404 0 0.0012239599999999998 0 0.00122406 3.3 0.00122398 3.3 0.00122408 0 0.0012239999999999998 0 0.0012240999999999999 3.3 0.00122402 3.3 0.00122412 0 0.00122404 0 0.00122414 3.3 0.00122406 3.3 0.00122416 0 0.00122408 0 0.00122418 3.3 0.0012240999999999999 3.3 0.0012242 0 0.00122412 0 0.00122422 3.3 0.0012241399999999999 3.3 0.00122424 0 0.00122416 0 0.00122426 3.3 0.0012241799999999998 3.3 0.00122428 0 0.0012242 0 0.0012243 3.3 0.0012242199999999998 3.3 0.0012243199999999999 0 0.00122424 0 0.00122434 3.3 0.00122426 3.3 0.00122436 0 0.00122428 0 0.00122438 3.3 0.0012243 3.3 0.0012244 0 0.0012243199999999999 0 0.00122442 3.3 0.00122434 3.3 0.00122444 0 0.0012243599999999999 0 0.00122446 3.3 0.00122438 3.3 0.00122448 0 0.0012243999999999998 0 0.0012245 3.3 0.00122442 3.3 0.00122452 0 0.0012244399999999998 0 0.0012245399999999999 3.3 0.00122446 3.3 0.00122456 0 0.00122448 0 0.00122458 3.3 0.0012245 3.3 0.0012246 0 0.00122452 0 0.00122462 3.3 0.0012245399999999999 3.3 0.00122464 0 0.00122456 0 0.00122466 3.3 0.0012245799999999999 3.3 0.00122468 0 0.0012246 0 0.0012247 3.3 0.0012246199999999998 3.3 0.0012247199999999999 0 0.00122464 0 0.00122474 3.3 0.0012246599999999998 3.3 0.0012247599999999999 0 0.00122468 0 0.00122478 3.3 0.0012247 3.3 0.0012248 0 0.0012247199999999999 0 0.00122482 3.3 0.00122474 3.3 0.00122484 0 0.0012247599999999999 0 0.00122486 3.3 0.00122478 3.3 0.00122488 0 0.0012247999999999998 0 0.0012249 3.3 0.00122482 3.3 0.00122492 0 0.0012248399999999998 0 0.0012249399999999999 3.3 0.00122486 3.3 0.00122496 0 0.00122488 0 0.00122498 3.3 0.0012249 3.3 0.001225 0 0.00122492 0 0.00122502 3.3 0.0012249399999999999 3.3 0.00122504 0 0.00122496 0 0.00122506 3.3 0.0012249799999999999 3.3 0.00122508 0 0.001225 0 0.0012251 3.3 0.0012250199999999998 3.3 0.00122512 0 0.00122504 0 0.00122514 3.3 0.0012250599999999998 3.3 0.0012251599999999999 0 0.00122508 0 0.00122518 3.3 0.0012251 3.3 0.0012252 0 0.00122512 0 0.00122522 3.3 0.00122514 3.3 0.00122524 0 0.0012251599999999999 0 0.00122526 3.3 0.00122518 3.3 0.00122528 0 0.0012251999999999999 0 0.0012253 3.3 0.00122522 3.3 0.00122532 0 0.0012252399999999998 0 0.00122534 3.3 0.00122526 3.3 0.00122536 0 0.0012252799999999998 0 0.0012253799999999999 3.3 0.0012253 3.3 0.0012254 0 0.00122532 0 0.00122542 3.3 0.00122534 3.3 0.00122544 0 0.00122536 0 0.00122546 3.3 0.0012253799999999999 3.3 0.00122548 0 0.0012254 0 0.0012255 3.3 0.0012254199999999999 3.3 0.00122552 0 0.00122544 0 0.00122554 3.3 0.0012254599999999998 3.3 0.0012255599999999999 0 0.00122548 0 0.00122558 3.3 0.0012255 3.3 0.0012256 0 0.00122552 0 0.00122562 3.3 0.00122554 3.3 0.00122564 0 0.0012255599999999999 0 0.00122566 3.3 0.00122558 3.3 0.00122568 0 0.0012255999999999999 0 0.0012257 3.3 0.00122562 3.3 0.00122572 0 0.0012256399999999998 0 0.00122574 3.3 0.00122566 3.3 0.00122576 0 0.0012256799999999998 0 0.0012257799999999999 3.3 0.0012257 3.3 0.0012258 0 0.00122572 0 0.00122582 3.3 0.00122574 3.3 0.00122584 0 0.00122576 0 0.00122586 3.3 0.0012257799999999999 3.3 0.00122588 0 0.0012258 0 0.0012259 3.3 0.0012258199999999999 3.3 0.00122592 0 0.00122584 0 0.00122594 3.3 0.0012258599999999998 3.3 0.00122596 0 0.00122588 0 0.00122598 3.3 0.0012258999999999998 3.3 0.0012259999999999999 0 0.00122592 0 0.00122602 3.3 0.00122594 3.3 0.00122604 0 0.00122596 0 0.00122606 3.3 0.00122598 3.3 0.00122608 0 0.0012259999999999999 0 0.0012261 3.3 0.00122602 3.3 0.00122612 0 0.0012260399999999999 0 0.00122614 3.3 0.00122606 3.3 0.00122616 0 0.0012260799999999998 0 0.0012261799999999999 3.3 0.0012261 3.3 0.0012262 0 0.0012261199999999998 0 0.0012262199999999999 3.3 0.00122614 3.3 0.00122624 0 0.00122616 0 0.00122626 3.3 0.0012261799999999999 3.3 0.00122628 0 0.0012262 0 0.0012263 3.3 0.0012262199999999999 3.3 0.00122632 0 0.00122624 0 0.00122634 3.3 0.0012262599999999999 3.3 0.00122636 0 0.00122628 0 0.00122638 3.3 0.0012262999999999998 3.3 0.0012263999999999999 0 0.00122632 0 0.00122642 3.3 0.00122634 3.3 0.00122644 0 0.00122636 0 0.00122646 3.3 0.00122638 3.3 0.00122648 0 0.0012263999999999999 0 0.0012265 3.3 0.00122642 3.3 0.00122652 0 0.0012264399999999999 0 0.00122654 3.3 0.00122646 3.3 0.00122656 0 0.0012264799999999998 0 0.00122658 3.3 0.0012265 3.3 0.0012266 0 0.0012265199999999998 0 0.0012266199999999999 3.3 0.00122654 3.3 0.00122664 0 0.00122656 0 0.00122666 3.3 0.00122658 3.3 0.00122668 0 0.0012266 0 0.0012267 3.3 0.0012266199999999999 3.3 0.00122672 0 0.00122664 0 0.00122674 3.3 0.0012266599999999999 3.3 0.00122676 0 0.00122668 0 0.00122678 3.3 0.0012266999999999998 3.3 0.0012268 0 0.00122672 0 0.00122682 3.3 0.0012267399999999998 3.3 0.0012268399999999999 0 0.00122676 0 0.00122686 3.3 0.00122678 3.3 0.00122688 0 0.0012268 0 0.0012269 3.3 0.00122682 3.3 0.00122692 0 0.0012268399999999999 0 0.00122694 3.3 0.00122686 3.3 0.00122696 0 0.0012268799999999999 0 0.00122698 3.3 0.0012269 3.3 0.001227 0 0.0012269199999999998 0 0.0012270199999999999 3.3 0.00122694 3.3 0.00122704 0 0.0012269599999999998 0 0.0012270599999999999 3.3 0.00122698 3.3 0.00122708 0 0.001227 0 0.0012271 3.3 0.0012270199999999999 3.3 0.00122712 0 0.00122704 0 0.00122714 3.3 0.0012270599999999999 3.3 0.00122716 0 0.00122708 0 0.00122718 3.3 0.0012270999999999998 3.3 0.0012272 0 0.00122712 0 0.00122722 3.3 0.0012271399999999998 3.3 0.0012272399999999999 0 0.00122716 0 0.00122726 3.3 0.00122718 3.3 0.00122728 0 0.0012272 0 0.0012273 3.3 0.00122722 3.3 0.00122732 0 0.0012272399999999999 0 0.00122734 3.3 0.00122726 3.3 0.00122736 0 0.0012272799999999999 0 0.00122738 3.3 0.0012273 3.3 0.0012274 0 0.0012273199999999998 0 0.00122742 3.3 0.00122734 3.3 0.00122744 0 0.0012273599999999998 0 0.0012274599999999999 3.3 0.00122738 3.3 0.00122748 0 0.0012274 0 0.0012275 3.3 0.00122742 3.3 0.00122752 0 0.00122744 0 0.00122754 3.3 0.0012274599999999999 3.3 0.00122756 0 0.00122748 0 0.00122758 3.3 0.0012274999999999999 3.3 0.0012276 0 0.00122752 0 0.00122762 3.3 0.0012275399999999998 3.3 0.00122764 0 0.00122756 0 0.00122766 3.3 0.0012275799999999998 3.3 0.0012276799999999999 0 0.0012276 0 0.0012277 3.3 0.00122762 3.3 0.00122772 0 0.00122764 0 0.00122774 3.3 0.00122766 3.3 0.00122776 0 0.0012276799999999999 0 0.00122778 3.3 0.0012277 3.3 0.0012278 0 0.0012277199999999999 0 0.00122782 3.3 0.00122774 3.3 0.00122784 0 0.0012277599999999998 0 0.0012278599999999999 3.3 0.00122778 3.3 0.00122788 0 0.0012277999999999998 0 0.0012278999999999999 3.3 0.00122782 3.3 0.00122792 0 0.00122784 0 0.00122794 3.3 0.0012278599999999999 3.3 0.00122796 0 0.00122788 0 0.00122798 3.3 0.0012278999999999999 3.3 0.001228 0 0.00122792 0 0.00122802 3.3 0.0012279399999999998 3.3 0.00122804 0 0.00122796 0 0.00122806 3.3 0.0012279799999999998 3.3 0.0012280799999999999 0 0.001228 0 0.0012281 3.3 0.00122802 3.3 0.00122812 0 0.00122804 0 0.00122814 3.3 0.00122806 3.3 0.00122816 0 0.0012280799999999999 0 0.00122818 3.3 0.0012281 3.3 0.0012282 0 0.0012281199999999999 0 0.00122822 3.3 0.00122814 3.3 0.00122824 0 0.0012281599999999998 0 0.00122826 3.3 0.00122818 3.3 0.00122828 0 0.0012281999999999998 0 0.0012282999999999999 3.3 0.00122822 3.3 0.00122832 0 0.00122824 0 0.00122834 3.3 0.00122826 3.3 0.00122836 0 0.00122828 0 0.00122838 3.3 0.0012282999999999999 3.3 0.0012284 0 0.00122832 0 0.00122842 3.3 0.0012283399999999999 3.3 0.00122844 0 0.00122836 0 0.00122846 3.3 0.0012283799999999998 3.3 0.00122848 0 0.0012284 0 0.0012285 3.3 0.0012284199999999998 3.3 0.0012285199999999999 0 0.00122844 0 0.00122854 3.3 0.00122846 3.3 0.00122856 0 0.00122848 0 0.00122858 3.3 0.0012285 3.3 0.0012286 0 0.0012285199999999999 0 0.00122862 3.3 0.00122854 3.3 0.00122864 0 0.0012285599999999999 0 0.00122866 3.3 0.00122858 3.3 0.00122868 0 0.0012285999999999998 0 0.0012286999999999999 3.3 0.00122862 3.3 0.00122872 0 0.0012286399999999998 0 0.0012287399999999999 3.3 0.00122866 3.3 0.00122876 0 0.00122868 0 0.00122878 3.3 0.0012286999999999999 3.3 0.0012288 0 0.00122872 0 0.00122882 3.3 0.0012287399999999999 3.3 0.00122884 0 0.00122876 0 0.00122886 3.3 0.0012287799999999998 3.3 0.00122888 0 0.0012288 0 0.0012289 3.3 0.0012288199999999998 3.3 0.0012289199999999999 0 0.00122884 0 0.00122894 3.3 0.00122886 3.3 0.00122896 0 0.00122888 0 0.00122898 3.3 0.0012289 3.3 0.001229 0 0.0012289199999999999 0 0.00122902 3.3 0.00122894 3.3 0.00122904 0 0.0012289599999999999 0 0.00122906 3.3 0.00122898 3.3 0.00122908 0 0.0012289999999999998 0 0.0012291 3.3 0.00122902 3.3 0.00122912 0 0.0012290399999999998 0 0.0012291399999999999 3.3 0.00122906 3.3 0.00122916 0 0.00122908 0 0.00122918 3.3 0.0012291 3.3 0.0012292 0 0.00122912 0 0.00122922 3.3 0.0012291399999999999 3.3 0.00122924 0 0.00122916 0 0.00122926 3.3 0.0012291799999999999 3.3 0.00122928 0 0.0012292 0 0.0012293 3.3 0.0012292199999999998 3.3 0.00122932 0 0.00122924 0 0.00122934 3.3 0.0012292599999999998 3.3 0.0012293599999999999 0 0.00122928 0 0.00122938 3.3 0.0012293 3.3 0.0012294 0 0.00122932 0 0.00122942 3.3 0.00122934 3.3 0.00122944 0 0.0012293599999999999 0 0.00122946 3.3 0.00122938 3.3 0.00122948 0 0.0012293999999999999 0 0.0012295 3.3 0.00122942 3.3 0.00122952 0 0.0012294399999999998 0 0.0012295399999999999 3.3 0.00122946 3.3 0.00122956 0 0.00122948 0 0.00122958 3.3 0.0012295 3.3 0.0012296 0 0.00122952 0 0.00122962 3.3 0.0012295399999999999 3.3 0.00122964 0 0.00122956 0 0.00122966 3.3 0.0012295799999999999 3.3 0.00122968 0 0.0012296 0 0.0012297 3.3 0.0012296199999999998 3.3 0.00122972 0 0.00122964 0 0.00122974 3.3 0.0012296599999999998 3.3 0.0012297599999999999 0 0.00122968 0 0.00122978 3.3 0.0012297 3.3 0.0012298 0 0.00122972 0 0.00122982 3.3 0.00122974 3.3 0.00122984 0 0.0012297599999999999 0 0.00122986 3.3 0.00122978 3.3 0.00122988 0 0.0012297999999999999 0 0.0012299 3.3 0.00122982 3.3 0.00122992 0 0.0012298399999999998 0 0.00122994 3.3 0.00122986 3.3 0.00122996 0 0.0012298799999999998 0 0.0012299799999999999 3.3 0.0012299 3.3 0.00123 0 0.00122992 0 0.00123002 3.3 0.00122994 3.3 0.00123004 0 0.00122996 0 0.00123006 3.3 0.0012299799999999999 3.3 0.00123008 0 0.00123 0 0.0012301 3.3 0.0012300199999999999 3.3 0.00123012 0 0.00123004 0 0.00123014 3.3 0.0012300599999999998 3.3 0.0012301599999999999 0 0.00123008 0 0.00123018 3.3 0.0012300999999999998 3.3 0.0012301999999999999 0 0.00123012 0 0.00123022 3.3 0.00123014 3.3 0.00123024 0 0.0012301599999999999 0 0.00123026 3.3 0.00123018 3.3 0.00123028 0 0.0012301999999999999 0 0.0012303 3.3 0.00123022 3.3 0.00123032 0 0.0012302399999999998 0 0.00123034 3.3 0.00123026 3.3 0.00123036 0 0.0012302799999999998 0 0.0012303799999999999 3.3 0.0012303 3.3 0.0012304 0 0.00123032 0 0.00123042 3.3 0.00123034 3.3 0.00123044 0 0.00123036 0 0.00123046 3.3 0.0012303799999999999 3.3 0.00123048 0 0.0012304 0 0.0012305 3.3 0.0012304199999999999 3.3 0.00123052 0 0.00123044 0 0.00123054 3.3 0.0012304599999999998 3.3 0.00123056 0 0.00123048 0 0.00123058 3.3 0.0012304999999999998 3.3 0.0012305999999999999 0 0.00123052 0 0.00123062 3.3 0.00123054 3.3 0.00123064 0 0.00123056 0 0.00123066 3.3 0.00123058 3.3 0.00123068 0 0.0012305999999999999 0 0.0012307 3.3 0.00123062 3.3 0.00123072 0 0.0012306399999999999 0 0.00123074 3.3 0.00123066 3.3 0.00123076 0 0.0012306799999999998 0 0.00123078 3.3 0.0012307 3.3 0.0012308 0 0.0012307199999999998 0 0.0012308199999999999 3.3 0.00123074 3.3 0.00123084 0 0.00123076 0 0.00123086 3.3 0.00123078 3.3 0.00123088 0 0.0012308 0 0.0012309 3.3 0.0012308199999999999 3.3 0.00123092 0 0.00123084 0 0.00123094 3.3 0.0012308599999999999 3.3 0.00123096 0 0.00123088 0 0.00123098 3.3 0.0012308999999999998 3.3 0.0012309999999999999 0 0.00123092 0 0.00123102 3.3 0.0012309399999999998 3.3 0.0012310399999999999 0 0.00123096 0 0.00123106 3.3 0.00123098 3.3 0.00123108 0 0.0012309999999999999 0 0.0012311 3.3 0.00123102 3.3 0.00123112 0 0.0012310399999999999 0 0.00123114 3.3 0.00123106 3.3 0.00123116 0 0.0012310799999999998 0 0.00123118 3.3 0.0012311 3.3 0.0012312 0 0.0012311199999999998 0 0.0012312199999999999 3.3 0.00123114 3.3 0.00123124 0 0.00123116 0 0.00123126 3.3 0.00123118 3.3 0.00123128 0 0.0012312 0 0.0012313 3.3 0.0012312199999999999 3.3 0.00123132 0 0.00123124 0 0.00123134 3.3 0.0012312599999999999 3.3 0.00123136 0 0.00123128 0 0.00123138 3.3 0.0012312999999999998 3.3 0.0012314 0 0.00123132 0 0.00123142 3.3 0.0012313399999999998 3.3 0.0012314399999999999 0 0.00123136 0 0.00123146 3.3 0.00123138 3.3 0.00123148 0 0.0012314 0 0.0012315 3.3 0.00123142 3.3 0.00123152 0 0.0012314399999999999 0 0.00123154 3.3 0.00123146 3.3 0.00123156 0 0.0012314799999999999 0 0.00123158 3.3 0.0012315 3.3 0.0012316 0 0.0012315199999999998 0 0.00123162 3.3 0.00123154 3.3 0.00123164 0 0.0012315599999999998 0 0.0012316599999999999 3.3 0.00123158 3.3 0.00123168 0 0.0012316 0 0.0012317 3.3 0.00123162 3.3 0.00123172 0 0.00123164 0 0.00123174 3.3 0.0012316599999999999 3.3 0.00123176 0 0.00123168 0 0.00123178 3.3 0.0012316999999999999 3.3 0.0012318 0 0.00123172 0 0.00123182 3.3 0.0012317399999999998 3.3 0.0012318399999999999 0 0.00123176 0 0.00123186 3.3 0.0012317799999999998 3.3 0.0012318799999999999 0 0.0012318 0 0.0012319 3.3 0.00123182 3.3 0.00123192 0 0.0012318399999999999 0 0.00123194 3.3 0.00123186 3.3 0.00123196 0 0.0012318799999999999 0 0.00123198 3.3 0.0012319 3.3 0.001232 0 0.0012319199999999998 0 0.00123202 3.3 0.00123194 3.3 0.00123204 0 0.0012319599999999998 0 0.0012320599999999999 3.3 0.00123198 3.3 0.00123208 0 0.001232 0 0.0012321 3.3 0.00123202 3.3 0.00123212 0 0.00123204 0 0.00123214 3.3 0.0012320599999999999 3.3 0.00123216 0 0.00123208 0 0.00123218 3.3 0.0012320999999999999 3.3 0.0012322 0 0.00123212 0 0.00123222 3.3 0.0012321399999999998 3.3 0.00123224 0 0.00123216 0 0.00123226 3.3 0.0012321799999999998 3.3 0.0012322799999999999 0 0.0012322 0 0.0012323 3.3 0.00123222 3.3 0.00123232 0 0.00123224 0 0.00123234 3.3 0.00123226 3.3 0.00123236 0 0.0012322799999999999 0 0.00123238 3.3 0.0012323 3.3 0.0012324 0 0.0012323199999999999 0 0.00123242 3.3 0.00123234 3.3 0.00123244 0 0.0012323599999999998 0 0.00123246 3.3 0.00123238 3.3 0.00123248 0 0.0012323999999999998 0 0.0012324999999999999 3.3 0.00123242 3.3 0.00123252 0 0.00123244 0 0.00123254 3.3 0.00123246 3.3 0.00123256 0 0.00123248 0 0.00123258 3.3 0.0012324999999999999 3.3 0.0012326 0 0.00123252 0 0.00123262 3.3 0.0012325399999999999 3.3 0.00123264 0 0.00123256 0 0.00123266 3.3 0.0012325799999999998 3.3 0.0012326799999999999 0 0.0012326 0 0.0012327 3.3 0.00123262 3.3 0.00123272 0 0.00123264 0 0.00123274 3.3 0.00123266 3.3 0.00123276 0 0.0012326799999999999 0 0.00123278 3.3 0.0012327 3.3 0.0012328 0 0.0012327199999999999 0 0.00123282 3.3 0.00123274 3.3 0.00123284 0 0.0012327599999999998 0 0.00123286 3.3 0.00123278 3.3 0.00123288 0 0.0012327999999999998 0 0.0012328999999999999 3.3 0.00123282 3.3 0.00123292 0 0.00123284 0 0.00123294 3.3 0.00123286 3.3 0.00123296 0 0.00123288 0 0.00123298 3.3 0.0012328999999999999 3.3 0.001233 0 0.00123292 0 0.00123302 3.3 0.0012329399999999999 3.3 0.00123304 0 0.00123296 0 0.00123306 3.3 0.0012329799999999998 3.3 0.00123308 0 0.001233 0 0.0012331 3.3 0.0012330199999999998 3.3 0.0012331199999999999 0 0.00123304 0 0.00123314 3.3 0.00123306 3.3 0.00123316 0 0.00123308 0 0.00123318 3.3 0.0012331 3.3 0.0012332 0 0.0012331199999999999 0 0.00123322 3.3 0.00123314 3.3 0.00123324 0 0.0012331599999999999 0 0.00123326 3.3 0.00123318 3.3 0.00123328 0 0.0012331999999999998 0 0.0012332999999999999 3.3 0.00123322 3.3 0.00123332 0 0.0012332399999999998 0 0.0012333399999999999 3.3 0.00123326 3.3 0.00123336 0 0.00123328 0 0.00123338 3.3 0.0012332999999999999 3.3 0.0012334 0 0.00123332 0 0.00123342 3.3 0.0012333399999999999 3.3 0.00123344 0 0.00123336 0 0.00123346 3.3 0.0012333799999999998 3.3 0.00123348 0 0.0012334 0 0.0012335 3.3 0.0012334199999999998 3.3 0.0012335199999999999 0 0.00123344 0 0.00123354 3.3 0.00123346 3.3 0.00123356 0 0.00123348 0 0.00123358 3.3 0.0012335 3.3 0.0012336 0 0.0012335199999999999 0 0.00123362 3.3 0.00123354 3.3 0.00123364 0 0.0012335599999999999 0 0.00123366 3.3 0.00123358 3.3 0.00123368 0 0.0012335999999999998 0 0.0012337 3.3 0.00123362 3.3 0.00123372 0 0.0012336399999999998 0 0.0012337399999999999 3.3 0.00123366 3.3 0.00123376 0 0.00123368 0 0.00123378 3.3 0.0012337 3.3 0.0012338 0 0.00123372 0 0.00123382 3.3 0.0012337399999999999 3.3 0.00123384 0 0.00123376 0 0.00123386 3.3 0.0012337799999999999 3.3 0.00123388 0 0.0012338 0 0.0012339 3.3 0.0012338199999999998 3.3 0.00123392 0 0.00123384 0 0.00123394 3.3 0.0012338599999999998 3.3 0.0012339599999999999 0 0.00123388 0 0.00123398 3.3 0.0012339 3.3 0.001234 0 0.00123392 0 0.00123402 3.3 0.00123394 3.3 0.00123404 0 0.0012339599999999999 0 0.00123406 3.3 0.00123398 3.3 0.00123408 0 0.0012339999999999999 0 0.0012341 3.3 0.00123402 3.3 0.00123412 0 0.0012340399999999998 0 0.0012341399999999999 3.3 0.00123406 3.3 0.00123416 0 0.0012340799999999998 0 0.0012341799999999999 3.3 0.0012341 3.3 0.0012342 0 0.00123412 0 0.00123422 3.3 0.0012341399999999999 3.3 0.00123424 0 0.00123416 0 0.00123426 3.3 0.0012341799999999999 3.3 0.00123428 0 0.0012342 0 0.0012343 3.3 0.0012342199999999998 3.3 0.00123432 0 0.00123424 0 0.00123434 3.3 0.0012342599999999998 3.3 0.0012343599999999999 0 0.00123428 0 0.00123438 3.3 0.0012343 3.3 0.0012344 0 0.00123432 0 0.00123442 3.3 0.00123434 3.3 0.00123444 0 0.0012343599999999999 0 0.00123446 3.3 0.00123438 3.3 0.00123448 0 0.0012343999999999999 0 0.0012345 3.3 0.00123442 3.3 0.00123452 0 0.0012344399999999998 0 0.00123454 3.3 0.00123446 3.3 0.00123456 0 0.0012344799999999998 0 0.0012345799999999999 3.3 0.0012345 3.3 0.0012346 0 0.00123452 0 0.00123462 3.3 0.00123454 3.3 0.00123464 0 0.00123456 0 0.00123466 3.3 0.0012345799999999999 3.3 0.00123468 0 0.0012346 0 0.0012347 3.3 0.0012346199999999999 3.3 0.00123472 0 0.00123464 0 0.00123474 3.3 0.0012346599999999998 3.3 0.00123476 0 0.00123468 0 0.00123478 3.3 0.0012346999999999998 3.3 0.0012347999999999999 0 0.00123472 0 0.00123482 3.3 0.00123474 3.3 0.00123484 0 0.00123476 0 0.00123486 3.3 0.00123478 3.3 0.00123488 0 0.0012347999999999999 0 0.0012349 3.3 0.00123482 3.3 0.00123492 0 0.0012348399999999999 0 0.00123494 3.3 0.00123486 3.3 0.00123496 0 0.0012348799999999998 0 0.0012349799999999999 3.3 0.0012349 3.3 0.001235 0 0.0012349199999999998 0 0.0012350199999999999 3.3 0.00123494 3.3 0.00123504 0 0.00123496 0 0.00123506 3.3 0.0012349799999999999 3.3 0.00123508 0 0.001235 0 0.0012351 3.3 0.0012350199999999999 3.3 0.00123512 0 0.00123504 0 0.00123514 3.3 0.0012350599999999998 3.3 0.00123516 0 0.00123508 0 0.00123518 3.3 0.0012350999999999998 3.3 0.0012351999999999999 0 0.00123512 0 0.00123522 3.3 0.00123514 3.3 0.00123524 0 0.00123516 0 0.00123526 3.3 0.00123518 3.3 0.00123528 0 0.0012351999999999999 0 0.0012353 3.3 0.00123522 3.3 0.00123532 0 0.0012352399999999999 0 0.00123534 3.3 0.00123526 3.3 0.00123536 0 0.0012352799999999998 0 0.00123538 3.3 0.0012353 3.3 0.0012354 0 0.0012353199999999998 0 0.0012354199999999999 3.3 0.00123534 3.3 0.00123544 0 0.00123536 0 0.00123546 3.3 0.00123538 3.3 0.00123548 0 0.0012354 0 0.0012355 3.3 0.0012354199999999999 3.3 0.00123552 0 0.00123544 0 0.00123554 3.3 0.0012354599999999999 3.3 0.00123556 0 0.00123548 0 0.00123558 3.3 0.0012354999999999998 3.3 0.0012356 0 0.00123552 0 0.00123562 3.3 0.0012355399999999998 3.3 0.0012356399999999999 0 0.00123556 0 0.00123566 3.3 0.00123558 3.3 0.00123568 0 0.0012356 0 0.0012357 3.3 0.00123562 3.3 0.00123572 0 0.0012356399999999999 0 0.00123574 3.3 0.00123566 3.3 0.00123576 0 0.0012356799999999999 0 0.00123578 3.3 0.0012357 3.3 0.0012358 0 0.0012357199999999998 0 0.0012358199999999999 3.3 0.00123574 3.3 0.00123584 0 0.00123576 0 0.00123586 3.3 0.00123578 3.3 0.00123588 0 0.0012358 0 0.0012359 3.3 0.0012358199999999999 3.3 0.00123592 0 0.00123584 0 0.00123594 3.3 0.0012358599999999999 3.3 0.00123596 0 0.00123588 0 0.00123598 3.3 0.0012358999999999998 3.3 0.001236 0 0.00123592 0 0.00123602 3.3 0.0012359399999999998 3.3 0.0012360399999999999 0 0.00123596 0 0.00123606 3.3 0.00123598 3.3 0.00123608 0 0.001236 0 0.0012361 3.3 0.00123602 3.3 0.00123612 0 0.0012360399999999999 0 0.00123614 3.3 0.00123606 3.3 0.00123616 0 0.0012360799999999999 0 0.00123618 3.3 0.0012361 3.3 0.0012362 0 0.0012361199999999998 0 0.00123622 3.3 0.00123614 3.3 0.00123624 0 0.0012361599999999998 0 0.0012362599999999999 3.3 0.00123618 3.3 0.00123628 0 0.0012362 0 0.0012363 3.3 0.00123622 3.3 0.00123632 0 0.00123624 0 0.00123634 3.3 0.0012362599999999999 3.3 0.00123636 0 0.00123628 0 0.00123638 3.3 0.0012362999999999999 3.3 0.0012364 0 0.00123632 0 0.00123642 3.3 0.0012363399999999998 3.3 0.0012364399999999999 0 0.00123636 0 0.00123646 3.3 0.0012363799999999998 3.3 0.0012364799999999999 0 0.0012364 0 0.0012365 3.3 0.00123642 3.3 0.00123652 0 0.0012364399999999999 0 0.00123654 3.3 0.00123646 3.3 0.00123656 0 0.0012364799999999999 0 0.00123658 3.3 0.0012365 3.3 0.0012366 0 0.0012365199999999999 0 0.00123662 3.3 0.00123654 3.3 0.00123664 0 0.0012365599999999998 0 0.0012366599999999999 3.3 0.00123658 3.3 0.00123668 0 0.0012366 0 0.0012367 3.3 0.00123662 3.3 0.00123672 0 0.00123664 0 0.00123674 3.3 0.0012366599999999999 3.3 0.00123676 0 0.00123668 0 0.00123678 3.3 0.0012366999999999999 3.3 0.0012368 0 0.00123672 0 0.00123682 3.3 0.0012367399999999998 3.3 0.00123684 0 0.00123676 0 0.00123686 3.3 0.0012367799999999998 3.3 0.0012368799999999999 0 0.0012368 0 0.0012369 3.3 0.00123682 3.3 0.00123692 0 0.00123684 0 0.00123694 3.3 0.00123686 3.3 0.00123696 0 0.0012368799999999999 0 0.00123698 3.3 0.0012369 3.3 0.001237 0 0.0012369199999999999 0 0.00123702 3.3 0.00123694 3.3 0.00123704 0 0.0012369599999999998 0 0.00123706 3.3 0.00123698 3.3 0.00123708 0 0.0012369999999999998 0 0.0012370999999999999 3.3 0.00123702 3.3 0.00123712 0 0.00123704 0 0.00123714 3.3 0.00123706 3.3 0.00123716 0 0.00123708 0 0.00123718 3.3 0.0012370999999999999 3.3 0.0012372 0 0.00123712 0 0.00123722 3.3 0.0012371399999999999 3.3 0.00123724 0 0.00123716 0 0.00123726 3.3 0.0012371799999999998 3.3 0.0012372799999999999 0 0.0012372 0 0.0012373 3.3 0.0012372199999999998 3.3 0.0012373199999999999 0 0.00123724 0 0.00123734 3.3 0.00123726 3.3 0.00123736 0 0.0012372799999999999 0 0.00123738 3.3 0.0012373 3.3 0.0012374 0 0.0012373199999999999 0 0.00123742 3.3 0.00123734 3.3 0.00123744 0 0.0012373599999999998 0 0.00123746 3.3 0.00123738 3.3 0.00123748 0 0.0012373999999999998 0 0.0012374999999999999 3.3 0.00123742 3.3 0.00123752 0 0.00123744 0 0.00123754 3.3 0.00123746 3.3 0.00123756 0 0.00123748 0 0.00123758 3.3 0.0012374999999999999 3.3 0.0012376 0 0.00123752 0 0.00123762 3.3 0.0012375399999999999 3.3 0.00123764 0 0.00123756 0 0.00123766 3.3 0.0012375799999999998 3.3 0.00123768 0 0.0012376 0 0.0012377 3.3 0.0012376199999999998 3.3 0.0012377199999999999 0 0.00123764 0 0.00123774 3.3 0.00123766 3.3 0.00123776 0 0.00123768 0 0.00123778 3.3 0.0012377 3.3 0.0012378 0 0.0012377199999999999 0 0.00123782 3.3 0.00123774 3.3 0.00123784 0 0.0012377599999999999 0 0.00123786 3.3 0.00123778 3.3 0.00123788 0 0.0012377999999999998 0 0.0012379 3.3 0.00123782 3.3 0.00123792 0 0.0012378399999999998 0 0.0012379399999999999 3.3 0.00123786 3.3 0.00123796 0 0.00123788 0 0.00123798 3.3 0.0012379 3.3 0.001238 0 0.00123792 0 0.00123802 3.3 0.0012379399999999999 3.3 0.00123804 0 0.00123796 0 0.00123806 3.3 0.0012379799999999999 3.3 0.00123808 0 0.001238 0 0.0012381 3.3 0.0012380199999999998 3.3 0.0012381199999999999 0 0.00123804 0 0.00123814 3.3 0.0012380599999999998 3.3 0.0012381599999999999 0 0.00123808 0 0.00123818 3.3 0.0012381 3.3 0.0012382 0 0.0012381199999999999 0 0.00123822 3.3 0.00123814 3.3 0.00123824 0 0.0012381599999999999 0 0.00123826 3.3 0.00123818 3.3 0.00123828 0 0.0012381999999999998 0 0.0012383 3.3 0.00123822 3.3 0.00123832 0 0.0012382399999999998 0 0.0012383399999999999 3.3 0.00123826 3.3 0.00123836 0 0.00123828 0 0.00123838 3.3 0.0012383 3.3 0.0012384 0 0.00123832 0 0.00123842 3.3 0.0012383399999999999 3.3 0.00123844 0 0.00123836 0 0.00123846 3.3 0.0012383799999999999 3.3 0.00123848 0 0.0012384 0 0.0012385 3.3 0.0012384199999999998 3.3 0.00123852 0 0.00123844 0 0.00123854 3.3 0.0012384599999999998 3.3 0.0012385599999999999 0 0.00123848 0 0.00123858 3.3 0.0012385 3.3 0.0012386 0 0.00123852 0 0.00123862 3.3 0.00123854 3.3 0.00123864 0 0.0012385599999999999 0 0.00123866 3.3 0.00123858 3.3 0.00123868 0 0.0012385999999999999 0 0.0012387 3.3 0.00123862 3.3 0.00123872 0 0.0012386399999999998 0 0.00123874 3.3 0.00123866 3.3 0.00123876 0 0.0012386799999999998 0 0.0012387799999999999 3.3 0.0012387 3.3 0.0012388 0 0.00123872 0 0.00123882 3.3 0.00123874 3.3 0.00123884 0 0.00123876 0 0.00123886 3.3 0.0012387799999999999 3.3 0.00123888 0 0.0012388 0 0.0012389 3.3 0.0012388199999999999 3.3 0.00123892 0 0.00123884 0 0.00123894 3.3 0.0012388599999999998 3.3 0.0012389599999999999 0 0.00123888 0 0.00123898 3.3 0.0012388999999999998 3.3 0.0012389999999999999 0 0.00123892 0 0.00123902 3.3 0.00123894 3.3 0.00123904 0 0.0012389599999999999 0 0.00123906 3.3 0.00123898 3.3 0.00123908 0 0.0012389999999999999 0 0.0012391 3.3 0.00123902 3.3 0.00123912 0 0.0012390399999999998 0 0.00123914 3.3 0.00123906 3.3 0.00123916 0 0.0012390799999999998 0 0.0012391799999999999 3.3 0.0012391 3.3 0.0012392 0 0.00123912 0 0.00123922 3.3 0.00123914 3.3 0.00123924 0 0.00123916 0 0.00123926 3.3 0.0012391799999999999 3.3 0.00123928 0 0.0012392 0 0.0012393 3.3 0.0012392199999999999 3.3 0.00123932 0 0.00123924 0 0.00123934 3.3 0.0012392599999999998 3.3 0.00123936 0 0.00123928 0 0.00123938 3.3 0.0012392999999999998 3.3 0.0012393999999999999 0 0.00123932 0 0.00123942 3.3 0.00123934 3.3 0.00123944 0 0.00123936 0 0.00123946 3.3 0.00123938 3.3 0.00123948 0 0.0012393999999999999 0 0.0012395 3.3 0.00123942 3.3 0.00123952 0 0.0012394399999999999 0 0.00123954 3.3 0.00123946 3.3 0.00123956 0 0.0012394799999999998 0 0.00123958 3.3 0.0012395 3.3 0.0012396 0 0.0012395199999999998 0 0.0012396199999999999 3.3 0.00123954 3.3 0.00123964 0 0.00123956 0 0.00123966 3.3 0.00123958 3.3 0.00123968 0 0.0012396 0 0.0012397 3.3 0.0012396199999999999 3.3 0.00123972 0 0.00123964 0 0.00123974 3.3 0.0012396599999999999 3.3 0.00123976 0 0.00123968 0 0.00123978 3.3 0.0012396999999999998 3.3 0.0012397999999999999 0 0.00123972 0 0.00123982 3.3 0.00123974 3.3 0.00123984 0 0.00123976 0 0.00123986 3.3 0.00123978 3.3 0.00123988 0 0.0012397999999999999 0 0.0012399 3.3 0.00123982 3.3 0.00123992 0 0.0012398399999999999 0 0.00123994 3.3 0.00123986 3.3 0.00123996 0 0.0012398799999999998 0 0.00123998 3.3 0.0012399 3.3 0.00124 0 0.0012399199999999998 0 0.0012400199999999999 3.3 0.00123994 3.3 0.00124004 0 0.00123996 0 0.00124006 3.3 0.00123998 3.3 0.00124008 0 0.00124 0 0.0012401 3.3 0.0012400199999999999 3.3 0.00124012 0 0.00124004 0 0.00124014 3.3 0.0012400599999999999 3.3 0.00124016 0 0.00124008 0 0.00124018 3.3 0.0012400999999999998 3.3 0.0012402 0 0.00124012 0 0.00124022 3.3 0.0012401399999999998 3.3 0.0012402399999999999 0 0.00124016 0 0.00124026 3.3 0.00124018 3.3 0.00124028 0 0.0012402 0 0.0012403 3.3 0.00124022 3.3 0.00124032 0 0.0012402399999999999 0 0.00124034 3.3 0.00124026 3.3 0.00124036 0 0.0012402799999999999 0 0.00124038 3.3 0.0012403 3.3 0.0012404 0 0.0012403199999999998 0 0.0012404199999999999 3.3 0.00124034 3.3 0.00124044 0 0.0012403599999999998 0 0.0012404599999999999 3.3 0.00124038 3.3 0.00124048 0 0.0012404 0 0.0012405 3.3 0.0012404199999999999 3.3 0.00124052 0 0.00124044 0 0.00124054 3.3 0.0012404599999999999 3.3 0.00124056 0 0.00124048 0 0.00124058 3.3 0.0012404999999999998 3.3 0.0012406 0 0.00124052 0 0.00124062 3.3 0.0012405399999999998 3.3 0.0012406399999999999 0 0.00124056 0 0.00124066 3.3 0.00124058 3.3 0.00124068 0 0.0012406 0 0.0012407 3.3 0.00124062 3.3 0.00124072 0 0.0012406399999999999 0 0.00124074 3.3 0.00124066 3.3 0.00124076 0 0.0012406799999999999 0 0.00124078 3.3 0.0012407 3.3 0.0012408 0 0.0012407199999999998 0 0.00124082 3.3 0.00124074 3.3 0.00124084 0 0.0012407599999999998 0 0.0012408599999999999 3.3 0.00124078 3.3 0.00124088 0 0.0012408 0 0.0012409 3.3 0.00124082 3.3 0.00124092 0 0.00124084 0 0.00124094 3.3 0.0012408599999999999 3.3 0.00124096 0 0.00124088 0 0.00124098 3.3 0.0012408999999999999 3.3 0.001241 0 0.00124092 0 0.00124102 3.3 0.0012409399999999998 3.3 0.00124104 0 0.00124096 0 0.00124106 3.3 0.0012409799999999998 3.3 0.0012410799999999999 0 0.001241 0 0.0012411 3.3 0.00124102 3.3 0.00124112 0 0.00124104 0 0.00124114 3.3 0.00124106 3.3 0.00124116 0 0.0012410799999999999 0 0.00124118 3.3 0.0012411 3.3 0.0012412 0 0.0012411199999999999 0 0.00124122 3.3 0.00124114 3.3 0.00124124 0 0.0012411599999999998 0 0.0012412599999999999 3.3 0.00124118 3.3 0.00124128 0 0.0012411999999999998 0 0.0012412999999999999 3.3 0.00124122 3.3 0.00124132 0 0.00124124 0 0.00124134 3.3 0.0012412599999999999 3.3 0.00124136 0 0.00124128 0 0.00124138 3.3 0.0012412999999999999 3.3 0.0012414 0 0.00124132 0 0.00124142 3.3 0.0012413399999999998 3.3 0.00124144 0 0.00124136 0 0.00124146 3.3 0.0012413799999999998 3.3 0.0012414799999999999 0 0.0012414 0 0.0012415 3.3 0.00124142 3.3 0.00124152 0 0.00124144 0 0.00124154 3.3 0.00124146 3.3 0.00124156 0 0.0012414799999999999 0 0.00124158 3.3 0.0012415 3.3 0.0012416 0 0.0012415199999999999 0 0.00124162 3.3 0.00124154 3.3 0.00124164 0 0.0012415599999999998 0 0.00124166 3.3 0.00124158 3.3 0.00124168 0 0.0012415999999999998 0 0.0012416999999999999 3.3 0.00124162 3.3 0.00124172 0 0.00124164 0 0.00124174 3.3 0.00124166 3.3 0.00124176 0 0.00124168 0 0.00124178 3.3 0.0012416999999999999 3.3 0.0012418 0 0.00124172 0 0.00124182 3.3 0.0012417399999999999 3.3 0.00124184 0 0.00124176 0 0.00124186 3.3 0.0012417799999999998 3.3 0.00124188 0 0.0012418 0 0.0012419 3.3 0.0012418199999999998 3.3 0.0012419199999999999 0 0.00124184 0 0.00124194 3.3 0.00124186 3.3 0.00124196 0 0.00124188 0 0.00124198 3.3 0.0012419 3.3 0.001242 0 0.0012419199999999999 0 0.00124202 3.3 0.00124194 3.3 0.00124204 0 0.0012419599999999999 0 0.00124206 3.3 0.00124198 3.3 0.00124208 0 0.0012419999999999998 0 0.0012420999999999999 3.3 0.00124202 3.3 0.00124212 0 0.0012420399999999998 0 0.0012421399999999999 3.3 0.00124206 3.3 0.00124216 0 0.00124208 0 0.00124218 3.3 0.0012420999999999999 3.3 0.0012422 0 0.00124212 0 0.00124222 3.3 0.0012421399999999999 3.3 0.00124224 0 0.00124216 0 0.00124226 3.3 0.0012421799999999998 3.3 0.00124228 0 0.0012422 0 0.0012423 3.3 0.0012422199999999998 3.3 0.0012423199999999999 0 0.00124224 0 0.00124234 3.3 0.00124226 3.3 0.00124236 0 0.00124228 0 0.00124238 3.3 0.0012423 3.3 0.0012424 0 0.0012423199999999999 0 0.00124242 3.3 0.00124234 3.3 0.00124244 0 0.0012423599999999999 0 0.00124246 3.3 0.00124238 3.3 0.00124248 0 0.0012423999999999998 0 0.0012425 3.3 0.00124242 3.3 0.00124252 0 0.0012424399999999998 0 0.0012425399999999999 3.3 0.00124246 3.3 0.00124256 0 0.00124248 0 0.00124258 3.3 0.0012425 3.3 0.0012426 0 0.00124252 0 0.00124262 3.3 0.0012425399999999999 3.3 0.00124264 0 0.00124256 0 0.00124266 3.3 0.0012425799999999999 3.3 0.00124268 0 0.0012426 0 0.0012427 3.3 0.0012426199999999998 3.3 0.00124272 0 0.00124264 0 0.00124274 3.3 0.0012426599999999998 3.3 0.0012427599999999999 0 0.00124268 0 0.00124278 3.3 0.0012427 3.3 0.0012428 0 0.00124272 0 0.00124282 3.3 0.00124274 3.3 0.00124284 0 0.0012427599999999999 0 0.00124286 3.3 0.00124278 3.3 0.00124288 0 0.0012427999999999999 0 0.0012429 3.3 0.00124282 3.3 0.00124292 0 0.0012428399999999998 0 0.0012429399999999999 3.3 0.00124286 3.3 0.00124296 0 0.00124288 0 0.00124298 3.3 0.0012429 3.3 0.001243 0 0.00124292 0 0.00124302 3.3 0.0012429399999999999 3.3 0.00124304 0 0.00124296 0 0.00124306 3.3 0.0012429799999999999 3.3 0.00124308 0 0.001243 0 0.0012431 3.3 0.0012430199999999998 3.3 0.00124312 0 0.00124304 0 0.00124314 3.3 0.0012430599999999998 3.3 0.0012431599999999999 0 0.00124308 0 0.00124318 3.3 0.0012431 3.3 0.0012432 0 0.00124312 0 0.00124322 3.3 0.00124314 3.3 0.00124324 0 0.0012431599999999999 0 0.00124326 3.3 0.00124318 3.3 0.00124328 0 0.0012431999999999999 0 0.0012433 3.3 0.00124322 3.3 0.00124332 0 0.0012432399999999998 0 0.00124334 3.3 0.00124326 3.3 0.00124336 0 0.0012432799999999998 0 0.0012433799999999999 3.3 0.0012433 3.3 0.0012434 0 0.00124332 0 0.00124342 3.3 0.00124334 3.3 0.00124344 0 0.00124336 0 0.00124346 3.3 0.0012433799999999999 3.3 0.00124348 0 0.0012434 0 0.0012435 3.3 0.0012434199999999999 3.3 0.00124352 0 0.00124344 0 0.00124354 3.3 0.0012434599999999998 3.3 0.0012435599999999999 0 0.00124348 0 0.00124358 3.3 0.0012434999999999998 3.3 0.0012435999999999999 0 0.00124352 0 0.00124362 3.3 0.00124354 3.3 0.00124364 0 0.0012435599999999999 0 0.00124366 3.3 0.00124358 3.3 0.00124368 0 0.0012435999999999999 0 0.0012437 3.3 0.00124362 3.3 0.00124372 0 0.0012436399999999998 0 0.00124374 3.3 0.00124366 3.3 0.00124376 0 0.0012436799999999998 0 0.0012437799999999999 3.3 0.0012437 3.3 0.0012438 0 0.00124372 0 0.00124382 3.3 0.00124374 3.3 0.00124384 0 0.00124376 0 0.00124386 3.3 0.0012437799999999999 3.3 0.00124388 0 0.0012438 0 0.0012439 3.3 0.0012438199999999999 3.3 0.00124392 0 0.00124384 0 0.00124394 3.3 0.0012438599999999998 3.3 0.00124396 0 0.00124388 0 0.00124398 3.3 0.0012438999999999998 3.3 0.0012439999999999999 0 0.00124392 0 0.00124402 3.3 0.00124394 3.3 0.00124404 0 0.00124396 0 0.00124406 3.3 0.00124398 3.3 0.00124408 0 0.0012439999999999999 0 0.0012441 3.3 0.00124402 3.3 0.00124412 0 0.0012440399999999999 0 0.00124414 3.3 0.00124406 3.3 0.00124416 0 0.0012440799999999998 0 0.00124418 3.3 0.0012441 3.3 0.0012442 0 0.0012441199999999998 0 0.0012442199999999999 3.3 0.00124414 3.3 0.00124424 0 0.00124416 0 0.00124426 3.3 0.00124418 3.3 0.00124428 0 0.0012442 0 0.0012443 3.3 0.0012442199999999999 3.3 0.00124432 0 0.00124424 0 0.00124434 3.3 0.0012442599999999999 3.3 0.00124436 0 0.00124428 0 0.00124438 3.3 0.0012442999999999998 3.3 0.0012443999999999999 0 0.00124432 0 0.00124442 3.3 0.0012443399999999998 3.3 0.0012444399999999999 0 0.00124436 0 0.00124446 3.3 0.00124438 3.3 0.00124448 0 0.0012443999999999999 0 0.0012445 3.3 0.00124442 3.3 0.00124452 0 0.0012444399999999999 0 0.00124454 3.3 0.00124446 3.3 0.00124456 0 0.0012444799999999998 0 0.00124458 3.3 0.0012445 3.3 0.0012446 0 0.0012445199999999998 0 0.0012446199999999999 3.3 0.00124454 3.3 0.00124464 0 0.00124456 0 0.00124466 3.3 0.00124458 3.3 0.00124468 0 0.0012446 0 0.0012447 3.3 0.0012446199999999999 3.3 0.00124472 0 0.00124464 0 0.00124474 3.3 0.0012446599999999999 3.3 0.00124476 0 0.00124468 0 0.00124478 3.3 0.0012446999999999998 3.3 0.0012448 0 0.00124472 0 0.00124482 3.3 0.0012447399999999998 3.3 0.0012448399999999999 0 0.00124476 0 0.00124486 3.3 0.00124478 3.3 0.00124488 0 0.0012448 0 0.0012449 3.3 0.00124482 3.3 0.00124492 0 0.0012448399999999999 0 0.00124494 3.3 0.00124486 3.3 0.00124496 0 0.0012448799999999999 0 0.00124498 3.3 0.0012449 3.3 0.001245 0 0.0012449199999999998 0 0.00124502 3.3 0.00124494 3.3 0.00124504 0 0.0012449599999999998 0 0.0012450599999999999 3.3 0.00124498 3.3 0.00124508 0 0.001245 0 0.0012451 3.3 0.00124502 3.3 0.00124512 0 0.00124504 0 0.00124514 3.3 0.0012450599999999999 3.3 0.00124516 0 0.00124508 0 0.00124518 3.3 0.0012450999999999999 3.3 0.0012452 0 0.00124512 0 0.00124522 3.3 0.0012451399999999998 3.3 0.0012452399999999999 0 0.00124516 0 0.00124526 3.3 0.0012451799999999998 3.3 0.0012452799999999999 0 0.0012452 0 0.0012453 3.3 0.00124522 3.3 0.00124532 0 0.0012452399999999999 0 0.00124534 3.3 0.00124526 3.3 0.00124536 0 0.0012452799999999999 0 0.00124538 3.3 0.0012453 3.3 0.0012454 0 0.0012453199999999998 0 0.00124542 3.3 0.00124534 3.3 0.00124544 0 0.0012453599999999998 0 0.0012454599999999999 3.3 0.00124538 3.3 0.00124548 0 0.0012454 0 0.0012455 3.3 0.00124542 3.3 0.00124552 0 0.00124544 0 0.00124554 3.3 0.0012454599999999999 3.3 0.00124556 0 0.00124548 0 0.00124558 3.3 0.0012454999999999999 3.3 0.0012456 0 0.00124552 0 0.00124562 3.3 0.0012455399999999998 3.3 0.00124564 0 0.00124556 0 0.00124566 3.3 0.0012455799999999998 3.3 0.0012456799999999999 0 0.0012456 0 0.0012457 3.3 0.00124562 3.3 0.00124572 0 0.00124564 0 0.00124574 3.3 0.00124566 3.3 0.00124576 0 0.0012456799999999999 0 0.00124578 3.3 0.0012457 3.3 0.0012458 0 0.0012457199999999999 0 0.00124582 3.3 0.00124574 3.3 0.00124584 0 0.0012457599999999998 0 0.00124586 3.3 0.00124578 3.3 0.00124588 0 0.0012457999999999998 0 0.0012458999999999999 3.3 0.00124582 3.3 0.00124592 0 0.00124584 0 0.00124594 3.3 0.00124586 3.3 0.00124596 0 0.00124588 0 0.00124598 3.3 0.0012458999999999999 3.3 0.001246 0 0.00124592 0 0.00124602 3.3 0.0012459399999999999 3.3 0.00124604 0 0.00124596 0 0.00124606 3.3 0.0012459799999999998 3.3 0.0012460799999999999 0 0.001246 0 0.0012461 3.3 0.0012460199999999998 3.3 0.0012461199999999999 0 0.00124604 0 0.00124614 3.3 0.00124606 3.3 0.00124616 0 0.0012460799999999999 0 0.00124618 3.3 0.0012461 3.3 0.0012462 0 0.0012461199999999999 0 0.00124622 3.3 0.00124614 3.3 0.00124624 0 0.0012461599999999998 0 0.00124626 3.3 0.00124618 3.3 0.00124628 0 0.0012461999999999998 0 0.0012462999999999999 3.3 0.00124622 3.3 0.00124632 0 0.00124624 0 0.00124634 3.3 0.00124626 3.3 0.00124636 0 0.00124628 0 0.00124638 3.3 0.0012462999999999999 3.3 0.0012464 0 0.00124632 0 0.00124642 3.3 0.0012463399999999999 3.3 0.00124644 0 0.00124636 0 0.00124646 3.3 0.0012463799999999998 3.3 0.00124648 0 0.0012464 0 0.0012465 3.3 0.0012464199999999998 3.3 0.0012465199999999999 0 0.00124644 0 0.00124654 3.3 0.00124646 3.3 0.00124656 0 0.00124648 0 0.00124658 3.3 0.0012465 3.3 0.0012466 0 0.0012465199999999999 0 0.00124662 3.3 0.00124654 3.3 0.00124664 0 0.0012465599999999999 0 0.00124666 3.3 0.00124658 3.3 0.00124668 0 0.0012465999999999998 0 0.0012467 3.3 0.00124662 3.3 0.00124672 0 0.0012466399999999998 0 0.0012467399999999999 3.3 0.00124666 3.3 0.00124676 0 0.00124668 0 0.00124678 3.3 0.0012467 3.3 0.0012468 0 0.00124672 0 0.00124682 3.3 0.0012467399999999999 3.3 0.00124684 0 0.00124676 0 0.00124686 3.3 0.0012467799999999999 3.3 0.00124688 0 0.0012468 0 0.0012469 3.3 0.0012468199999999998 3.3 0.0012469199999999999 0 0.00124684 0 0.00124694 3.3 0.00124686 3.3 0.00124696 0 0.00124688 0 0.00124698 3.3 0.0012469 3.3 0.001247 0 0.0012469199999999999 0 0.00124702 3.3 0.00124694 3.3 0.00124704 0 0.0012469599999999999 0 0.00124706 3.3 0.00124698 3.3 0.00124708 0 0.0012469999999999998 0 0.0012471 3.3 0.00124702 3.3 0.00124712 0 0.0012470399999999998 0 0.0012471399999999999 3.3 0.00124706 3.3 0.00124716 0 0.00124708 0 0.00124718 3.3 0.0012471 3.3 0.0012472 0 0.00124712 0 0.00124722 3.3 0.0012471399999999999 3.3 0.00124724 0 0.00124716 0 0.00124726 3.3 0.0012471799999999999 3.3 0.00124728 0 0.0012472 0 0.0012473 3.3 0.0012472199999999998 3.3 0.00124732 0 0.00124724 0 0.00124734 3.3 0.0012472599999999998 3.3 0.0012473599999999999 0 0.00124728 0 0.00124738 3.3 0.0012473 3.3 0.0012474 0 0.00124732 0 0.00124742 3.3 0.00124734 3.3 0.00124744 0 0.0012473599999999999 0 0.00124746 3.3 0.00124738 3.3 0.00124748 0 0.0012473999999999999 0 0.0012475 3.3 0.00124742 3.3 0.00124752 0 0.0012474399999999998 0 0.0012475399999999999 3.3 0.00124746 3.3 0.00124756 0 0.0012474799999999998 0 0.0012475799999999999 3.3 0.0012475 3.3 0.0012476 0 0.00124752 0 0.00124762 3.3 0.0012475399999999999 3.3 0.00124764 0 0.00124756 0 0.00124766 3.3 0.0012475799999999999 3.3 0.00124768 0 0.0012476 0 0.0012477 3.3 0.0012476199999999998 3.3 0.00124772 0 0.00124764 0 0.00124774 3.3 0.0012476599999999998 3.3 0.0012477599999999999 0 0.00124768 0 0.00124778 3.3 0.0012477 3.3 0.0012478 0 0.00124772 0 0.00124782 3.3 0.00124774 3.3 0.00124784 0 0.0012477599999999999 0 0.00124786 3.3 0.00124778 3.3 0.00124788 0 0.0012477999999999999 0 0.0012479 3.3 0.00124782 3.3 0.00124792 0 0.0012478399999999998 0 0.00124794 3.3 0.00124786 3.3 0.00124796 0 0.0012478799999999998 0 0.0012479799999999999 3.3 0.0012479 3.3 0.001248 0 0.00124792 0 0.00124802 3.3 0.00124794 3.3 0.00124804 0 0.00124796 0 0.00124806 3.3 0.0012479799999999999 3.3 0.00124808 0 0.001248 0 0.0012481 3.3 0.0012480199999999999 3.3 0.00124812 0 0.00124804 0 0.00124814 3.3 0.0012480599999999998 3.3 0.00124816 0 0.00124808 0 0.00124818 3.3 0.0012480999999999998 3.3 0.0012481999999999999 0 0.00124812 0 0.00124822 3.3 0.00124814 3.3 0.00124824 0 0.00124816 0 0.00124826 3.3 0.00124818 3.3 0.00124828 0 0.0012481999999999999 0 0.0012483 3.3 0.00124822 3.3 0.00124832 0 0.0012482399999999999 0 0.00124834 3.3 0.00124826 3.3 0.00124836 0 0.0012482799999999998 0 0.0012483799999999999 3.3 0.0012483 3.3 0.0012484 0 0.0012483199999999998 0 0.0012484199999999999 3.3 0.00124834 3.3 0.00124844 0 0.00124836 0 0.00124846 3.3 0.0012483799999999999 3.3 0.00124848 0 0.0012484 0 0.0012485 3.3 0.0012484199999999999 3.3 0.00124852 0 0.00124844 0 0.00124854 3.3 0.0012484599999999998 3.3 0.00124856 0 0.00124848 0 0.00124858 3.3 0.0012484999999999998 3.3 0.0012485999999999999 0 0.00124852 0 0.00124862 3.3 0.00124854 3.3 0.00124864 0 0.00124856 0 0.00124866 3.3 0.00124858 3.3 0.00124868 0 0.0012485999999999999 0 0.0012487 3.3 0.00124862 3.3 0.00124872 0 0.0012486399999999999 0 0.00124874 3.3 0.00124866 3.3 0.00124876 0 0.0012486799999999998 0 0.00124878 3.3 0.0012487 3.3 0.0012488 0 0.0012487199999999998 0 0.0012488199999999999 3.3 0.00124874 3.3 0.00124884 0 0.00124876 0 0.00124886 3.3 0.00124878 3.3 0.00124888 0 0.0012488 0 0.0012489 3.3 0.0012488199999999999 3.3 0.00124892 0 0.00124884 0 0.00124894 3.3 0.0012488599999999999 3.3 0.00124896 0 0.00124888 0 0.00124898 3.3 0.0012488999999999998 3.3 0.001249 0 0.00124892 0 0.00124902 3.3 0.0012489399999999998 3.3 0.0012490399999999999 0 0.00124896 0 0.00124906 3.3 0.00124898 3.3 0.00124908 0 0.001249 0 0.0012491 3.3 0.00124902 3.3 0.00124912 0 0.0012490399999999999 0 0.00124914 3.3 0.00124906 3.3 0.00124916 0 0.0012490799999999999 0 0.00124918 3.3 0.0012491 3.3 0.0012492 0 0.0012491199999999998 0 0.0012492199999999999 3.3 0.00124914 3.3 0.00124924 0 0.0012491599999999998 0 0.0012492599999999999 3.3 0.00124918 3.3 0.00124928 0 0.0012492 0 0.0012493 3.3 0.0012492199999999999 3.3 0.00124932 0 0.00124924 0 0.00124934 3.3 0.0012492599999999999 3.3 0.00124936 0 0.00124928 0 0.00124938 3.3 0.0012492999999999998 3.3 0.0012494 0 0.00124932 0 0.00124942 3.3 0.0012493399999999998 3.3 0.0012494399999999999 0 0.00124936 0 0.00124946 3.3 0.00124938 3.3 0.00124948 0 0.0012494 0 0.0012495 3.3 0.00124942 3.3 0.00124952 0 0.0012494399999999999 0 0.00124954 3.3 0.00124946 3.3 0.00124956 0 0.0012494799999999999 0 0.00124958 3.3 0.0012495 3.3 0.0012496 0 0.0012495199999999998 0 0.00124962 3.3 0.00124954 3.3 0.00124964 0 0.0012495599999999998 0 0.0012496599999999999 3.3 0.00124958 3.3 0.00124968 0 0.0012496 0 0.0012497 3.3 0.00124962 3.3 0.00124972 0 0.00124964 0 0.00124974 3.3 0.0012496599999999999 3.3 0.00124976 0 0.00124968 0 0.00124978 3.3 0.0012496999999999999 3.3 0.0012498 0 0.00124972 0 0.00124982 3.3 0.0012497399999999998 3.3 0.00124984 0 0.00124976 0 0.00124986 3.3 0.0012497799999999998 3.3 0.0012498799999999999 0 0.0012498 0 0.0012499 3.3 0.00124982 3.3 0.00124992 0 0.00124984 0 0.00124994 3.3 0.00124986 3.3 0.00124996 0 0.0012498799999999999 0 0.00124998 3.3 0.0012499 3.3 0.00125 0 0.0012499199999999999 0 0.00125002 3.3 0.00124994 3.3 0.00125004 0 0.0012499599999999998 0 0.0012500599999999999 3.3 0.00124998 3.3 0.00125008 0 0.00125 0 0.0012501 3.3 0.00125002 3.3 0.00125012 0 0.00125004 0 0.00125014 3.3 0.0012500599999999999 3.3 0.00125016 0 0.00125008 0 0.00125018 3.3 0.0012500999999999999 3.3 0.0012502 0 0.00125012 0 0.00125022 3.3 0.0012501399999999998 3.3 0.00125024 0 0.00125016 0 0.00125026 3.3 0.0012501799999999998 3.3 0.0012502799999999999 0 0.0012502 0 0.0012503 3.3 0.00125022 3.3 0.00125032 0 0.00125024 0 0.00125034 3.3 0.00125026 3.3 0.00125036 0 0.0012502799999999999 0 0.00125038 3.3 0.0012503 3.3 0.0012504 0 0.0012503199999999999 0 0.00125042 3.3 0.00125034 3.3 0.00125044 0 0.0012503599999999998 0 0.00125046 3.3 0.00125038 3.3 0.00125048 0 0.0012503999999999998 0 0.0012504999999999999 3.3 0.00125042 3.3 0.00125052 0 0.00125044 0 0.00125054 3.3 0.00125046 3.3 0.00125056 0 0.00125048 0 0.00125058 3.3 0.0012504999999999999 3.3 0.0012506 0 0.00125052 0 0.00125062 3.3 0.0012505399999999999 3.3 0.00125064 0 0.00125056 0 0.00125066 3.3 0.0012505799999999998 3.3 0.0012506799999999999 0 0.0012506 0 0.0012507 3.3 0.0012506199999999998 3.3 0.0012507199999999999 0 0.00125064 0 0.00125074 3.3 0.00125066 3.3 0.00125076 0 0.0012506799999999999 0 0.00125078 3.3 0.0012507 3.3 0.0012508 0 0.0012507199999999999 0 0.00125082 3.3 0.00125074 3.3 0.00125084 0 0.0012507599999999998 0 0.00125086 3.3 0.00125078 3.3 0.00125088 0 0.0012507999999999998 0 0.0012508999999999999 3.3 0.00125082 3.3 0.00125092 0 0.00125084 0 0.00125094 3.3 0.00125086 3.3 0.00125096 0 0.00125088 0 0.00125098 3.3 0.0012508999999999999 3.3 0.001251 0 0.00125092 0 0.00125102 3.3 0.0012509399999999999 3.3 0.00125104 0 0.00125096 0 0.00125106 3.3 0.0012509799999999998 3.3 0.00125108 0 0.001251 0 0.0012511 3.3 0.0012510199999999998 3.3 0.0012511199999999999 0 0.00125104 0 0.00125114 3.3 0.00125106 3.3 0.00125116 0 0.00125108 0 0.00125118 3.3 0.0012511 3.3 0.0012512 0 0.0012511199999999999 0 0.00125122 3.3 0.00125114 3.3 0.00125124 0 0.0012511599999999999 0 0.00125126 3.3 0.00125118 3.3 0.00125128 0 0.0012511999999999998 0 0.0012513 3.3 0.00125122 3.3 0.00125132 0 0.0012512399999999998 0 0.0012513399999999999 3.3 0.00125126 3.3 0.00125136 0 0.00125128 0 0.00125138 3.3 0.0012513 3.3 0.0012514 0 0.00125132 0 0.00125142 3.3 0.0012513399999999999 3.3 0.00125144 0 0.00125136 0 0.00125146 3.3 0.0012513799999999999 3.3 0.00125148 0 0.0012514 0 0.0012515 3.3 0.0012514199999999998 3.3 0.0012515199999999999 0 0.00125144 0 0.00125154 3.3 0.0012514599999999998 3.3 0.0012515599999999999 0 0.00125148 0 0.00125158 3.3 0.0012515 3.3 0.0012516 0 0.0012515199999999999 0 0.00125162 3.3 0.00125154 3.3 0.00125164 0 0.0012515599999999999 0 0.00125166 3.3 0.00125158 3.3 0.00125168 0 0.0012515999999999998 0 0.0012517 3.3 0.00125162 3.3 0.00125172 0 0.0012516399999999998 0 0.0012517399999999999 3.3 0.00125166 3.3 0.00125176 0 0.00125168 0 0.00125178 3.3 0.0012517 3.3 0.0012518 0 0.00125172 0 0.00125182 3.3 0.0012517399999999999 3.3 0.00125184 0 0.00125176 0 0.00125186 3.3 0.0012517799999999999 3.3 0.00125188 0 0.0012518 0 0.0012519 3.3 0.0012518199999999998 3.3 0.00125192 0 0.00125184 0 0.00125194 3.3 0.0012518599999999998 3.3 0.0012519599999999999 0 0.00125188 0 0.00125198 3.3 0.0012519 3.3 0.001252 0 0.00125192 0 0.00125202 3.3 0.00125194 3.3 0.00125204 0 0.0012519599999999999 0 0.00125206 3.3 0.00125198 3.3 0.00125208 0 0.0012519999999999999 0 0.0012521 3.3 0.00125202 3.3 0.00125212 0 0.0012520399999999998 0 0.00125214 3.3 0.00125206 3.3 0.00125216 0 0.0012520799999999998 0 0.0012521799999999999 3.3 0.0012521 3.3 0.0012522 0 0.00125212 0 0.00125222 3.3 0.00125214 3.3 0.00125224 0 0.00125216 0 0.00125226 3.3 0.0012521799999999999 3.3 0.00125228 0 0.0012522 0 0.0012523 3.3 0.0012522199999999999 3.3 0.00125232 0 0.00125224 0 0.00125234 3.3 0.0012522599999999998 3.3 0.0012523599999999999 0 0.00125228 0 0.00125238 3.3 0.0012522999999999998 3.3 0.0012523999999999999 0 0.00125232 0 0.00125242 3.3 0.00125234 3.3 0.00125244 0 0.0012523599999999999 0 0.00125246 3.3 0.00125238 3.3 0.00125248 0 0.0012523999999999999 0 0.0012525 3.3 0.00125242 3.3 0.00125252 0 0.0012524399999999998 0 0.00125254 3.3 0.00125246 3.3 0.00125256 0 0.0012524799999999998 0 0.0012525799999999999 3.3 0.0012525 3.3 0.0012526 0 0.00125252 0 0.00125262 3.3 0.00125254 3.3 0.00125264 0 0.00125256 0 0.00125266 3.3 0.0012525799999999999 3.3 0.00125268 0 0.0012526 0 0.0012527 3.3 0.0012526199999999999 3.3 0.00125272 0 0.00125264 0 0.00125274 3.3 0.0012526599999999998 3.3 0.00125276 0 0.00125268 0 0.00125278 3.3 0.0012526999999999998 3.3 0.0012527999999999999 0 0.00125272 0 0.00125282 3.3 0.00125274 3.3 0.00125284 0 0.00125276 0 0.00125286 3.3 0.00125278 3.3 0.00125288 0 0.0012527999999999999 0 0.0012529 3.3 0.00125282 3.3 0.00125292 0 0.0012528399999999999 0 0.00125294 3.3 0.00125286 3.3 0.00125296 0 0.0012528799999999998 0 0.00125298 3.3 0.0012529 3.3 0.001253 0 0.0012529199999999998 0 0.0012530199999999999 3.3 0.00125294 3.3 0.00125304 0 0.00125296 0 0.00125306 3.3 0.00125298 3.3 0.00125308 0 0.001253 0 0.0012531 3.3 0.0012530199999999999 3.3 0.00125312 0 0.00125304 0 0.00125314 3.3 0.0012530599999999999 3.3 0.00125316 0 0.00125308 0 0.00125318 3.3 0.0012530999999999998 3.3 0.0012531999999999999 0 0.00125312 0 0.00125322 3.3 0.00125314 3.3 0.00125324 0 0.00125316 0 0.00125326 3.3 0.00125318 3.3 0.00125328 0 0.0012531999999999999 0 0.0012533 3.3 0.00125322 3.3 0.00125332 0 0.0012532399999999999 0 0.00125334 3.3 0.00125326 3.3 0.00125336 0 0.0012532799999999998 0 0.00125338 3.3 0.0012533 3.3 0.0012534 0 0.0012533199999999998 0 0.0012534199999999999 3.3 0.00125334 3.3 0.00125344 0 0.00125336 0 0.00125346 3.3 0.00125338 3.3 0.00125348 0 0.0012534 0 0.0012535 3.3 0.0012534199999999999 3.3 0.00125352 0 0.00125344 0 0.00125354 3.3 0.0012534599999999999 3.3 0.00125356 0 0.00125348 0 0.00125358 3.3 0.0012534999999999998 3.3 0.0012536 0 0.00125352 0 0.00125362 3.3 0.0012535399999999998 3.3 0.0012536399999999999 0 0.00125356 0 0.00125366 3.3 0.00125358 3.3 0.00125368 0 0.0012536 0 0.0012537 3.3 0.00125362 3.3 0.00125372 0 0.0012536399999999999 0 0.00125374 3.3 0.00125366 3.3 0.00125376 0 0.0012536799999999999 0 0.00125378 3.3 0.0012537 3.3 0.0012538 0 0.0012537199999999998 0 0.0012538199999999999 3.3 0.00125374 3.3 0.00125384 0 0.0012537599999999998 0 0.0012538599999999999 3.3 0.00125378 3.3 0.00125388 0 0.0012538 0 0.0012539 3.3 0.0012538199999999999 3.3 0.00125392 0 0.00125384 0 0.00125394 3.3 0.0012538599999999999 3.3 0.00125396 0 0.00125388 0 0.00125398 3.3 0.0012538999999999998 3.3 0.001254 0 0.00125392 0 0.00125402 3.3 0.0012539399999999998 3.3 0.0012540399999999999 0 0.00125396 0 0.00125406 3.3 0.00125398 3.3 0.00125408 0 0.001254 0 0.0012541 3.3 0.00125402 3.3 0.00125412 0 0.0012540399999999999 0 0.00125414 3.3 0.00125406 3.3 0.00125416 0 0.0012540799999999999 0 0.00125418 3.3 0.0012541 3.3 0.0012542 0 0.0012541199999999998 0 0.00125422 3.3 0.00125414 3.3 0.00125424 0 0.0012541599999999998 0 0.0012542599999999999 3.3 0.00125418 3.3 0.00125428 0 0.0012542 0 0.0012543 3.3 0.00125422 3.3 0.00125432 0 0.00125424 0 0.00125434 3.3 0.0012542599999999999 3.3 0.00125436 0 0.00125428 0 0.00125438 3.3 0.0012542999999999999 3.3 0.0012544 0 0.00125432 0 0.00125442 3.3 0.0012543399999999998 3.3 0.00125444 0 0.00125436 0 0.00125446 3.3 0.0012543799999999998 3.3 0.0012544799999999999 0 0.0012544 0 0.0012545 3.3 0.00125442 3.3 0.00125452 0 0.00125444 0 0.00125454 3.3 0.00125446 3.3 0.00125456 0 0.0012544799999999999 0 0.00125458 3.3 0.0012545 3.3 0.0012546 0 0.0012545199999999999 0 0.00125462 3.3 0.00125454 3.3 0.00125464 0 0.0012545599999999998 0 0.0012546599999999999 3.3 0.00125458 3.3 0.00125468 0 0.0012545999999999998 0 0.0012546999999999999 3.3 0.00125462 3.3 0.00125472 0 0.00125464 0 0.00125474 3.3 0.0012546599999999999 3.3 0.00125476 0 0.00125468 0 0.00125478 3.3 0.0012546999999999999 3.3 0.0012548 0 0.00125472 0 0.00125482 3.3 0.0012547399999999998 3.3 0.00125484 0 0.00125476 0 0.00125486 3.3 0.0012547799999999998 3.3 0.0012548799999999999 0 0.0012548 0 0.0012549 3.3 0.00125482 3.3 0.00125492 0 0.00125484 0 0.00125494 3.3 0.00125486 3.3 0.00125496 0 0.0012548799999999999 0 0.00125498 3.3 0.0012549 3.3 0.001255 0 0.0012549199999999999 0 0.00125502 3.3 0.00125494 3.3 0.00125504 0 0.0012549599999999998 0 0.00125506 3.3 0.00125498 3.3 0.00125508 0 0.0012549999999999998 0 0.0012550999999999999 3.3 0.00125502 3.3 0.00125512 0 0.00125504 0 0.00125514 3.3 0.00125506 3.3 0.00125516 0 0.00125508 0 0.00125518 3.3 0.0012550999999999999 3.3 0.0012552 0 0.00125512 0 0.00125522 3.3 0.0012551399999999999 3.3 0.00125524 0 0.00125516 0 0.00125526 3.3 0.0012551799999999998 3.3 0.00125528 0 0.0012552 0 0.0012553 3.3 0.0012552199999999998 3.3 0.0012553199999999999 0 0.00125524 0 0.00125534 3.3 0.00125526 3.3 0.00125536 0 0.00125528 0 0.00125538 3.3 0.0012553 3.3 0.0012554 0 0.0012553199999999999 0 0.00125542 3.3 0.00125534 3.3 0.00125544 0 0.0012553599999999999 0 0.00125546 3.3 0.00125538 3.3 0.00125548 0 0.0012553999999999998 0 0.0012554999999999999 3.3 0.00125542 3.3 0.00125552 0 0.0012554399999999998 0 0.0012555399999999999 3.3 0.00125546 3.3 0.00125556 0 0.00125548 0 0.00125558 3.3 0.0012554999999999999 3.3 0.0012556 0 0.00125552 0 0.00125562 3.3 0.0012555399999999999 3.3 0.00125564 0 0.00125556 0 0.00125566 3.3 0.0012555799999999998 3.3 0.00125568 0 0.0012556 0 0.0012557 3.3 0.0012556199999999998 3.3 0.0012557199999999999 0 0.00125564 0 0.00125574 3.3 0.00125566 3.3 0.00125576 0 0.00125568 0 0.00125578 3.3 0.0012557 3.3 0.0012558 0 0.0012557199999999999 0 0.00125582 3.3 0.00125574 3.3 0.00125584 0 0.0012557599999999999 0 0.00125586 3.3 0.00125578 3.3 0.00125588 0 0.0012557999999999998 0 0.0012559 3.3 0.00125582 3.3 0.00125592 0 0.0012558399999999998 0 0.0012559399999999999 3.3 0.00125586 3.3 0.00125596 0 0.00125588 0 0.00125598 3.3 0.0012559 3.3 0.001256 0 0.00125592 0 0.00125602 3.3 0.0012559399999999999 3.3 0.00125604 0 0.00125596 0 0.00125606 3.3 0.0012559799999999999 3.3 0.00125608 0 0.001256 0 0.0012561 3.3 0.0012560199999999998 3.3 0.00125612 0 0.00125604 0 0.00125614 3.3 0.0012560599999999998 3.3 0.0012561599999999999 0 0.00125608 0 0.00125618 3.3 0.0012561 3.3 0.0012562 0 0.00125612 0 0.00125622 3.3 0.00125614 3.3 0.00125624 0 0.0012561599999999999 0 0.00125626 3.3 0.00125618 3.3 0.00125628 0 0.0012561999999999999 0 0.0012563 3.3 0.00125622 3.3 0.00125632 0 0.0012562399999999998 0 0.0012563399999999999 3.3 0.00125626 3.3 0.00125636 0 0.0012562799999999998 0 0.0012563799999999999 3.3 0.0012563 3.3 0.0012564 0 0.00125632 0 0.00125642 3.3 0.0012563399999999999 3.3 0.00125644 0 0.00125636 0 0.00125646 3.3 0.0012563799999999999 3.3 0.00125648 0 0.0012564 0 0.0012565 3.3 0.0012564199999999998 3.3 0.00125652 0 0.00125644 0 0.00125654 3.3 0.0012564599999999998 3.3 0.0012565599999999999 0 0.00125648 0 0.00125658 3.3 0.0012565 3.3 0.0012566 0 0.00125652 0 0.00125662 3.3 0.00125654 3.3 0.00125664 0 0.0012565599999999999 0 0.00125666 3.3 0.00125658 3.3 0.00125668 0 0.0012565999999999999 0 0.0012567 3.3 0.00125662 3.3 0.00125672 0 0.0012566399999999998 0 0.00125674 3.3 0.00125666 3.3 0.00125676 0 0.0012566799999999998 0 0.0012567799999999999 3.3 0.0012567 3.3 0.0012568 0 0.00125672 0 0.00125682 3.3 0.00125674 3.3 0.00125684 0 0.00125676 0 0.00125686 3.3 0.0012567799999999999 3.3 0.00125688 0 0.0012568 0 0.0012569 3.3 0.0012568199999999999 3.3 0.00125692 0 0.00125684 0 0.00125694 3.3 0.0012568599999999998 3.3 0.00125696 0 0.00125688 0 0.00125698 3.3 0.0012568999999999998 3.3 0.0012569999999999999 0 0.00125692 0 0.00125702 3.3 0.00125694 3.3 0.00125704 0 0.00125696 0 0.00125706 3.3 0.00125698 3.3 0.00125708 0 0.0012569999999999999 0 0.0012571 3.3 0.00125702 3.3 0.00125712 0 0.0012570399999999999 0 0.00125714 3.3 0.00125706 3.3 0.00125716 0 0.0012570799999999998 0 0.0012571799999999999 3.3 0.0012571 3.3 0.0012572 0 0.00125712 0 0.00125722 3.3 0.00125714 3.3 0.00125724 0 0.00125716 0 0.00125726 3.3 0.0012571799999999999 3.3 0.00125728 0 0.0012572 0 0.0012573 3.3 0.0012572199999999999 3.3 0.00125732 0 0.00125724 0 0.00125734 3.3 0.0012572599999999998 3.3 0.00125736 0 0.00125728 0 0.00125738 3.3 0.0012572999999999998 3.3 0.0012573999999999999 0 0.00125732 0 0.00125742 3.3 0.00125734 3.3 0.00125744 0 0.00125736 0 0.00125746 3.3 0.00125738 3.3 0.00125748 0 0.0012573999999999999 0 0.0012575 3.3 0.00125742 3.3 0.00125752 0 0.0012574399999999999 0 0.00125754 3.3 0.00125746 3.3 0.00125756 0 0.0012574799999999998 0 0.00125758 3.3 0.0012575 3.3 0.0012576 0 0.0012575199999999998 0 0.0012576199999999999 3.3 0.00125754 3.3 0.00125764 0 0.00125756 0 0.00125766 3.3 0.00125758 3.3 0.00125768 0 0.0012576 0 0.0012577 3.3 0.0012576199999999999 3.3 0.00125772 0 0.00125764 0 0.00125774 3.3 0.0012576599999999999 3.3 0.00125776 0 0.00125768 0 0.00125778 3.3 0.0012576999999999998 3.3 0.0012577999999999999 0 0.00125772 0 0.00125782 3.3 0.0012577399999999998 3.3 0.0012578399999999999 0 0.00125776 0 0.00125786 3.3 0.00125778 3.3 0.00125788 0 0.0012577999999999999 0 0.0012579 3.3 0.00125782 3.3 0.00125792 0 0.0012578399999999999 0 0.00125794 3.3 0.00125786 3.3 0.00125796 0 0.0012578799999999998 0 0.00125798 3.3 0.0012579 3.3 0.001258 0 0.0012579199999999998 0 0.0012580199999999999 3.3 0.00125794 3.3 0.00125804 0 0.00125796 0 0.00125806 3.3 0.00125798 3.3 0.00125808 0 0.001258 0 0.0012581 3.3 0.0012580199999999999 3.3 0.00125812 0 0.00125804 0 0.00125814 3.3 0.0012580599999999999 3.3 0.00125816 0 0.00125808 0 0.00125818 3.3 0.0012580999999999998 3.3 0.0012582 0 0.00125812 0 0.00125822 3.3 0.0012581399999999998 3.3 0.0012582399999999999 0 0.00125816 0 0.00125826 3.3 0.00125818 3.3 0.00125828 0 0.0012582 0 0.0012583 3.3 0.00125822 3.3 0.00125832 0 0.0012582399999999999 0 0.00125834 3.3 0.00125826 3.3 0.00125836 0 0.0012582799999999999 0 0.00125838 3.3 0.0012583 3.3 0.0012584 0 0.0012583199999999998 0 0.00125842 3.3 0.00125834 3.3 0.00125844 0 0.0012583599999999998 0 0.0012584599999999999 3.3 0.00125838 3.3 0.00125848 0 0.0012584 0 0.0012585 3.3 0.00125842 3.3 0.00125852 0 0.00125844 0 0.00125854 3.3 0.0012584599999999999 3.3 0.00125856 0 0.00125848 0 0.00125858 3.3 0.0012584999999999999 3.3 0.0012586 0 0.00125852 0 0.00125862 3.3 0.0012585399999999998 3.3 0.0012586399999999999 0 0.00125856 0 0.00125866 3.3 0.0012585799999999998 3.3 0.0012586799999999999 0 0.0012586 0 0.0012587 3.3 0.00125862 3.3 0.00125872 0 0.0012586399999999999 0 0.00125874 3.3 0.00125866 3.3 0.00125876 0 0.0012586799999999999 0 0.00125878 3.3 0.0012587 3.3 0.0012588 0 0.0012587199999999998 0 0.00125882 3.3 0.00125874 3.3 0.00125884 0 0.0012587599999999998 0 0.0012588599999999999 3.3 0.00125878 3.3 0.00125888 0 0.0012588 0 0.0012589 3.3 0.00125882 3.3 0.00125892 0 0.00125884 0 0.00125894 3.3 0.0012588599999999999 3.3 0.00125896 0 0.00125888 0 0.00125898 3.3 0.0012588999999999999 3.3 0.001259 0 0.00125892 0 0.00125902 3.3 0.0012589399999999998 3.3 0.00125904 0 0.00125896 0 0.00125906 3.3 0.0012589799999999998 3.3 0.0012590799999999999 0 0.001259 0 0.0012591 3.3 0.00125902 3.3 0.00125912 0 0.00125904 0 0.00125914 3.3 0.00125906 3.3 0.00125916 0 0.0012590799999999999 0 0.00125918 3.3 0.0012591 3.3 0.0012592 0 0.0012591199999999999 0 0.00125922 3.3 0.00125914 3.3 0.00125924 0 0.0012591599999999998 0 0.00125926 3.3 0.00125918 3.3 0.00125928 0 0.0012591999999999998 0 0.0012592999999999999 3.3 0.00125922 3.3 0.00125932 0 0.00125924 0 0.00125934 3.3 0.00125926 3.3 0.00125936 0 0.00125928 0 0.00125938 3.3 0.0012592999999999999 3.3 0.0012594 0 0.00125932 0 0.00125942 3.3 0.0012593399999999999 3.3 0.00125944 0 0.00125936 0 0.00125946 3.3 0.0012593799999999998 3.3 0.0012594799999999999 0 0.0012594 0 0.0012595 3.3 0.0012594199999999998 3.3 0.0012595199999999999 0 0.00125944 0 0.00125954 3.3 0.00125946 3.3 0.00125956 0 0.0012594799999999999 0 0.00125958 3.3 0.0012595 3.3 0.0012596 0 0.0012595199999999999 0 0.00125962 3.3 0.00125954 3.3 0.00125964 0 0.0012595599999999998 0 0.00125966 3.3 0.00125958 3.3 0.00125968 0 0.0012595999999999998 0 0.0012596999999999999 3.3 0.00125962 3.3 0.00125972 0 0.00125964 0 0.00125974 3.3 0.00125966 3.3 0.00125976 0 0.00125968 0 0.00125978 3.3 0.0012596999999999999 3.3 0.0012598 0 0.00125972 0 0.00125982 3.3 0.0012597399999999999 3.3 0.00125984 0 0.00125976 0 0.00125986 3.3 0.0012597799999999998 3.3 0.00125988 0 0.0012598 0 0.0012599 3.3 0.0012598199999999998 3.3 0.0012599199999999999 0 0.00125984 0 0.00125994 3.3 0.00125986 3.3 0.00125996 0 0.00125988 0 0.00125998 3.3 0.0012599 3.3 0.00126 0 0.0012599199999999999 0 0.00126002 3.3 0.00125994 3.3 0.00126004 0 0.0012599599999999999 0 0.00126006 3.3 0.00125998 3.3 0.00126008 0 0.0012599999999999998 0 0.0012601 3.3 0.00126002 3.3 0.00126012 0 0.0012600399999999998 0 0.0012601399999999999 3.3 0.00126006 3.3 0.00126016 0 0.00126008 0 0.00126018 3.3 0.0012601 3.3 0.0012602 0 0.00126012 0 0.00126022 3.3 0.0012601399999999999 3.3 0.00126024 0 0.00126016 0 0.00126026 3.3 0.0012601799999999999 3.3 0.00126028 0 0.0012602 0 0.0012603 3.3 0.0012602199999999998 3.3 0.0012603199999999999 0 0.00126024 0 0.00126034 3.3 0.00126026 3.3 0.00126036 0 0.00126028 0 0.00126038 3.3 0.0012603 3.3 0.0012604 0 0.0012603199999999999 0 0.00126042 3.3 0.00126034 3.3 0.00126044 0 0.0012603599999999999 0 0.00126046 3.3 0.00126038 3.3 0.00126048 0 0.0012603999999999998 0 0.0012605 3.3 0.00126042 3.3 0.00126052 0 0.0012604399999999998 0 0.0012605399999999999 3.3 0.00126046 3.3 0.00126056 0 0.00126048 0 0.00126058 3.3 0.0012605 3.3 0.0012606 0 0.00126052 0 0.00126062 3.3 0.0012605399999999999 3.3 0.00126064 0 0.00126056 0 0.00126066 3.3 0.0012605799999999999 3.3 0.00126068 0 0.0012606 0 0.0012607 3.3 0.0012606199999999998 3.3 0.00126072 0 0.00126064 0 0.00126074 3.3 0.0012606599999999998 3.3 0.0012607599999999999 0 0.00126068 0 0.00126078 3.3 0.0012607 3.3 0.0012608 0 0.00126072 0 0.00126082 3.3 0.00126074 3.3 0.00126084 0 0.0012607599999999999 0 0.00126086 3.3 0.00126078 3.3 0.00126088 0 0.0012607999999999999 0 0.0012609 3.3 0.00126082 3.3 0.00126092 0 0.0012608399999999998 0 0.0012609399999999999 3.3 0.00126086 3.3 0.00126096 0 0.0012608799999999998 0 0.0012609799999999999 3.3 0.0012609 3.3 0.001261 0 0.00126092 0 0.00126102 3.3 0.0012609399999999999 3.3 0.00126104 0 0.00126096 0 0.00126106 3.3 0.0012609799999999999 3.3 0.00126108 0 0.001261 0 0.0012611 3.3 0.0012610199999999998 3.3 0.00126112 0 0.00126104 0 0.00126114 3.3 0.0012610599999999998 3.3 0.0012611599999999999 0 0.00126108 0 0.00126118 3.3 0.0012611 3.3 0.0012612 0 0.00126112 0 0.00126122 3.3 0.00126114 3.3 0.00126124 0 0.0012611599999999999 0 0.00126126 3.3 0.00126118 3.3 0.00126128 0 0.0012611999999999999 0 0.0012613 3.3 0.00126122 3.3 0.00126132 0 0.0012612399999999998 0 0.00126134 3.3 0.00126126 3.3 0.00126136 0 0.0012612799999999998 0 0.0012613799999999999 3.3 0.0012613 3.3 0.0012614 0 0.00126132 0 0.00126142 3.3 0.00126134 3.3 0.00126144 0 0.00126136 0 0.00126146 3.3 0.0012613799999999999 3.3 0.00126148 0 0.0012614 0 0.0012615 3.3 0.0012614199999999999 3.3 0.00126152 0 0.00126144 0 0.00126154 3.3 0.0012614599999999998 3.3 0.00126156 0 0.00126148 0 0.00126158 3.3 0.0012614999999999998 3.3 0.0012615999999999999 0 0.00126152 0 0.00126162 3.3 0.00126154 3.3 0.00126164 0 0.00126156 0 0.00126166 3.3 0.00126158 3.3 0.00126168 0 0.0012615999999999999 0 0.0012617 3.3 0.00126162 3.3 0.00126172 0 0.0012616399999999999 0 0.00126174 3.3 0.00126166 3.3 0.00126176 0 0.0012616799999999998 0 0.0012617799999999999 3.3 0.0012617 3.3 0.0012618 0 0.0012617199999999998 0 0.0012618199999999999 3.3 0.00126174 3.3 0.00126184 0 0.00126176 0 0.00126186 3.3 0.0012617799999999999 3.3 0.00126188 0 0.0012618 0 0.0012619 3.3 0.0012618199999999999 3.3 0.00126192 0 0.00126184 0 0.00126194 3.3 0.0012618599999999998 3.3 0.00126196 0 0.00126188 0 0.00126198 3.3 0.0012618999999999998 3.3 0.0012619999999999999 0 0.00126192 0 0.00126202 3.3 0.00126194 3.3 0.00126204 0 0.00126196 0 0.00126206 3.3 0.00126198 3.3 0.00126208 0 0.0012619999999999999 0 0.0012621 3.3 0.00126202 3.3 0.00126212 0 0.0012620399999999999 0 0.00126214 3.3 0.00126206 3.3 0.00126216 0 0.0012620799999999998 0 0.00126218 3.3 0.0012621 3.3 0.0012622 0 0.0012621199999999998 0 0.0012622199999999999 3.3 0.00126214 3.3 0.00126224 0 0.00126216 0 0.00126226 3.3 0.00126218 3.3 0.00126228 0 0.0012622 0 0.0012623 3.3 0.0012622199999999999 3.3 0.00126232 0 0.00126224 0 0.00126234 3.3 0.0012622599999999999 3.3 0.00126236 0 0.00126228 0 0.00126238 3.3 0.0012622999999999998 3.3 0.0012624 0 0.00126232 0 0.00126242 3.3 0.0012623399999999998 3.3 0.0012624399999999999 0 0.00126236 0 0.00126246 3.3 0.00126238 3.3 0.00126248 0 0.0012624 0 0.0012625 3.3 0.00126242 3.3 0.00126252 0 0.0012624399999999999 0 0.00126254 3.3 0.00126246 3.3 0.00126256 0 0.0012624799999999999 0 0.00126258 3.3 0.0012625 3.3 0.0012626 0 0.0012625199999999998 0 0.0012626199999999999 3.3 0.00126254 3.3 0.00126264 0 0.0012625599999999998 0 0.0012626599999999999 3.3 0.00126258 3.3 0.00126268 0 0.0012626 0 0.0012627 3.3 0.0012626199999999999 3.3 0.00126272 0 0.00126264 0 0.00126274 3.3 0.0012626599999999999 3.3 0.00126276 0 0.00126268 0 0.00126278 3.3 0.0012626999999999998 3.3 0.0012628 0 0.00126272 0 0.00126282 3.3 0.0012627399999999998 3.3 0.0012628399999999999 0 0.00126276 0 0.00126286 3.3 0.00126278 3.3 0.00126288 0 0.0012628 0 0.0012629 3.3 0.00126282 3.3 0.00126292 0 0.0012628399999999999 0 0.00126294 3.3 0.00126286 3.3 0.00126296 0 0.0012628799999999999 0 0.00126298 3.3 0.0012629 3.3 0.001263 0 0.0012629199999999998 0 0.00126302 3.3 0.00126294 3.3 0.00126304 0 0.0012629599999999998 0 0.0012630599999999999 3.3 0.00126298 3.3 0.00126308 0 0.001263 0 0.0012631 3.3 0.00126302 3.3 0.00126312 0 0.00126304 0 0.00126314 3.3 0.0012630599999999999 3.3 0.00126316 0 0.00126308 0 0.00126318 3.3 0.0012630999999999999 3.3 0.0012632 0 0.00126312 0 0.00126322 3.3 0.0012631399999999998 3.3 0.00126324 0 0.00126316 0 0.00126326 3.3 0.0012631799999999998 3.3 0.0012632799999999999 0 0.0012632 0 0.0012633 3.3 0.00126322 3.3 0.00126332 0 0.00126324 0 0.00126334 3.3 0.00126326 3.3 0.00126336 0 0.0012632799999999999 0 0.00126338 3.3 0.0012633 3.3 0.0012634 0 0.0012633199999999999 0 0.00126342 3.3 0.00126334 3.3 0.00126344 0 0.0012633599999999998 0 0.0012634599999999999 3.3 0.00126338 3.3 0.00126348 0 0.0012633999999999998 0 0.0012634999999999999 3.3 0.00126342 3.3 0.00126352 0 0.00126344 0 0.00126354 3.3 0.0012634599999999999 3.3 0.00126356 0 0.00126348 0 0.00126358 3.3 0.0012634999999999999 3.3 0.0012636 0 0.00126352 0 0.00126362 3.3 0.0012635399999999998 3.3 0.00126364 0 0.00126356 0 0.00126366 3.3 0.0012635799999999998 3.3 0.0012636799999999999 0 0.0012636 0 0.0012637 3.3 0.00126362 3.3 0.00126372 0 0.00126364 0 0.00126374 3.3 0.00126366 3.3 0.00126376 0 0.0012636799999999999 0 0.00126378 3.3 0.0012637 3.3 0.0012638 0 0.0012637199999999999 0 0.00126382 3.3 0.00126374 3.3 0.00126384 0 0.0012637599999999998 0 0.00126386 3.3 0.00126378 3.3 0.00126388 0 0.0012637999999999998 0 0.0012638999999999999 3.3 0.00126382 3.3 0.00126392 0 0.00126384 0 0.00126394 3.3 0.00126386 3.3 0.00126396 0 0.00126388 0 0.00126398 3.3 0.0012638999999999999 3.3 0.001264 0 0.00126392 0 0.00126402 3.3 0.0012639399999999999 3.3 0.00126404 0 0.00126396 0 0.00126406 3.3 0.0012639799999999998 3.3 0.0012640799999999999 0 0.001264 0 0.0012641 3.3 0.0012640199999999998 3.3 0.0012641199999999999 0 0.00126404 0 0.00126414 3.3 0.00126406 3.3 0.00126416 0 0.0012640799999999999 0 0.00126418 3.3 0.0012641 3.3 0.0012642 0 0.0012641199999999999 0 0.00126422 3.3 0.00126414 3.3 0.00126424 0 0.0012641599999999998 0 0.00126426 3.3 0.00126418 3.3 0.00126428 0 0.0012641999999999998 0 0.0012642999999999999 3.3 0.00126422 3.3 0.00126432 0 0.00126424 0 0.00126434 3.3 0.00126426 3.3 0.00126436 0 0.00126428 0 0.00126438 3.3 0.0012642999999999999 3.3 0.0012644 0 0.00126432 0 0.00126442 3.3 0.0012643399999999999 3.3 0.00126444 0 0.00126436 0 0.00126446 3.3 0.0012643799999999998 3.3 0.00126448 0 0.0012644 0 0.0012645 3.3 0.0012644199999999998 3.3 0.0012645199999999999 0 0.00126444 0 0.00126454 3.3 0.00126446 3.3 0.00126456 0 0.00126448 0 0.00126458 3.3 0.0012645 3.3 0.0012646 0 0.0012645199999999999 0 0.00126462 3.3 0.00126454 3.3 0.00126464 0 0.0012645599999999999 0 0.00126466 3.3 0.00126458 3.3 0.00126468 0 0.0012645999999999998 0 0.0012647 3.3 0.00126462 3.3 0.00126472 0 0.0012646399999999998 0 0.0012647399999999999 3.3 0.00126466 3.3 0.00126476 0 0.00126468 0 0.00126478 3.3 0.0012647 3.3 0.0012648 0 0.00126472 0 0.00126482 3.3 0.0012647399999999999 3.3 0.00126484 0 0.00126476 0 0.00126486 3.3 0.0012647799999999999 3.3 0.00126488 0 0.0012648 0 0.0012649 3.3 0.0012648199999999998 3.3 0.0012649199999999999 0 0.00126484 0 0.00126494 3.3 0.0012648599999999998 3.3 0.0012649599999999999 0 0.00126488 0 0.00126498 3.3 0.0012649 3.3 0.001265 0 0.0012649199999999999 0 0.00126502 3.3 0.00126494 3.3 0.00126504 0 0.0012649599999999999 0 0.00126506 3.3 0.00126498 3.3 0.00126508 0 0.0012649999999999998 0 0.0012651 3.3 0.00126502 3.3 0.00126512 0 0.0012650399999999998 0 0.0012651399999999999 3.3 0.00126506 3.3 0.00126516 0 0.00126508 0 0.00126518 3.3 0.0012651 3.3 0.0012652 0 0.00126512 0 0.00126522 3.3 0.0012651399999999999 3.3 0.00126524 0 0.00126516 0 0.00126526 3.3 0.0012651799999999999 3.3 0.00126528 0 0.0012652 0 0.0012653 3.3 0.0012652199999999998 3.3 0.00126532 0 0.00126524 0 0.00126534 3.3 0.0012652599999999998 3.3 0.0012653599999999999 0 0.00126528 0 0.00126538 3.3 0.0012653 3.3 0.0012654 0 0.00126532 0 0.00126542 3.3 0.00126534 3.3 0.00126544 0 0.0012653599999999999 0 0.00126546 3.3 0.00126538 3.3 0.00126548 0 0.0012653999999999999 0 0.0012655 3.3 0.00126542 3.3 0.00126552 0 0.0012654399999999998 0 0.00126554 3.3 0.00126546 3.3 0.00126556 0 0.0012654799999999998 0 0.0012655799999999999 3.3 0.0012655 3.3 0.0012656 0 0.00126552 0 0.00126562 3.3 0.00126554 3.3 0.00126564 0 0.00126556 0 0.00126566 3.3 0.0012655799999999999 3.3 0.00126568 0 0.0012656 0 0.0012657 3.3 0.0012656199999999999 3.3 0.00126572 0 0.00126564 0 0.00126574 3.3 0.0012656599999999998 3.3 0.0012657599999999999 0 0.00126568 0 0.00126578 3.3 0.0012656999999999998 3.3 0.0012657999999999999 0 0.00126572 0 0.00126582 3.3 0.00126574 3.3 0.00126584 0 0.0012657599999999999 0 0.00126586 3.3 0.00126578 3.3 0.00126588 0 0.0012657999999999999 0 0.0012659 3.3 0.00126582 3.3 0.00126592 0 0.0012658399999999998 0 0.00126594 3.3 0.00126586 3.3 0.00126596 0 0.0012658799999999998 0 0.0012659799999999999 3.3 0.0012659 3.3 0.001266 0 0.00126592 0 0.00126602 3.3 0.00126594 3.3 0.00126604 0 0.00126596 0 0.00126606 3.3 0.0012659799999999999 3.3 0.00126608 0 0.001266 0 0.0012661 3.3 0.0012660199999999999 3.3 0.00126612 0 0.00126604 0 0.00126614 3.3 0.0012660599999999998 3.3 0.00126616 0 0.00126608 0 0.00126618 3.3 0.0012660999999999998 3.3 0.0012661999999999999 0 0.00126612 0 0.00126622 3.3 0.00126614 3.3 0.00126624 0 0.00126616 0 0.00126626 3.3 0.00126618 3.3 0.00126628 0 0.0012661999999999999 0 0.0012663 3.3 0.00126622 3.3 0.00126632 0 0.0012662399999999999 0 0.00126634 3.3 0.00126626 3.3 0.00126636 0 0.0012662799999999998 0 0.00126638 3.3 0.0012663 3.3 0.0012664 0 0.0012663199999999998 0 0.0012664199999999999 3.3 0.00126634 3.3 0.00126644 0 0.00126636 0 0.00126646 3.3 0.00126638 3.3 0.00126648 0 0.0012664 0 0.0012665 3.3 0.0012664199999999999 3.3 0.00126652 0 0.00126644 0 0.00126654 3.3 0.0012664599999999999 3.3 0.00126656 0 0.00126648 0 0.00126658 3.3 0.0012664999999999998 3.3 0.0012665999999999999 0 0.00126652 0 0.00126662 3.3 0.0012665399999999998 3.3 0.0012666399999999999 0 0.00126656 0 0.00126666 3.3 0.00126658 3.3 0.00126668 0 0.0012665999999999999 0 0.0012667 3.3 0.00126662 3.3 0.00126672 0 0.0012666399999999999 0 0.00126674 3.3 0.00126666 3.3 0.00126676 0 0.0012666799999999998 0 0.00126678 3.3 0.0012667 3.3 0.0012668 0 0.0012667199999999998 0 0.0012668199999999999 3.3 0.00126674 3.3 0.00126684 0 0.00126676 0 0.00126686 3.3 0.00126678 3.3 0.00126688 0 0.0012668 0 0.0012669 3.3 0.0012668199999999999 3.3 0.00126692 0 0.00126684 0 0.00126694 3.3 0.0012668599999999999 3.3 0.00126696 0 0.00126688 0 0.00126698 3.3 0.0012668999999999998 3.3 0.001267 0 0.00126692 0 0.00126702 3.3 0.0012669399999999998 3.3 0.0012670399999999999 0 0.00126696 0 0.00126706 3.3 0.00126698 3.3 0.00126708 0 0.001267 0 0.0012671 3.3 0.00126702 3.3 0.00126712 0 0.0012670399999999999 0 0.00126714 3.3 0.00126706 3.3 0.00126716 0 0.0012670799999999999 0 0.00126718 3.3 0.0012671 3.3 0.0012672 0 0.0012671199999999998 0 0.00126722 3.3 0.00126714 3.3 0.00126724 0 0.0012671599999999998 0 0.0012672599999999999 3.3 0.00126718 3.3 0.00126728 0 0.0012672 0 0.0012673 3.3 0.00126722 3.3 0.00126732 0 0.00126724 0 0.00126734 3.3 0.0012672599999999999 3.3 0.00126736 0 0.00126728 0 0.00126738 3.3 0.0012672999999999999 3.3 0.0012674 0 0.00126732 0 0.00126742 3.3 0.0012673399999999998 3.3 0.0012674399999999999 0 0.00126736 0 0.00126746 3.3 0.00126738 3.3 0.00126748 0 0.0012674 0 0.0012675 3.3 0.00126742 3.3 0.00126752 0 0.0012674399999999999 0 0.00126754 3.3 0.00126746 3.3 0.00126756 0 0.0012674799999999999 0 0.00126758 3.3 0.0012675 3.3 0.0012676 0 0.0012675199999999998 0 0.00126762 3.3 0.00126754 3.3 0.00126764 0 0.0012675599999999998 0 0.0012676599999999999 3.3 0.00126758 3.3 0.00126768 0 0.0012676 0 0.0012677 3.3 0.00126762 3.3 0.00126772 0 0.00126764 0 0.00126774 3.3 0.0012676599999999999 3.3 0.00126776 0 0.00126768 0 0.00126778 3.3 0.0012676999999999999 3.3 0.0012678 0 0.00126772 0 0.00126782 3.3 0.0012677399999999998 3.3 0.00126784 0 0.00126776 0 0.00126786 3.3 0.0012677799999999998 3.3 0.0012678799999999999 0 0.0012678 0 0.0012679 3.3 0.00126782 3.3 0.00126792 0 0.00126784 0 0.00126794 3.3 0.00126786 3.3 0.00126796 0 0.0012678799999999999 0 0.00126798 3.3 0.0012679 3.3 0.001268 0 0.0012679199999999999 0 0.00126802 3.3 0.00126794 3.3 0.00126804 0 0.0012679599999999998 0 0.0012680599999999999 3.3 0.00126798 3.3 0.00126808 0 0.0012679999999999998 0 0.0012680999999999999 3.3 0.00126802 3.3 0.00126812 0 0.00126804 0 0.00126814 3.3 0.0012680599999999999 3.3 0.00126816 0 0.00126808 0 0.00126818 3.3 0.0012680999999999999 3.3 0.0012682 0 0.00126812 0 0.00126822 3.3 0.0012681399999999998 3.3 0.00126824 0 0.00126816 0 0.00126826 3.3 0.0012681799999999998 3.3 0.0012682799999999999 0 0.0012682 0 0.0012683 3.3 0.00126822 3.3 0.00126832 0 0.00126824 0 0.00126834 3.3 0.00126826 3.3 0.00126836 0 0.0012682799999999999 0 0.00126838 3.3 0.0012683 3.3 0.0012684 0 0.0012683199999999999 0 0.00126842 3.3 0.00126834 3.3 0.00126844 0 0.0012683599999999998 0 0.00126846 3.3 0.00126838 3.3 0.00126848 0 0.0012683999999999998 0 0.0012684999999999999 3.3 0.00126842 3.3 0.00126852 0 0.00126844 0 0.00126854 3.3 0.00126846 3.3 0.00126856 0 0.00126848 0 0.00126858 3.3 0.0012684999999999999 3.3 0.0012686 0 0.00126852 0 0.00126862 3.3 0.0012685399999999999 3.3 0.00126864 0 0.00126856 0 0.00126866 3.3 0.0012685799999999998 3.3 0.00126868 0 0.0012686 0 0.0012687 3.3 0.0012686199999999998 3.3 0.0012687199999999999 0 0.00126864 0 0.00126874 3.3 0.00126866 3.3 0.00126876 0 0.00126868 0 0.00126878 3.3 0.0012687 3.3 0.0012688 0 0.0012687199999999999 0 0.00126882 3.3 0.00126874 3.3 0.00126884 0 0.0012687599999999999 0 0.00126886 3.3 0.00126878 3.3 0.00126888 0 0.0012687999999999998 0 0.0012688999999999999 3.3 0.00126882 3.3 0.00126892 0 0.0012688399999999998 0 0.0012689399999999999 3.3 0.00126886 3.3 0.00126896 0 0.00126888 0 0.00126898 3.3 0.0012688999999999999 3.3 0.001269 0 0.00126892 0 0.00126902 3.3 0.0012689399999999999 3.3 0.00126904 0 0.00126896 0 0.00126906 3.3 0.0012689799999999998 3.3 0.00126908 0 0.001269 0 0.0012691 3.3 0.0012690199999999998 3.3 0.0012691199999999999 0 0.00126904 0 0.00126914 3.3 0.00126906 3.3 0.00126916 0 0.00126908 0 0.00126918 3.3 0.0012691 3.3 0.0012692 0 0.0012691199999999999 0 0.00126922 3.3 0.00126914 3.3 0.00126924 0 0.0012691599999999999 0 0.00126926 3.3 0.00126918 3.3 0.00126928 0 0.0012691999999999998 0 0.0012693 3.3 0.00126922 3.3 0.00126932 0 0.0012692399999999998 0 0.0012693399999999999 3.3 0.00126926 3.3 0.00126936 0 0.00126928 0 0.00126938 3.3 0.0012693 3.3 0.0012694 0 0.00126932 0 0.00126942 3.3 0.0012693399999999999 3.3 0.00126944 0 0.00126936 0 0.00126946 3.3 0.0012693799999999999 3.3 0.00126948 0 0.0012694 0 0.0012695 3.3 0.0012694199999999998 3.3 0.00126952 0 0.00126944 0 0.00126954 3.3 0.0012694599999999998 3.3 0.0012695599999999999 0 0.00126948 0 0.00126958 3.3 0.0012695 3.3 0.0012696 0 0.00126952 0 0.00126962 3.3 0.00126954 3.3 0.00126964 0 0.0012695599999999999 0 0.00126966 3.3 0.00126958 3.3 0.00126968 0 0.0012695999999999999 0 0.0012697 3.3 0.00126962 3.3 0.00126972 0 0.0012696399999999998 0 0.0012697399999999999 3.3 0.00126966 3.3 0.00126976 0 0.0012696799999999998 0 0.0012697799999999999 3.3 0.0012697 3.3 0.0012698 0 0.00126972 0 0.00126982 3.3 0.0012697399999999999 3.3 0.00126984 0 0.00126976 0 0.00126986 3.3 0.0012697799999999999 3.3 0.00126988 0 0.0012698 0 0.0012699 3.3 0.0012698199999999998 3.3 0.00126992 0 0.00126984 0 0.00126994 3.3 0.0012698599999999998 3.3 0.0012699599999999999 0 0.00126988 0 0.00126998 3.3 0.0012699 3.3 0.00127 0 0.00126992 0 0.00127002 3.3 0.00126994 3.3 0.00127004 0 0.0012699599999999999 0 0.00127006 3.3 0.00126998 3.3 0.00127008 0 0.0012699999999999999 0 0.0012701 3.3 0.00127002 3.3 0.00127012 0 0.0012700399999999998 0 0.00127014 3.3 0.00127006 3.3 0.00127016 0 0.0012700799999999998 0 0.0012701799999999999 3.3 0.0012701 3.3 0.0012702 0 0.00127012 0 0.00127022 3.3 0.00127014 3.3 0.00127024 0 0.00127016 0 0.00127026 3.3 0.0012701799999999999 3.3 0.00127028 0 0.0012702 0 0.0012703 3.3 0.0012702199999999999 3.3 0.00127032 0 0.00127024 0 0.00127034 3.3 0.0012702599999999998 3.3 0.00127036 0 0.00127028 0 0.00127038 3.3 0.0012702999999999998 3.3 0.0012703999999999999 0 0.00127032 0 0.00127042 3.3 0.00127034 3.3 0.00127044 0 0.00127036 0 0.00127046 3.3 0.00127038 3.3 0.00127048 0 0.0012703999999999999 0 0.0012705 3.3 0.00127042 3.3 0.00127052 0 0.0012704399999999999 0 0.00127054 3.3 0.00127046 3.3 0.00127056 0 0.0012704799999999998 0 0.0012705799999999999 3.3 0.0012705 3.3 0.0012706 0 0.00127052 0 0.00127062 3.3 0.00127054 3.3 0.00127064 0 0.00127056 0 0.00127066 3.3 0.0012705799999999999 3.3 0.00127068 0 0.0012706 0 0.0012707 3.3 0.0012706199999999999 3.3 0.00127072 0 0.00127064 0 0.00127074 3.3 0.0012706599999999998 3.3 0.00127076 0 0.00127068 0 0.00127078 3.3 0.0012706999999999998 3.3 0.0012707999999999999 0 0.00127072 0 0.00127082 3.3 0.00127074 3.3 0.00127084 0 0.00127076 0 0.00127086 3.3 0.00127078 3.3 0.00127088 0 0.0012707999999999999 0 0.0012709 3.3 0.00127082 3.3 0.00127092 0 0.0012708399999999999 0 0.00127094 3.3 0.00127086 3.3 0.00127096 0 0.0012708799999999998 0 0.00127098 3.3 0.0012709 3.3 0.001271 0 0.0012709199999999998 0 0.0012710199999999999 3.3 0.00127094 3.3 0.00127104 0 0.00127096 0 0.00127106 3.3 0.00127098 3.3 0.00127108 0 0.001271 0 0.0012711 3.3 0.0012710199999999999 3.3 0.00127112 0 0.00127104 0 0.00127114 3.3 0.0012710599999999999 3.3 0.00127116 0 0.00127108 0 0.00127118 3.3 0.0012710999999999998 3.3 0.0012711999999999999 0 0.00127112 0 0.00127122 3.3 0.0012711399999999998 3.3 0.0012712399999999999 0 0.00127116 0 0.00127126 3.3 0.00127118 3.3 0.00127128 0 0.0012711999999999999 0 0.0012713 3.3 0.00127122 3.3 0.00127132 0 0.0012712399999999999 0 0.00127134 3.3 0.00127126 3.3 0.00127136 0 0.0012712799999999998 0 0.00127138 3.3 0.0012713 3.3 0.0012714 0 0.0012713199999999998 0 0.0012714199999999999 3.3 0.00127134 3.3 0.00127144 0 0.00127136 0 0.00127146 3.3 0.00127138 3.3 0.00127148 0 0.0012714 0 0.0012715 3.3 0.0012714199999999999 3.3 0.00127152 0 0.00127144 0 0.00127154 3.3 0.0012714599999999999 3.3 0.00127156 0 0.00127148 0 0.00127158 3.3 0.0012714999999999998 3.3 0.0012716 0 0.00127152 0 0.00127162 3.3 0.0012715399999999998 3.3 0.0012716399999999999 0 0.00127156 0 0.00127166 3.3 0.00127158 3.3 0.00127168 0 0.0012716 0 0.0012717 3.3 0.00127162 3.3 0.00127172 0 0.0012716399999999999 0 0.00127174 3.3 0.00127166 3.3 0.00127176 0 0.0012716799999999999 0 0.00127178 3.3 0.0012717 3.3 0.0012718 0 0.0012717199999999998 0 0.00127182 3.3 0.00127174 3.3 0.00127184 0 0.0012717599999999998 0 0.0012718599999999999 3.3 0.00127178 3.3 0.00127188 0 0.0012718 0 0.0012719 3.3 0.00127182 3.3 0.00127192 0 0.00127184 0 0.00127194 3.3 0.0012718599999999999 3.3 0.00127196 0 0.00127188 0 0.00127198 3.3 0.0012718999999999999 3.3 0.001272 0 0.00127192 0 0.00127202 3.3 0.0012719399999999998 3.3 0.0012720399999999999 0 0.00127196 0 0.00127206 3.3 0.0012719799999999998 3.3 0.0012720799999999999 0 0.001272 0 0.0012721 3.3 0.00127202 3.3 0.00127212 0 0.0012720399999999999 0 0.00127214 3.3 0.00127206 3.3 0.00127216 0 0.0012720799999999999 0 0.00127218 3.3 0.0012721 3.3 0.0012722 0 0.0012721199999999998 0 0.00127222 3.3 0.00127214 3.3 0.00127224 0 0.0012721599999999998 0 0.0012722599999999999 3.3 0.00127218 3.3 0.00127228 0 0.0012722 0 0.0012723 3.3 0.00127222 3.3 0.00127232 0 0.00127224 0 0.00127234 3.3 0.0012722599999999999 3.3 0.00127236 0 0.00127228 0 0.00127238 3.3 0.0012722999999999999 3.3 0.0012724 0 0.00127232 0 0.00127242 3.3 0.0012723399999999998 3.3 0.00127244 0 0.00127236 0 0.00127246 3.3 0.0012723799999999998 3.3 0.0012724799999999999 0 0.0012724 0 0.0012725 3.3 0.00127242 3.3 0.00127252 0 0.00127244 0 0.00127254 3.3 0.00127246 3.3 0.00127256 0 0.0012724799999999999 0 0.00127258 3.3 0.0012725 3.3 0.0012726 0 0.0012725199999999999 0 0.00127262 3.3 0.00127254 3.3 0.00127264 0 0.0012725599999999998 0 0.00127266 3.3 0.00127258 3.3 0.00127268 0 0.0012725999999999998 0 0.0012726999999999999 3.3 0.00127262 3.3 0.00127272 0 0.00127264 0 0.00127274 3.3 0.00127266 3.3 0.00127276 0 0.00127268 0 0.00127278 3.3 0.0012726999999999999 3.3 0.0012728 0 0.00127272 0 0.00127282 3.3 0.0012727399999999999 3.3 0.00127284 0 0.00127276 0 0.00127286 3.3 0.0012727799999999998 3.3 0.0012728799999999999 0 0.0012728 0 0.0012729 3.3 0.0012728199999999998 3.3 0.0012729199999999999 0 0.00127284 0 0.00127294 3.3 0.00127286 3.3 0.00127296 0 0.0012728799999999999 0 0.00127298 3.3 0.0012729 3.3 0.001273 0 0.0012729199999999999 0 0.00127302 3.3 0.00127294 3.3 0.00127304 0 0.0012729599999999998 0 0.00127306 3.3 0.00127298 3.3 0.00127308 0 0.0012729999999999998 0 0.0012730999999999999 3.3 0.00127302 3.3 0.00127312 0 0.00127304 0 0.00127314 3.3 0.00127306 3.3 0.00127316 0 0.00127308 0 0.00127318 3.3 0.0012730999999999999 3.3 0.0012732 0 0.00127312 0 0.00127322 3.3 0.0012731399999999999 3.3 0.00127324 0 0.00127316 0 0.00127326 3.3 0.0012731799999999998 3.3 0.00127328 0 0.0012732 0 0.0012733 3.3 0.0012732199999999998 3.3 0.0012733199999999999 0 0.00127324 0 0.00127334 3.3 0.00127326 3.3 0.00127336 0 0.00127328 0 0.00127338 3.3 0.0012733 3.3 0.0012734 0 0.0012733199999999999 0 0.00127342 3.3 0.00127334 3.3 0.00127344 0 0.0012733599999999999 0 0.00127346 3.3 0.00127338 3.3 0.00127348 0 0.0012733999999999998 0 0.0012735 3.3 0.00127342 3.3 0.00127352 0 0.0012734399999999998 0 0.0012735399999999999 3.3 0.00127346 3.3 0.00127356 0 0.00127348 0 0.00127358 3.3 0.0012735 3.3 0.0012736 0 0.00127352 0 0.00127362 3.3 0.0012735399999999999 3.3 0.00127364 0 0.00127356 0 0.00127366 3.3 0.0012735799999999999 3.3 0.00127368 0 0.0012736 0 0.0012737 3.3 0.0012736199999999998 3.3 0.0012737199999999999 0 0.00127364 0 0.00127374 3.3 0.0012736599999999998 3.3 0.0012737599999999999 0 0.00127368 0 0.00127378 3.3 0.0012737 3.3 0.0012738 0 0.0012737199999999999 0 0.00127382 3.3 0.00127374 3.3 0.00127384 0 0.0012737599999999999 0 0.00127386 3.3 0.00127378 3.3 0.00127388 0 0.0012737999999999998 0 0.0012739 3.3 0.00127382 3.3 0.00127392 0 0.0012738399999999998 0 0.0012739399999999999 3.3 0.00127386 3.3 0.00127396 0 0.00127388 0 0.00127398 3.3 0.0012739 3.3 0.001274 0 0.00127392 0 0.00127402 3.3 0.0012739399999999999 3.3 0.00127404 0 0.00127396 0 0.00127406 3.3 0.0012739799999999999 3.3 0.00127408 0 0.001274 0 0.0012741 3.3 0.0012740199999999998 3.3 0.00127412 0 0.00127404 0 0.00127414 3.3 0.0012740599999999998 3.3 0.0012741599999999999 0 0.00127408 0 0.00127418 3.3 0.0012741 3.3 0.0012742 0 0.00127412 0 0.00127422 3.3 0.00127414 3.3 0.00127424 0 0.0012741599999999999 0 0.00127426 3.3 0.00127418 3.3 0.00127428 0 0.0012741999999999999 0 0.0012743 3.3 0.00127422 3.3 0.00127432 0 0.0012742399999999998 0 0.0012743399999999999 3.3 0.00127426 3.3 0.00127436 0 0.0012742799999999998 0 0.0012743799999999999 3.3 0.0012743 3.3 0.0012744 0 0.00127432 0 0.00127442 3.3 0.0012743399999999999 3.3 0.00127444 0 0.00127436 0 0.00127446 3.3 0.0012743799999999999 3.3 0.00127448 0 0.0012744 0 0.0012745 3.3 0.0012744199999999998 3.3 0.00127452 0 0.00127444 0 0.00127454 3.3 0.0012744599999999998 3.3 0.0012745599999999999 0 0.00127448 0 0.00127458 3.3 0.0012745 3.3 0.0012746 0 0.00127452 0 0.00127462 3.3 0.00127454 3.3 0.00127464 0 0.0012745599999999999 0 0.00127466 3.3 0.00127458 3.3 0.00127468 0 0.0012745999999999999 0 0.0012747 3.3 0.00127462 3.3 0.00127472 0 0.0012746399999999998 0 0.00127474 3.3 0.00127466 3.3 0.00127476 0 0.0012746799999999998 0 0.0012747799999999999 3.3 0.0012747 3.3 0.0012748 0 0.00127472 0 0.00127482 3.3 0.00127474 3.3 0.00127484 0 0.00127476 0 0.00127486 3.3 0.0012747799999999999 3.3 0.00127488 0 0.0012748 0 0.0012749 3.3 0.0012748199999999999 3.3 0.00127492 0 0.00127484 0 0.00127494 3.3 0.0012748599999999998 3.3 0.00127496 0 0.00127488 0 0.00127498 3.3 0.0012748999999999998 3.3 0.0012749999999999999 0 0.00127492 0 0.00127502 3.3 0.00127494 3.3 0.00127504 0 0.00127496 0 0.00127506 3.3 0.00127498 3.3 0.00127508 0 0.0012749999999999999 0 0.0012751 3.3 0.00127502 3.3 0.00127512 0 0.0012750399999999999 0 0.00127514 3.3 0.00127506 3.3 0.00127516 0 0.0012750799999999998 0 0.0012751799999999999 3.3 0.0012751 3.3 0.0012752 0 0.0012751199999999998 0 0.0012752199999999999 3.3 0.00127514 3.3 0.00127524 0 0.00127516 0 0.00127526 3.3 0.0012751799999999999 3.3 0.00127528 0 0.0012752 0 0.0012753 3.3 0.0012752199999999999 3.3 0.00127532 0 0.00127524 0 0.00127534 3.3 0.0012752599999999998 3.3 0.00127536 0 0.00127528 0 0.00127538 3.3 0.0012752999999999998 3.3 0.0012753999999999999 0 0.00127532 0 0.00127542 3.3 0.00127534 3.3 0.00127544 0 0.00127536 0 0.00127546 3.3 0.00127538 3.3 0.00127548 0 0.0012753999999999999 0 0.0012755 3.3 0.00127542 3.3 0.00127552 0 0.0012754399999999999 0 0.00127554 3.3 0.00127546 3.3 0.00127556 0 0.0012754799999999998 0 0.00127558 3.3 0.0012755 3.3 0.0012756 0 0.0012755199999999998 0 0.0012756199999999999 3.3 0.00127554 3.3 0.00127564 0 0.00127556 0 0.00127566 3.3 0.00127558 3.3 0.00127568 0 0.0012756 0 0.0012757 3.3 0.0012756199999999999 3.3 0.00127572 0 0.00127564 0 0.00127574 3.3 0.0012756599999999999 3.3 0.00127576 0 0.00127568 0 0.00127578 3.3 0.0012756999999999998 3.3 0.0012758 0 0.00127572 0 0.00127582 3.3 0.0012757399999999998 3.3 0.0012758399999999999 0 0.00127576 0 0.00127586 3.3 0.00127578 3.3 0.00127588 0 0.0012758 0 0.0012759 3.3 0.00127582 3.3 0.00127592 0 0.0012758399999999999 0 0.00127594 3.3 0.00127586 3.3 0.00127596 0 0.0012758799999999999 0 0.00127598 3.3 0.0012759 3.3 0.001276 0 0.0012759199999999998 0 0.0012760199999999999 3.3 0.00127594 3.3 0.00127604 0 0.0012759599999999998 0 0.0012760599999999999 3.3 0.00127598 3.3 0.00127608 0 0.001276 0 0.0012761 3.3 0.0012760199999999999 3.3 0.00127612 0 0.00127604 0 0.00127614 3.3 0.0012760599999999999 3.3 0.00127616 0 0.00127608 0 0.00127618 3.3 0.0012760999999999998 3.3 0.0012762 0 0.00127612 0 0.00127622 3.3 0.0012761399999999998 3.3 0.0012762399999999999 0 0.00127616 0 0.00127626 3.3 0.00127618 3.3 0.00127628 0 0.0012762 0 0.0012763 3.3 0.00127622 3.3 0.00127632 0 0.0012762399999999999 0 0.00127634 3.3 0.00127626 3.3 0.00127636 0 0.0012762799999999999 0 0.00127638 3.3 0.0012763 3.3 0.0012764 0 0.0012763199999999998 0 0.00127642 3.3 0.00127634 3.3 0.00127644 0 0.0012763599999999998 0 0.0012764599999999999 3.3 0.00127638 3.3 0.00127648 0 0.0012764 0 0.0012765 3.3 0.00127642 3.3 0.00127652 0 0.00127644 0 0.00127654 3.3 0.0012764599999999999 3.3 0.00127656 0 0.00127648 0 0.00127658 3.3 0.0012764999999999999 3.3 0.0012766 0 0.00127652 0 0.00127662 3.3 0.0012765399999999998 3.3 0.00127664 0 0.00127656 0 0.00127666 3.3 0.0012765799999999998 3.3 0.0012766799999999999 0 0.0012766 0 0.0012767 3.3 0.00127662 3.3 0.00127672 0 0.00127664 0 0.00127674 3.3 0.00127666 3.3 0.00127676 0 0.0012766799999999999 0 0.00127678 3.3 0.0012767 3.3 0.0012768 0 0.0012767199999999999 0 0.00127682 3.3 0.00127674 3.3 0.00127684 0 0.0012767599999999998 0 0.0012768599999999999 3.3 0.00127678 3.3 0.00127688 0 0.0012767999999999998 0 0.0012768999999999999 3.3 0.00127682 3.3 0.00127692 0 0.00127684 0 0.00127694 3.3 0.0012768599999999999 3.3 0.00127696 0 0.00127688 0 0.00127698 3.3 0.0012768999999999999 3.3 0.001277 0 0.00127692 0 0.00127702 3.3 0.0012769399999999998 3.3 0.00127704 0 0.00127696 0 0.00127706 3.3 0.0012769799999999998 3.3 0.0012770799999999999 0 0.001277 0 0.0012771 3.3 0.00127702 3.3 0.00127712 0 0.00127704 0 0.00127714 3.3 0.00127706 3.3 0.00127716 0 0.0012770799999999999 0 0.00127718 3.3 0.0012771 3.3 0.0012772 0 0.0012771199999999999 0 0.00127722 3.3 0.00127714 3.3 0.00127724 0 0.0012771599999999998 0 0.00127726 3.3 0.00127718 3.3 0.00127728 0 0.0012771999999999998 0 0.0012772999999999999 3.3 0.00127722 3.3 0.00127732 0 0.00127724 0 0.00127734 3.3 0.00127726 3.3 0.00127736 0 0.00127728 0 0.00127738 3.3 0.0012772999999999999 3.3 0.0012774 0 0.00127732 0 0.00127742 3.3 0.0012773399999999999 3.3 0.00127744 0 0.00127736 0 0.00127746 3.3 0.0012773799999999998 3.3 0.00127748 0 0.0012774 0 0.0012775 3.3 0.0012774199999999998 3.3 0.0012775199999999999 0 0.00127744 0 0.00127754 3.3 0.00127746 3.3 0.00127756 0 0.00127748 0 0.00127758 3.3 0.0012775 3.3 0.0012776 0 0.0012775199999999999 0 0.00127762 3.3 0.00127754 3.3 0.00127764 0 0.0012775599999999999 0 0.00127766 3.3 0.00127758 3.3 0.00127768 0 0.0012775999999999998 0 0.0012776999999999999 3.3 0.00127762 3.3 0.00127772 0 0.00127764 0 0.00127774 3.3 0.00127766 3.3 0.00127776 0 0.00127768 0 0.00127778 3.3 0.0012776999999999999 3.3 0.0012778 0 0.00127772 0 0.00127782 3.3 0.0012777399999999999 3.3 0.00127784 0 0.00127776 0 0.00127786 3.3 0.0012777799999999998 3.3 0.00127788 0 0.0012778 0 0.0012779 3.3 0.0012778199999999998 3.3 0.0012779199999999999 0 0.00127784 0 0.00127794 3.3 0.00127786 3.3 0.00127796 0 0.00127788 0 0.00127798 3.3 0.0012779 3.3 0.001278 0 0.0012779199999999999 0 0.00127802 3.3 0.00127794 3.3 0.00127804 0 0.0012779599999999999 0 0.00127806 3.3 0.00127798 3.3 0.00127808 0 0.0012779999999999998 0 0.0012781 3.3 0.00127802 3.3 0.00127812 0 0.0012780399999999998 0 0.0012781399999999999 3.3 0.00127806 3.3 0.00127816 0 0.00127808 0 0.00127818 3.3 0.0012781 3.3 0.0012782 0 0.00127812 0 0.00127822 3.3 0.0012781399999999999 3.3 0.00127824 0 0.00127816 0 0.00127826 3.3 0.0012781799999999999 3.3 0.00127828 0 0.0012782 0 0.0012783 3.3 0.0012782199999999998 3.3 0.0012783199999999999 0 0.00127824 0 0.00127834 3.3 0.0012782599999999998 3.3 0.0012783599999999999 0 0.00127828 0 0.00127838 3.3 0.0012783 3.3 0.0012784 0 0.0012783199999999999 0 0.00127842 3.3 0.00127834 3.3 0.00127844 0 0.0012783599999999999 0 0.00127846 3.3 0.00127838 3.3 0.00127848 0 0.0012783999999999998 0 0.0012785 3.3 0.00127842 3.3 0.00127852 0 0.0012784399999999998 0 0.0012785399999999999 3.3 0.00127846 3.3 0.00127856 0 0.00127848 0 0.00127858 3.3 0.0012785 3.3 0.0012786 0 0.00127852 0 0.00127862 3.3 0.0012785399999999999 3.3 0.00127864 0 0.00127856 0 0.00127866 3.3 0.0012785799999999999 3.3 0.00127868 0 0.0012786 0 0.0012787 3.3 0.0012786199999999998 3.3 0.00127872 0 0.00127864 0 0.00127874 3.3 0.0012786599999999998 3.3 0.0012787599999999999 0 0.00127868 0 0.00127878 3.3 0.0012787 3.3 0.0012788 0 0.00127872 0 0.00127882 3.3 0.00127874 3.3 0.00127884 0 0.0012787599999999999 0 0.00127886 3.3 0.00127878 3.3 0.00127888 0 0.0012787999999999999 0 0.0012789 3.3 0.00127882 3.3 0.00127892 0 0.0012788399999999998 0 0.00127894 3.3 0.00127886 3.3 0.00127896 0 0.0012788799999999998 0 0.0012789799999999999 3.3 0.0012789 3.3 0.001279 0 0.00127892 0 0.00127902 3.3 0.00127894 3.3 0.00127904 0 0.00127896 0 0.00127906 3.3 0.0012789799999999999 3.3 0.00127908 0 0.001279 0 0.0012791 3.3 0.0012790199999999999 3.3 0.00127912 0 0.00127904 0 0.00127914 3.3 0.0012790599999999998 3.3 0.0012791599999999999 0 0.00127908 0 0.00127918 3.3 0.0012790999999999998 3.3 0.0012791999999999999 0 0.00127912 0 0.00127922 3.3 0.00127914 3.3 0.00127924 0 0.0012791599999999999 0 0.00127926 3.3 0.00127918 3.3 0.00127928 0 0.0012791999999999999 0 0.0012793 3.3 0.00127922 3.3 0.00127932 0 0.0012792399999999998 0 0.00127934 3.3 0.00127926 3.3 0.00127936 0 0.0012792799999999998 0 0.0012793799999999999 3.3 0.0012793 3.3 0.0012794 0 0.00127932 0 0.00127942 3.3 0.00127934 3.3 0.00127944 0 0.00127936 0 0.00127946 3.3 0.0012793799999999999 3.3 0.00127948 0 0.0012794 0 0.0012795 3.3 0.0012794199999999999 3.3 0.00127952 0 0.00127944 0 0.00127954 3.3 0.0012794599999999998 3.3 0.00127956 0 0.00127948 0 0.00127958 3.3 0.0012794999999999998 3.3 0.0012795999999999999 0 0.00127952 0 0.00127962 3.3 0.00127954 3.3 0.00127964 0 0.00127956 0 0.00127966 3.3 0.00127958 3.3 0.00127968 0 0.0012795999999999999 0 0.0012797 3.3 0.00127962 3.3 0.00127972 0 0.0012796399999999999 0 0.00127974 3.3 0.00127966 3.3 0.00127976 0 0.0012796799999999998 0 0.00127978 3.3 0.0012797 3.3 0.0012798 0 0.0012797199999999998 0 0.0012798199999999999 3.3 0.00127974 3.3 0.00127984 0 0.00127976 0 0.00127986 3.3 0.00127978 3.3 0.00127988 0 0.0012798 0 0.0012799 3.3 0.0012798199999999999 3.3 0.00127992 0 0.00127984 0 0.00127994 3.3 0.0012798599999999999 3.3 0.00127996 0 0.00127988 0 0.00127998 3.3 0.0012798999999999998 3.3 0.0012799999999999999 0 0.00127992 0 0.00128002 3.3 0.0012799399999999998 3.3 0.0012800399999999999 0 0.00127996 0 0.00128006 3.3 0.00127998 3.3 0.00128008 0 0.0012799999999999999 0 0.0012801 3.3 0.00128002 3.3 0.00128012 0 0.0012800399999999999 0 0.00128014 3.3 0.00128006 3.3 0.00128016 0 0.0012800799999999998 0 0.00128018 3.3 0.0012801 3.3 0.0012802 0 0.0012801199999999998 0 0.0012802199999999999 3.3 0.00128014 3.3 0.00128024 0 0.00128016 0 0.00128026 3.3 0.00128018 3.3 0.00128028 0 0.0012802 0 0.0012803 3.3 0.0012802199999999999 3.3 0.00128032 0 0.00128024 0 0.00128034 3.3 0.0012802599999999999 3.3 0.00128036 0 0.00128028 0 0.00128038 3.3 0.0012802999999999998 3.3 0.0012804 0 0.00128032 0 0.00128042 3.3 0.0012803399999999998 3.3 0.0012804399999999999 0 0.00128036 0 0.00128046 3.3 0.00128038 3.3 0.00128048 0 0.0012804 0 0.0012805 3.3 0.00128042 3.3 0.00128052 0 0.0012804399999999999 0 0.00128054 3.3 0.00128046 3.3 0.00128056 0 0.0012804799999999999 0 0.00128058 3.3 0.0012805 3.3 0.0012806 0 0.0012805199999999998 0 0.00128062 3.3 0.00128054 3.3 0.00128064 0 0.0012805599999999998 0 0.0012806599999999999 3.3 0.00128058 3.3 0.00128068 0 0.0012806 0 0.0012807 3.3 0.00128062 3.3 0.00128072 0 0.00128064 0 0.00128074 3.3 0.0012806599999999999 3.3 0.00128076 0 0.00128068 0 0.00128078 3.3 0.0012806999999999999 3.3 0.0012808 0 0.00128072 0 0.00128082 3.3 0.0012807399999999998 3.3 0.0012808399999999999 0 0.00128076 0 0.00128086 3.3 0.0012807799999999998 3.3 0.0012808799999999999 0 0.0012808 0 0.0012809 3.3 0.00128082 3.3 0.00128092 0 0.0012808399999999999 0 0.00128094 3.3 0.00128086 3.3 0.00128096 0 0.0012808799999999999 0 0.00128098 3.3 0.0012809 3.3 0.001281 0 0.0012809199999999998 0 0.00128102 3.3 0.00128094 3.3 0.00128104 0 0.0012809599999999998 0 0.0012810599999999999 3.3 0.00128098 3.3 0.00128108 0 0.001281 0 0.0012811 3.3 0.00128102 3.3 0.00128112 0 0.00128104 0 0.00128114 3.3 0.0012810599999999999 3.3 0.00128116 0 0.00128108 0 0.00128118 3.3 0.0012810999999999999 3.3 0.0012812 0 0.00128112 0 0.00128122 3.3 0.0012811399999999998 3.3 0.00128124 0 0.00128116 0 0.00128126 3.3 0.0012811799999999998 3.3 0.0012812799999999999 0 0.0012812 0 0.0012813 3.3 0.00128122 3.3 0.00128132 0 0.00128124 0 0.00128134 3.3 0.00128126 3.3 0.00128136 0 0.0012812799999999999 0 0.00128138 3.3 0.0012813 3.3 0.0012814 0 0.0012813199999999999 0 0.00128142 3.3 0.00128134 3.3 0.00128144 0 0.0012813599999999998 0 0.0012814599999999999 3.3 0.00128138 3.3 0.00128148 0 0.0012813999999999998 0 0.0012814999999999999 3.3 0.00128142 3.3 0.00128152 0 0.00128144 0 0.00128154 3.3 0.0012814599999999999 3.3 0.00128156 0 0.00128148 0 0.00128158 3.3 0.0012814999999999999 3.3 0.0012816 0 0.00128152 0 0.00128162 3.3 0.0012815399999999998 3.3 0.00128164 0 0.00128156 0 0.00128166 3.3 0.0012815799999999998 3.3 0.0012816799999999999 0 0.0012816 0 0.0012817 3.3 0.00128162 3.3 0.00128172 0 0.00128164 0 0.00128174 3.3 0.00128166 3.3 0.00128176 0 0.0012816799999999999 0 0.00128178 3.3 0.0012817 3.3 0.0012818 0 0.0012817199999999999 0 0.00128182 3.3 0.00128174 3.3 0.00128184 0 0.0012817599999999998 0 0.00128186 3.3 0.00128178 3.3 0.00128188 0 0.0012817999999999998 0 0.0012818999999999999 3.3 0.00128182 3.3 0.00128192 0 0.00128184 0 0.00128194 3.3 0.00128186 3.3 0.00128196 0 0.00128188 0 0.00128198 3.3 0.0012818999999999999 3.3 0.001282 0 0.00128192 0 0.00128202 3.3 0.0012819399999999999 3.3 0.00128204 0 0.00128196 0 0.00128206 3.3 0.0012819799999999998 3.3 0.00128208 0 0.001282 0 0.0012821 3.3 0.0012820199999999998 3.3 0.0012821199999999999 0 0.00128204 0 0.00128214 3.3 0.00128206 3.3 0.00128216 0 0.00128208 0 0.00128218 3.3 0.0012821 3.3 0.0012822 0 0.0012821199999999999 0 0.00128222 3.3 0.00128214 3.3 0.00128224 0 0.0012821599999999999 0 0.00128226 3.3 0.00128218 3.3 0.00128228 0 0.0012821999999999998 0 0.0012822999999999999 3.3 0.00128222 3.3 0.00128232 0 0.0012822399999999998 0 0.0012823399999999999 3.3 0.00128226 3.3 0.00128236 0 0.00128228 0 0.00128238 3.3 0.0012822999999999999 3.3 0.0012824 0 0.00128232 0 0.00128242 3.3 0.0012823399999999999 3.3 0.00128244 0 0.00128236 0 0.00128246 3.3 0.0012823799999999998 3.3 0.00128248 0 0.0012824 0 0.0012825 3.3 0.0012824199999999998 3.3 0.0012825199999999999 0 0.00128244 0 0.00128254 3.3 0.00128246 3.3 0.00128256 0 0.00128248 0 0.00128258 3.3 0.0012825 3.3 0.0012826 0 0.0012825199999999999 0 0.00128262 3.3 0.00128254 3.3 0.00128264 0 0.0012825599999999999 0 0.00128266 3.3 0.00128258 3.3 0.00128268 0 0.0012825999999999998 0 0.0012827 3.3 0.00128262 3.3 0.00128272 0 0.0012826399999999998 0 0.0012827399999999999 3.3 0.00128266 3.3 0.00128276 0 0.00128268 0 0.00128278 3.3 0.0012827 3.3 0.0012828 0 0.00128272 0 0.00128282 3.3 0.0012827399999999999 3.3 0.00128284 0 0.00128276 0 0.00128286 3.3 0.0012827799999999999 3.3 0.00128288 0 0.0012828 0 0.0012829 3.3 0.0012828199999999998 3.3 0.00128292 0 0.00128284 0 0.00128294 3.3 0.0012828599999999998 3.3 0.0012829599999999999 0 0.00128288 0 0.00128298 3.3 0.0012829 3.3 0.001283 0 0.00128292 0 0.00128302 3.3 0.00128294 3.3 0.00128304 0 0.0012829599999999999 0 0.00128306 3.3 0.00128298 3.3 0.00128308 0 0.0012829999999999999 0 0.0012831 3.3 0.00128302 3.3 0.00128312 0 0.0012830399999999998 0 0.0012831399999999999 3.3 0.00128306 3.3 0.00128316 0 0.0012830799999999998 0 0.0012831799999999999 3.3 0.0012831 3.3 0.0012832 0 0.00128312 0 0.00128322 3.3 0.0012831399999999999 3.3 0.00128324 0 0.00128316 0 0.00128326 3.3 0.0012831799999999999 3.3 0.00128328 0 0.0012832 0 0.0012833 3.3 0.0012832199999999998 3.3 0.00128332 0 0.00128324 0 0.00128334 3.3 0.0012832599999999998 3.3 0.0012833599999999999 0 0.00128328 0 0.00128338 3.3 0.0012833 3.3 0.0012834 0 0.00128332 0 0.00128342 3.3 0.00128334 3.3 0.00128344 0 0.0012833599999999999 0 0.00128346 3.3 0.00128338 3.3 0.00128348 0 0.0012833999999999999 0 0.0012835 3.3 0.00128342 3.3 0.00128352 0 0.0012834399999999998 0 0.00128354 3.3 0.00128346 3.3 0.00128356 0 0.0012834799999999998 0 0.0012835799999999999 3.3 0.0012835 3.3 0.0012836 0 0.00128352 0 0.00128362 3.3 0.00128354 3.3 0.00128364 0 0.00128356 0 0.00128366 3.3 0.0012835799999999999 3.3 0.00128368 0 0.0012836 0 0.0012837 3.3 0.0012836199999999999 3.3 0.00128372 0 0.00128364 0 0.00128374 3.3 0.0012836599999999998 3.3 0.00128376 0 0.00128368 0 0.00128378 3.3 0.0012836999999999998 3.3 0.0012837999999999999 0 0.00128372 0 0.00128382 3.3 0.00128374 3.3 0.00128384 0 0.00128376 0 0.00128386 3.3 0.00128378 3.3 0.00128388 0 0.0012837999999999999 0 0.0012839 3.3 0.00128382 3.3 0.00128392 0 0.0012838399999999999 0 0.00128394 3.3 0.00128386 3.3 0.00128396 0 0.0012838799999999998 0 0.0012839799999999999 3.3 0.0012839 3.3 0.001284 0 0.0012839199999999998 0 0.0012840199999999999 3.3 0.00128394 3.3 0.00128404 0 0.00128396 0 0.00128406 3.3 0.0012839799999999999 3.3 0.00128408 0 0.001284 0 0.0012841 3.3 0.0012840199999999999 3.3 0.00128412 0 0.00128404 0 0.00128414 3.3 0.0012840599999999998 3.3 0.00128416 0 0.00128408 0 0.00128418 3.3 0.0012840999999999998 3.3 0.0012841999999999999 0 0.00128412 0 0.00128422 3.3 0.00128414 3.3 0.00128424 0 0.00128416 0 0.00128426 3.3 0.00128418 3.3 0.00128428 0 0.0012841999999999999 0 0.0012843 3.3 0.00128422 3.3 0.00128432 0 0.0012842399999999999 0 0.00128434 3.3 0.00128426 3.3 0.00128436 0 0.0012842799999999998 0 0.00128438 3.3 0.0012843 3.3 0.0012844 0 0.0012843199999999998 0 0.0012844199999999999 3.3 0.00128434 3.3 0.00128444 0 0.00128436 0 0.00128446 3.3 0.00128438 3.3 0.00128448 0 0.0012844 0 0.0012845 3.3 0.0012844199999999999 3.3 0.00128452 0 0.00128444 0 0.00128454 3.3 0.0012844599999999999 3.3 0.00128456 0 0.00128448 0 0.00128458 3.3 0.0012844999999999998 3.3 0.0012845999999999999 0 0.00128452 0 0.00128462 3.3 0.0012845399999999998 3.3 0.0012846399999999999 0 0.00128456 0 0.00128466 3.3 0.00128458 3.3 0.00128468 0 0.0012845999999999999 0 0.0012847 3.3 0.00128462 3.3 0.00128472 0 0.0012846399999999999 0 0.00128474 3.3 0.00128466 3.3 0.00128476 0 0.0012846799999999998 0 0.00128478 3.3 0.0012847 3.3 0.0012848 0 0.0012847199999999998 0 0.0012848199999999999 3.3 0.00128474 3.3 0.00128484 0 0.00128476 0 0.00128486 3.3 0.00128478 3.3 0.00128488 0 0.0012848 0 0.0012849 3.3 0.0012848199999999999 3.3 0.00128492 0 0.00128484 0 0.00128494 3.3 0.0012848599999999999 3.3 0.00128496 0 0.00128488 0 0.00128498 3.3 0.0012848999999999998 3.3 0.001285 0 0.00128492 0 0.00128502 3.3 0.0012849399999999998 3.3 0.0012850399999999999 0 0.00128496 0 0.00128506 3.3 0.00128498 3.3 0.00128508 0 0.001285 0 0.0012851 3.3 0.00128502 3.3 0.00128512 0 0.0012850399999999999 0 0.00128514 3.3 0.00128506 3.3 0.00128516 0 0.0012850799999999999 0 0.00128518 3.3 0.0012851 3.3 0.0012852 0 0.0012851199999999998 0 0.00128522 3.3 0.00128514 3.3 0.00128524 0 0.0012851599999999998 0 0.0012852599999999999 3.3 0.00128518 3.3 0.00128528 0 0.0012852 0 0.0012853 3.3 0.00128522 3.3 0.00128532 0 0.00128524 0 0.00128534 3.3 0.0012852599999999999 3.3 0.00128536 0 0.00128528 0 0.00128538 3.3 0.0012852999999999999 3.3 0.0012854 0 0.00128532 0 0.00128542 3.3 0.0012853399999999998 3.3 0.0012854399999999999 0 0.00128536 0 0.00128546 3.3 0.0012853799999999998 3.3 0.0012854799999999999 0 0.0012854 0 0.0012855 3.3 0.00128542 3.3 0.00128552 0 0.0012854399999999999 0 0.00128554 3.3 0.00128546 3.3 0.00128556 0 0.0012854799999999999 0 0.00128558 3.3 0.0012855 3.3 0.0012856 0 0.0012855199999999998 0 0.00128562 3.3 0.00128554 3.3 0.00128564 0 0.0012855599999999998 0 0.0012856599999999999 3.3 0.00128558 3.3 0.00128568 0 0.0012856 0 0.0012857 3.3 0.00128562 3.3 0.00128572 0 0.00128564 0 0.00128574 3.3 0.0012856599999999999 3.3 0.00128576 0 0.00128568 0 0.00128578 3.3 0.0012856999999999999 3.3 0.0012858 0 0.00128572 0 0.00128582 3.3 0.0012857399999999998 3.3 0.00128584 0 0.00128576 0 0.00128586 3.3 0.0012857799999999998 3.3 0.0012858799999999999 0 0.0012858 0 0.0012859 3.3 0.00128582 3.3 0.00128592 0 0.00128584 0 0.00128594 3.3 0.00128586 3.3 0.00128596 0 0.0012858799999999999 0 0.00128598 3.3 0.0012859 3.3 0.001286 0 0.0012859199999999999 0 0.00128602 3.3 0.00128594 3.3 0.00128604 0 0.0012859599999999998 0 0.00128606 3.3 0.00128598 3.3 0.00128608 0 0.0012859999999999998 0 0.0012860999999999999 3.3 0.00128602 3.3 0.00128612 0 0.00128604 0 0.00128614 3.3 0.00128606 3.3 0.00128616 0 0.00128608 0 0.00128618 3.3 0.0012860999999999999 3.3 0.0012862 0 0.00128612 0 0.00128622 3.3 0.0012861399999999999 3.3 0.00128624 0 0.00128616 0 0.00128626 3.3 0.0012861799999999998 3.3 0.0012862799999999999 0 0.0012862 0 0.0012863 3.3 0.0012862199999999998 3.3 0.0012863199999999999 0 0.00128624 0 0.00128634 3.3 0.00128626 3.3 0.00128636 0 0.0012862799999999999 0 0.00128638 3.3 0.0012863 3.3 0.0012864 0 0.0012863199999999999 0 0.00128642 3.3 0.00128634 3.3 0.00128644 0 0.0012863599999999998 0 0.00128646 3.3 0.00128638 3.3 0.00128648 0 0.0012863999999999998 0 0.0012864999999999999 3.3 0.00128642 3.3 0.00128652 0 0.00128644 0 0.00128654 3.3 0.00128646 3.3 0.00128656 0 0.00128648 0 0.00128658 3.3 0.0012864999999999999 3.3 0.0012866 0 0.00128652 0 0.00128662 3.3 0.0012865399999999999 3.3 0.00128664 0 0.00128656 0 0.00128666 3.3 0.0012865799999999998 3.3 0.00128668 0 0.0012866 0 0.0012867 3.3 0.0012866199999999998 3.3 0.0012867199999999999 0 0.00128664 0 0.00128674 3.3 0.00128666 3.3 0.00128676 0 0.00128668 0 0.00128678 3.3 0.0012867 3.3 0.0012868 0 0.0012867199999999999 0 0.00128682 3.3 0.00128674 3.3 0.00128684 0 0.0012867599999999999 0 0.00128686 3.3 0.00128678 3.3 0.00128688 0 0.0012867999999999998 0 0.0012869 3.3 0.00128682 3.3 0.00128692 0 0.0012868399999999998 0 0.0012869399999999999 3.3 0.00128686 3.3 0.00128696 0 0.00128688 0 0.00128698 3.3 0.0012869 3.3 0.001287 0 0.00128692 0 0.00128702 3.3 0.0012869399999999999 3.3 0.00128704 0 0.00128696 0 0.00128706 3.3 0.0012869799999999999 3.3 0.00128708 0 0.001287 0 0.0012871 3.3 0.0012870199999999998 3.3 0.0012871199999999999 0 0.00128704 0 0.00128714 3.3 0.0012870599999999998 3.3 0.0012871599999999999 0 0.00128708 0 0.00128718 3.3 0.0012871 3.3 0.0012872 0 0.0012871199999999999 0 0.00128722 3.3 0.00128714 3.3 0.00128724 0 0.0012871599999999999 0 0.00128726 3.3 0.00128718 3.3 0.00128728 0 0.0012871999999999998 0 0.0012873 3.3 0.00128722 3.3 0.00128732 0 0.0012872399999999998 0 0.0012873399999999999 3.3 0.00128726 3.3 0.00128736 0 0.00128728 0 0.00128738 3.3 0.0012873 3.3 0.0012874 0 0.00128732 0 0.00128742 3.3 0.0012873399999999999 3.3 0.00128744 0 0.00128736 0 0.00128746 3.3 0.0012873799999999999 3.3 0.00128748 0 0.0012874 0 0.0012875 3.3 0.0012874199999999998 3.3 0.00128752 0 0.00128744 0 0.00128754 3.3 0.0012874599999999998 3.3 0.0012875599999999999 0 0.00128748 0 0.00128758 3.3 0.0012875 3.3 0.0012876 0 0.00128752 0 0.00128762 3.3 0.00128754 3.3 0.00128764 0 0.0012875599999999999 0 0.00128766 3.3 0.00128758 3.3 0.00128768 0 0.0012875999999999999 0 0.0012877 3.3 0.00128762 3.3 0.00128772 0 0.0012876399999999998 0 0.00128774 3.3 0.00128766 3.3 0.00128776 0 0.0012876799999999998 0 0.0012877799999999999 3.3 0.0012877 3.3 0.0012878 0 0.00128772 0 0.00128782 3.3 0.00128774 3.3 0.00128784 0 0.00128776 0 0.00128786 3.3 0.0012877799999999999 3.3 0.00128788 0 0.0012878 0 0.0012879 3.3 0.0012878199999999999 3.3 0.00128792 0 0.00128784 0 0.00128794 3.3 0.0012878599999999998 3.3 0.0012879599999999999 0 0.00128788 0 0.00128798 3.3 0.0012879 3.3 0.001288 0 0.00128792 0 0.00128802 3.3 0.00128794 3.3 0.00128804 0 0.0012879599999999999 0 0.00128806 3.3 0.00128798 3.3 0.00128808 0 0.0012879999999999999 0 0.0012881 3.3 0.00128802 3.3 0.00128812 0 0.0012880399999999998 0 0.00128814 3.3 0.00128806 3.3 0.00128816 0 0.0012880799999999998 0 0.0012881799999999999 3.3 0.0012881 3.3 0.0012882 0 0.00128812 0 0.00128822 3.3 0.00128814 3.3 0.00128824 0 0.00128816 0 0.00128826 3.3 0.0012881799999999999 3.3 0.00128828 0 0.0012882 0 0.0012883 3.3 0.0012882199999999999 3.3 0.00128832 0 0.00128824 0 0.00128834 3.3 0.0012882599999999998 3.3 0.00128836 0 0.00128828 0 0.00128838 3.3 0.0012882999999999998 3.3 0.0012883999999999999 0 0.00128832 0 0.00128842 3.3 0.00128834 3.3 0.00128844 0 0.00128836 0 0.00128846 3.3 0.00128838 3.3 0.00128848 0 0.0012883999999999999 0 0.0012885 3.3 0.00128842 3.3 0.00128852 0 0.0012884399999999999 0 0.00128854 3.3 0.00128846 3.3 0.00128856 0 0.0012884799999999998 0 0.0012885799999999999 3.3 0.0012885 3.3 0.0012886 0 0.0012885199999999998 0 0.0012886199999999999 3.3 0.00128854 3.3 0.00128864 0 0.00128856 0 0.00128866 3.3 0.0012885799999999999 3.3 0.00128868 0 0.0012886 0 0.0012887 3.3 0.0012886199999999999 3.3 0.00128872 0 0.00128864 0 0.00128874 3.3 0.0012886599999999998 3.3 0.00128876 0 0.00128868 0 0.00128878 3.3 0.0012886999999999998 3.3 0.0012887999999999999 0 0.00128872 0 0.00128882 3.3 0.00128874 3.3 0.00128884 0 0.00128876 0 0.00128886 3.3 0.00128878 3.3 0.00128888 0 0.0012887999999999999 0 0.0012889 3.3 0.00128882 3.3 0.00128892 0 0.0012888399999999999 0 0.00128894 3.3 0.00128886 3.3 0.00128896 0 0.0012888799999999998 0 0.00128898 3.3 0.0012889 3.3 0.001289 0 0.0012889199999999998 0 0.0012890199999999999 3.3 0.00128894 3.3 0.00128904 0 0.00128896 0 0.00128906 3.3 0.00128898 3.3 0.00128908 0 0.001289 0 0.0012891 3.3 0.0012890199999999999 3.3 0.00128912 0 0.00128904 0 0.00128914 3.3 0.0012890599999999999 3.3 0.00128916 0 0.00128908 0 0.00128918 3.3 0.0012890999999999998 3.3 0.0012892 0 0.00128912 0 0.00128922 3.3 0.0012891399999999998 3.3 0.0012892399999999999 0 0.00128916 0 0.00128926 3.3 0.00128918 3.3 0.00128928 0 0.0012892 0 0.0012893 3.3 0.00128922 3.3 0.00128932 0 0.0012892399999999999 0 0.00128934 3.3 0.00128926 3.3 0.00128936 0 0.0012892799999999999 0 0.00128938 3.3 0.0012893 3.3 0.0012894 0 0.0012893199999999998 0 0.0012894199999999999 3.3 0.00128934 3.3 0.00128944 0 0.0012893599999999998 0 0.0012894599999999999 3.3 0.00128938 3.3 0.00128948 0 0.0012894 0 0.0012895 3.3 0.0012894199999999999 3.3 0.00128952 0 0.00128944 0 0.00128954 3.3 0.0012894599999999999 3.3 0.00128956 0 0.00128948 0 0.00128958 3.3 0.0012894999999999998 3.3 0.0012896 0 0.00128952 0 0.00128962 3.3 0.0012895399999999998 3.3 0.0012896399999999999 0 0.00128956 0 0.00128966 3.3 0.00128958 3.3 0.00128968 0 0.0012896 0 0.0012897 3.3 0.00128962 3.3 0.00128972 0 0.0012896399999999999 0 0.00128974 3.3 0.00128966 3.3 0.00128976 0 0.0012896799999999999 0 0.00128978 3.3 0.0012897 3.3 0.0012898 0 0.0012897199999999998 0 0.00128982 3.3 0.00128974 3.3 0.00128984 0 0.0012897599999999998 0 0.0012898599999999999 3.3 0.00128978 3.3 0.00128988 0 0.0012898 0 0.0012899 3.3 0.00128982 3.3 0.00128992 0 0.00128984 0 0.00128994 3.3 0.0012898599999999999 3.3 0.00128996 0 0.00128988 0 0.00128998 3.3 0.0012898999999999999 3.3 0.00129 0 0.00128992 0 0.00129002 3.3 0.0012899399999999998 3.3 0.00129004 0 0.00128996 0 0.00129006 3.3 0.0012899799999999998 3.3 0.0012900799999999999 0 0.00129 0 0.0012901 3.3 0.00129002 3.3 0.00129012 0 0.00129004 0 0.00129014 3.3 0.00129006 3.3 0.00129016 0 0.0012900799999999999 0 0.00129018 3.3 0.0012901 3.3 0.0012902 0 0.0012901199999999999 0 0.00129022 3.3 0.00129014 3.3 0.00129024 0 0.0012901599999999998 0 0.0012902599999999999 3.3 0.00129018 3.3 0.00129028 0 0.0012901999999999998 0 0.0012902999999999999 3.3 0.00129022 3.3 0.00129032 0 0.00129024 0 0.00129034 3.3 0.0012902599999999999 3.3 0.00129036 0 0.00129028 0 0.00129038 3.3 0.0012902999999999999 3.3 0.0012904 0 0.00129032 0 0.00129042 3.3 0.0012903399999999998 3.3 0.00129044 0 0.00129036 0 0.00129046 3.3 0.0012903799999999998 3.3 0.0012904799999999999 0 0.0012904 0 0.0012905 3.3 0.00129042 3.3 0.00129052 0 0.00129044 0 0.00129054 3.3 0.00129046 3.3 0.00129056 0 0.0012904799999999999 0 0.00129058 3.3 0.0012905 3.3 0.0012906 0 0.0012905199999999999 0 0.00129062 3.3 0.00129054 3.3 0.00129064 0 0.0012905599999999998 0 0.00129066 3.3 0.00129058 3.3 0.00129068 0 0.0012905999999999998 0 0.0012906999999999999 3.3 0.00129062 3.3 0.00129072 0 0.00129064 0 0.00129074 3.3 0.00129066 3.3 0.00129076 0 0.00129068 0 0.00129078 3.3 0.0012906999999999999 3.3 0.0012908 0 0.00129072 0 0.00129082 3.3 0.0012907399999999999 3.3 0.00129084 0 0.00129076 0 0.00129086 3.3 0.0012907799999999998 3.3 0.00129088 0 0.0012908 0 0.0012909 3.3 0.0012908199999999998 3.3 0.0012909199999999999 0 0.00129084 0 0.00129094 3.3 0.00129086 3.3 0.00129096 0 0.00129088 0 0.00129098 3.3 0.0012909 3.3 0.001291 0 0.0012909199999999999 0 0.00129102 3.3 0.00129094 3.3 0.00129104 0 0.0012909599999999999 0 0.00129106 3.3 0.00129098 3.3 0.00129108 0 0.0012909999999999998 0 0.0012910999999999999 3.3 0.00129102 3.3 0.00129112 0 0.0012910399999999998 0 0.0012911399999999999 3.3 0.00129106 3.3 0.00129116 0 0.00129108 0 0.00129118 3.3 0.0012910999999999999 3.3 0.0012912 0 0.00129112 0 0.00129122 3.3 0.0012911399999999999 3.3 0.00129124 0 0.00129116 0 0.00129126 3.3 0.0012911799999999998 3.3 0.00129128 0 0.0012912 0 0.0012913 3.3 0.0012912199999999998 3.3 0.0012913199999999999 0 0.00129124 0 0.00129134 3.3 0.00129126 3.3 0.00129136 0 0.00129128 0 0.00129138 3.3 0.0012913 3.3 0.0012914 0 0.0012913199999999999 0 0.00129142 3.3 0.00129134 3.3 0.00129144 0 0.0012913599999999999 0 0.00129146 3.3 0.00129138 3.3 0.00129148 0 0.0012913999999999998 0 0.0012915 3.3 0.00129142 3.3 0.00129152 0 0.0012914399999999998 0 0.0012915399999999999 3.3 0.00129146 3.3 0.00129156 0 0.00129148 0 0.00129158 3.3 0.0012915 3.3 0.0012916 0 0.00129152 0 0.00129162 3.3 0.0012915399999999999 3.3 0.00129164 0 0.00129156 0 0.00129166 3.3 0.0012915799999999999 3.3 0.00129168 0 0.0012916 0 0.0012917 3.3 0.0012916199999999998 3.3 0.0012917199999999999 0 0.00129164 0 0.00129174 3.3 0.0012916599999999998 3.3 0.0012917599999999999 0 0.00129168 0 0.00129178 3.3 0.0012917 3.3 0.0012918 0 0.0012917199999999999 0 0.00129182 3.3 0.00129174 3.3 0.00129184 0 0.0012917599999999999 0 0.00129186 3.3 0.00129178 3.3 0.00129188 0 0.0012917999999999998 0 0.0012919 3.3 0.00129182 3.3 0.00129192 0 0.0012918399999999998 0 0.0012919399999999999 3.3 0.00129186 3.3 0.00129196 0 0.00129188 0 0.00129198 3.3 0.0012919 3.3 0.001292 0 0.00129192 0 0.00129202 3.3 0.0012919399999999999 3.3 0.00129204 0 0.00129196 0 0.00129206 3.3 0.0012919799999999999 3.3 0.00129208 0 0.001292 0 0.0012921 3.3 0.0012920199999999998 3.3 0.00129212 0 0.00129204 0 0.00129214 3.3 0.0012920599999999998 3.3 0.0012921599999999999 0 0.00129208 0 0.00129218 3.3 0.0012921 3.3 0.0012922 0 0.00129212 0 0.00129222 3.3 0.00129214 3.3 0.00129224 0 0.0012921599999999999 0 0.00129226 3.3 0.00129218 3.3 0.00129228 0 0.0012921999999999999 0 0.0012923 3.3 0.00129222 3.3 0.00129232 0 0.0012922399999999998 0 0.00129234 3.3 0.00129226 3.3 0.00129236 0 0.0012922799999999998 0 0.0012923799999999999 3.3 0.0012923 3.3 0.0012924 0 0.00129232 0 0.00129242 3.3 0.00129234 3.3 0.00129244 0 0.00129236 0 0.00129246 3.3 0.0012923799999999999 3.3 0.00129248 0 0.0012924 0 0.0012925 3.3 0.0012924199999999999 3.3 0.00129252 0 0.00129244 0 0.00129254 3.3 0.0012924599999999998 3.3 0.0012925599999999999 0 0.00129248 0 0.00129258 3.3 0.0012924999999999998 3.3 0.0012925999999999999 0 0.00129252 0 0.00129262 3.3 0.00129254 3.3 0.00129264 0 0.0012925599999999999 0 0.00129266 3.3 0.00129258 3.3 0.00129268 0 0.0012925999999999999 0 0.0012927 3.3 0.00129262 3.3 0.00129272 0 0.0012926399999999998 0 0.00129274 3.3 0.00129266 3.3 0.00129276 0 0.0012926799999999998 0 0.0012927799999999999 3.3 0.0012927 3.3 0.0012928 0 0.00129272 0 0.00129282 3.3 0.00129274 3.3 0.00129284 0 0.00129276 0 0.00129286 3.3 0.0012927799999999999 3.3 0.00129288 0 0.0012928 0 0.0012929 3.3 0.0012928199999999999 3.3 0.00129292 0 0.00129284 0 0.00129294 3.3 0.0012928599999999998 3.3 0.00129296 0 0.00129288 0 0.00129298 3.3 0.0012928999999999998 3.3 0.0012929999999999999 0 0.00129292 0 0.00129302 3.3 0.00129294 3.3 0.00129304 0 0.00129296 0 0.00129306 3.3 0.00129298 3.3 0.00129308 0 0.0012929999999999999 0 0.0012931 3.3 0.00129302 3.3 0.00129312 0 0.0012930399999999999 0 0.00129314 3.3 0.00129306 3.3 0.00129316 0 0.0012930799999999998 0 0.00129318 3.3 0.0012931 3.3 0.0012932 0 0.0012931199999999998 0 0.0012932199999999999 3.3 0.00129314 3.3 0.00129324 0 0.00129316 0 0.00129326 3.3 0.00129318 3.3 0.00129328 0 0.0012932 0 0.0012933 3.3 0.0012932199999999999 3.3 0.00129332 0 0.00129324 0 0.00129334 3.3 0.0012932599999999999 3.3 0.00129336 0 0.00129328 0 0.00129338 3.3 0.0012932999999999998 3.3 0.0012933999999999999 0 0.00129332 0 0.00129342 3.3 0.0012933399999999998 3.3 0.0012934399999999999 0 0.00129336 0 0.00129346 3.3 0.00129338 3.3 0.00129348 0 0.0012933999999999999 0 0.0012935 3.3 0.00129342 3.3 0.00129352 0 0.0012934399999999999 0 0.00129354 3.3 0.00129346 3.3 0.00129356 0 0.0012934799999999998 0 0.00129358 3.3 0.0012935 3.3 0.0012936 0 0.0012935199999999998 0 0.0012936199999999999 3.3 0.00129354 3.3 0.00129364 0 0.00129356 0 0.00129366 3.3 0.00129358 3.3 0.00129368 0 0.0012936 0 0.0012937 3.3 0.0012936199999999999 3.3 0.00129372 0 0.00129364 0 0.00129374 3.3 0.0012936599999999999 3.3 0.00129376 0 0.00129368 0 0.00129378 3.3 0.0012936999999999998 3.3 0.0012938 0 0.00129372 0 0.00129382 3.3 0.0012937399999999998 3.3 0.0012938399999999999 0 0.00129376 0 0.00129386 3.3 0.00129378 3.3 0.00129388 0 0.0012938 0 0.0012939 3.3 0.00129382 3.3 0.00129392 0 0.0012938399999999999 0 0.00129394 3.3 0.00129386 3.3 0.00129396 0 0.0012938799999999999 0 0.00129398 3.3 0.0012939 3.3 0.001294 0 0.0012939199999999998 0 0.00129402 3.3 0.00129394 3.3 0.00129404 0 0.0012939599999999998 0 0.0012940599999999999 3.3 0.00129398 3.3 0.00129408 0 0.001294 0 0.0012941 3.3 0.00129402 3.3 0.00129412 0 0.00129404 0 0.00129414 3.3 0.0012940599999999999 3.3 0.00129416 0 0.00129408 0 0.00129418 3.3 0.0012940999999999999 3.3 0.0012942 0 0.00129412 0 0.00129422 3.3 0.0012941399999999998 3.3 0.0012942399999999999 0 0.00129416 0 0.00129426 3.3 0.0012941799999999998 3.3 0.0012942799999999999 0 0.0012942 0 0.0012943 3.3 0.00129422 3.3 0.00129432 0 0.0012942399999999999 0 0.00129434 3.3 0.00129426 3.3 0.00129436 0 0.0012942799999999999 0 0.00129438 3.3 0.0012943 3.3 0.0012944 0 0.0012943199999999998 0 0.00129442 3.3 0.00129434 3.3 0.00129444 0 0.0012943599999999998 0 0.0012944599999999999 3.3 0.00129438 3.3 0.00129448 0 0.0012944 0 0.0012945 3.3 0.00129442 3.3 0.00129452 0 0.00129444 0 0.00129454 3.3 0.0012944599999999999 3.3 0.00129456 0 0.00129448 0 0.00129458 3.3 0.0012944999999999999 3.3 0.0012946 0 0.00129452 0 0.00129462 3.3 0.0012945399999999998 3.3 0.00129464 0 0.00129456 0 0.00129466 3.3 0.0012945799999999998 3.3 0.0012946799999999999 0 0.0012946 0 0.0012947 3.3 0.00129462 3.3 0.00129472 0 0.00129464 0 0.00129474 3.3 0.00129466 3.3 0.00129476 0 0.0012946799999999999 0 0.00129478 3.3 0.0012947 3.3 0.0012948 0 0.0012947199999999999 0 0.00129482 3.3 0.00129474 3.3 0.00129484 0 0.0012947599999999998 0 0.0012948599999999999 3.3 0.00129478 3.3 0.00129488 0 0.0012947999999999998 0 0.0012948999999999999 3.3 0.00129482 3.3 0.00129492 0 0.00129484 0 0.00129494 3.3 0.0012948599999999999 3.3 0.00129496 0 0.00129488 0 0.00129498 3.3 0.0012948999999999999 3.3 0.001295 0 0.00129492 0 0.00129502 3.3 0.0012949399999999998 3.3 0.00129504 0 0.00129496 0 0.00129506 3.3 0.0012949799999999998 3.3 0.0012950799999999999 0 0.001295 0 0.0012951 3.3 0.00129502 3.3 0.00129512 0 0.00129504 0 0.00129514 3.3 0.00129506 3.3 0.00129516 0 0.0012950799999999999 0 0.00129518 3.3 0.0012951 3.3 0.0012952 0 0.0012951199999999999 0 0.00129522 3.3 0.00129514 3.3 0.00129524 0 0.0012951599999999998 0 0.00129526 3.3 0.00129518 3.3 0.00129528 0 0.0012951999999999998 0 0.0012952999999999999 3.3 0.00129522 3.3 0.00129532 0 0.00129524 0 0.00129534 3.3 0.00129526 3.3 0.00129536 0 0.00129528 0 0.00129538 3.3 0.0012952999999999999 3.3 0.0012954 0 0.00129532 0 0.00129542 3.3 0.0012953399999999999 3.3 0.00129544 0 0.00129536 0 0.00129546 3.3 0.0012953799999999998 3.3 0.00129548 0 0.0012954 0 0.0012955 3.3 0.0012954199999999998 3.3 0.0012955199999999999 0 0.00129544 0 0.00129554 3.3 0.00129546 3.3 0.00129556 0 0.00129548 0 0.00129558 3.3 0.0012955 3.3 0.0012956 0 0.0012955199999999999 0 0.00129562 3.3 0.00129554 3.3 0.00129564 0 0.0012955599999999999 0 0.00129566 3.3 0.00129558 3.3 0.00129568 0 0.0012955999999999998 0 0.0012956999999999999 3.3 0.00129562 3.3 0.00129572 0 0.0012956399999999998 0 0.0012957399999999999 3.3 0.00129566 3.3 0.00129576 0 0.00129568 0 0.00129578 3.3 0.0012956999999999999 3.3 0.0012958 0 0.00129572 0 0.00129582 3.3 0.0012957399999999999 3.3 0.00129584 0 0.00129576 0 0.00129586 3.3 0.0012957799999999998 3.3 0.00129588 0 0.0012958 0 0.0012959 3.3 0.0012958199999999998 3.3 0.0012959199999999999 0 0.00129584 0 0.00129594 3.3 0.00129586 3.3 0.00129596 0 0.00129588 0 0.00129598 3.3 0.0012959 3.3 0.001296 0 0.0012959199999999999 0 0.00129602 3.3 0.00129594 3.3 0.00129604 0 0.0012959599999999999 0 0.00129606 3.3 0.00129598 3.3 0.00129608 0 0.0012959999999999998 0 0.0012961 3.3 0.00129602 3.3 0.00129612 0 0.0012960399999999998 0 0.0012961399999999999 3.3 0.00129606 3.3 0.00129616 0 0.00129608 0 0.00129618 3.3 0.0012961 3.3 0.0012962 0 0.00129612 0 0.00129622 3.3 0.0012961399999999999 3.3 0.00129624 0 0.00129616 0 0.00129626 3.3 0.0012961799999999999 3.3 0.00129628 0 0.0012962 0 0.0012963 3.3 0.0012962199999999998 3.3 0.00129632 0 0.00129624 0 0.00129634 3.3 0.0012962599999999998 3.3 0.0012963599999999999 0 0.00129628 0 0.00129638 3.3 0.0012963 3.3 0.0012964 0 0.00129632 0 0.00129642 3.3 0.00129634 3.3 0.00129644 0 0.0012963599999999999 0 0.00129646 3.3 0.00129638 3.3 0.00129648 0 0.0012963999999999999 0 0.0012965 3.3 0.00129642 3.3 0.00129652 0 0.0012964399999999998 0 0.0012965399999999999 3.3 0.00129646 3.3 0.00129656 0 0.0012964799999999998 0 0.0012965799999999999 3.3 0.0012965 3.3 0.0012966 0 0.00129652 0 0.00129662 3.3 0.0012965399999999999 3.3 0.00129664 0 0.00129656 0 0.00129666 3.3 0.0012965799999999999 3.3 0.00129668 0 0.0012966 0 0.0012967 3.3 0.0012966199999999998 3.3 0.00129672 0 0.00129664 0 0.00129674 3.3 0.0012966599999999998 3.3 0.0012967599999999999 0 0.00129668 0 0.00129678 3.3 0.0012967 3.3 0.0012968 0 0.00129672 0 0.00129682 3.3 0.00129674 3.3 0.00129684 0 0.0012967599999999999 0 0.00129686 3.3 0.00129678 3.3 0.00129688 0 0.0012967999999999999 0 0.0012969 3.3 0.00129682 3.3 0.00129692 0 0.0012968399999999998 0 0.00129694 3.3 0.00129686 3.3 0.00129696 0 0.0012968799999999998 0 0.0012969799999999999 3.3 0.0012969 3.3 0.001297 0 0.00129692 0 0.00129702 3.3 0.00129694 3.3 0.00129704 0 0.00129696 0 0.00129706 3.3 0.0012969799999999999 3.3 0.00129708 0 0.001297 0 0.0012971 3.3 0.0012970199999999999 3.3 0.00129712 0 0.00129704 0 0.00129714 3.3 0.0012970599999999998 3.3 0.00129716 0 0.00129708 0 0.00129718 3.3 0.0012970999999999998 3.3 0.0012971999999999999 0 0.00129712 0 0.00129722 3.3 0.00129714 3.3 0.00129724 0 0.00129716 0 0.00129726 3.3 0.00129718 3.3 0.00129728 0 0.0012971999999999999 0 0.0012973 3.3 0.00129722 3.3 0.00129732 0 0.0012972399999999999 0 0.00129734 3.3 0.00129726 3.3 0.00129736 0 0.0012972799999999998 0 0.0012973799999999999 3.3 0.0012973 3.3 0.0012974 0 0.0012973199999999998 0 0.0012974199999999999 3.3 0.00129734 3.3 0.00129744 0 0.00129736 0 0.00129746 3.3 0.0012973799999999999 3.3 0.00129748 0 0.0012974 0 0.0012975 3.3 0.0012974199999999999 3.3 0.00129752 0 0.00129744 0 0.00129754 3.3 0.0012974599999999998 3.3 0.00129756 0 0.00129748 0 0.00129758 3.3 0.0012974999999999998 3.3 0.0012975999999999999 0 0.00129752 0 0.00129762 3.3 0.00129754 3.3 0.00129764 0 0.00129756 0 0.00129766 3.3 0.00129758 3.3 0.00129768 0 0.0012975999999999999 0 0.0012977 3.3 0.00129762 3.3 0.00129772 0 0.0012976399999999999 0 0.00129774 3.3 0.00129766 3.3 0.00129776 0 0.0012976799999999998 0 0.00129778 3.3 0.0012977 3.3 0.0012978 0 0.0012977199999999998 0 0.0012978199999999999 3.3 0.00129774 3.3 0.00129784 0 0.00129776 0 0.00129786 3.3 0.00129778 3.3 0.00129788 0 0.0012978 0 0.0012979 3.3 0.0012978199999999999 3.3 0.00129792 0 0.00129784 0 0.00129794 3.3 0.0012978599999999999 3.3 0.00129796 0 0.00129788 0 0.00129798 3.3 0.0012978999999999998 3.3 0.001298 0 0.00129792 0 0.00129802 3.3 0.0012979399999999998 3.3 0.0012980399999999999 0 0.00129796 0 0.00129806 3.3 0.00129798 3.3 0.00129808 0 0.001298 0 0.0012981 3.3 0.00129802 3.3 0.00129812 0 0.0012980399999999999 0 0.00129814 3.3 0.00129806 3.3 0.00129816 0 0.0012980799999999999 0 0.00129818 3.3 0.0012981 3.3 0.0012982 0 0.0012981199999999998 0 0.0012982199999999999 3.3 0.00129814 3.3 0.00129824 0 0.0012981599999999998 0 0.0012982599999999999 3.3 0.00129818 3.3 0.00129828 0 0.0012982 0 0.0012983 3.3 0.0012982199999999999 3.3 0.00129832 0 0.00129824 0 0.00129834 3.3 0.0012982599999999999 3.3 0.00129836 0 0.00129828 0 0.00129838 3.3 0.0012982999999999998 3.3 0.0012984 0 0.00129832 0 0.00129842 3.3 0.0012983399999999998 3.3 0.0012984399999999999 0 0.00129836 0 0.00129846 3.3 0.00129838 3.3 0.00129848 0 0.0012984 0 0.0012985 3.3 0.00129842 3.3 0.00129852 0 0.0012984399999999999 0 0.00129854 3.3 0.00129846 3.3 0.00129856 0 0.0012984799999999999 0 0.00129858 3.3 0.0012985 3.3 0.0012986 0 0.0012985199999999998 0 0.00129862 3.3 0.00129854 3.3 0.00129864 0 0.0012985599999999998 0 0.0012986599999999999 3.3 0.00129858 3.3 0.00129868 0 0.0012986 0 0.0012987 3.3 0.00129862 3.3 0.00129872 0 0.00129864 0 0.00129874 3.3 0.0012986599999999999 3.3 0.00129876 0 0.00129868 0 0.00129878 3.3 0.0012986999999999999 3.3 0.0012988 0 0.00129872 0 0.00129882 3.3 0.0012987399999999998 3.3 0.0012988399999999999 0 0.00129876 0 0.00129886 3.3 0.0012987799999999998 3.3 0.0012988799999999999 0 0.0012988 0 0.0012989 3.3 0.00129882 3.3 0.00129892 0 0.0012988399999999999 0 0.00129894 3.3 0.00129886 3.3 0.00129896 0 0.0012988799999999999 0 0.00129898 3.3 0.0012989 3.3 0.001299 0 0.0012989199999999998 0 0.00129902 3.3 0.00129894 3.3 0.00129904 0 0.0012989599999999998 0 0.0012990599999999999 3.3 0.00129898 3.3 0.00129908 0 0.001299 0 0.0012991 3.3 0.00129902 3.3 0.00129912 0 0.00129904 0 0.00129914 3.3 0.0012990599999999999 3.3 0.00129916 0 0.00129908 0 0.00129918 3.3 0.0012990999999999999 3.3 0.0012992 0 0.00129912 0 0.00129922 3.3 0.0012991399999999998 3.3 0.00129924 0 0.00129916 0 0.00129926 3.3 0.0012991799999999998 3.3 0.0012992799999999999 0 0.0012992 0 0.0012993 3.3 0.00129922 3.3 0.00129932 0 0.00129924 0 0.00129934 3.3 0.00129926 3.3 0.00129936 0 0.0012992799999999999 0 0.00129938 3.3 0.0012993 3.3 0.0012994 0 0.0012993199999999999 0 0.00129942 3.3 0.00129934 3.3 0.00129944 0 0.0012993599999999998 0 0.00129946 3.3 0.00129938 3.3 0.00129948 0 0.0012993999999999998 0 0.0012994999999999999 3.3 0.00129942 3.3 0.00129952 0 0.00129944 0 0.00129954 3.3 0.00129946 3.3 0.00129956 0 0.00129948 0 0.00129958 3.3 0.0012994999999999999 3.3 0.0012996 0 0.00129952 0 0.00129962 3.3 0.0012995399999999999 3.3 0.00129964 0 0.00129956 0 0.00129966 3.3 0.0012995799999999998 3.3 0.0012996799999999999 0 0.0012996 0 0.0012997 3.3 0.0012996199999999998 3.3 0.0012997199999999999 0 0.00129964 0 0.00129974 3.3 0.00129966 3.3 0.00129976 0 0.0012996799999999999 0 0.00129978 3.3 0.0012997 3.3 0.0012998 0 0.0012997199999999999 0 0.00129982 3.3 0.00129974 3.3 0.00129984 0 0.0012997599999999998 0 0.00129986 3.3 0.00129978 3.3 0.00129988 0 0.0012997999999999998 0 0.0012998999999999999 3.3 0.00129982 3.3 0.00129992 0 0.00129984 0 0.00129994 3.3 0.00129986 3.3 0.00129996 0 0.00129988 0 0.00129998 3.3 0.0012998999999999999 3.3 0.0013 0 0.00129992 0 0.00130002 3.3 0.0012999399999999999 3.3 0.00130004 0 0.00129996 0 0.00130006 3.3 0.0012999799999999998 3.3 0.00130008 0 0.0013 0 0.0013001 3.3 0.0013000199999999998 3.3 0.0013001199999999999 0 0.00130004 0 0.00130014 3.3 0.00130006 3.3 0.00130016 0 0.00130008 0 0.00130018 3.3 0.0013001 3.3 0.0013002 0 0.0013001199999999999 0 0.00130022 3.3 0.00130014 3.3 0.00130024 0 0.0013001599999999999 0 0.00130026 3.3 0.00130018 3.3 0.00130028 0 0.0013001999999999998 0 0.0013003 3.3 0.00130022 3.3 0.00130032 0 0.0013002399999999998 0 0.0013003399999999999 3.3 0.00130026 3.3 0.00130036 0 0.00130028 0 0.00130038 3.3 0.0013003 3.3 0.0013004 0 0.00130032 0 0.00130042 3.3 0.0013003399999999999 3.3 0.00130044 0 0.00130036 0 0.00130046 3.3 0.0013003799999999999 3.3 0.00130048 0 0.0013004 0 0.0013005 3.3 0.0013004199999999998 3.3 0.0013005199999999999 0 0.00130044 0 0.00130054 3.3 0.0013004599999999998 3.3 0.0013005599999999999 0 0.00130048 0 0.00130058 3.3 0.0013005 3.3 0.0013006 0 0.0013005199999999999 0 0.00130062 3.3 0.00130054 3.3 0.00130064 0 0.0013005599999999999 0 0.00130066 3.3 0.00130058 3.3 0.00130068 0 0.0013005999999999998 0 0.0013007 3.3 0.00130062 3.3 0.00130072 0 0.0013006399999999998 0 0.0013007399999999999 3.3 0.00130066 3.3 0.00130076 0 0.00130068 0 0.00130078 3.3 0.0013007 3.3 0.0013008 0 0.00130072 0 0.00130082 3.3 0.0013007399999999999 3.3 0.00130084 0 0.00130076 0 0.00130086 3.3 0.0013007799999999999 3.3 0.00130088 0 0.0013008 0 0.0013009 3.3 0.0013008199999999998 3.3 0.00130092 0 0.00130084 0 0.00130094 3.3 0.0013008599999999998 3.3 0.0013009599999999999 0 0.00130088 0 0.00130098 3.3 0.0013009 3.3 0.001301 0 0.00130092 0 0.00130102 3.3 0.00130094 3.3 0.00130104 0 0.0013009599999999999 0 0.00130106 3.3 0.00130098 3.3 0.00130108 0 0.0013009999999999999 0 0.0013011 3.3 0.00130102 3.3 0.00130112 0 0.0013010399999999998 0 0.00130114 3.3 0.00130106 3.3 0.00130116 0 0.0013010799999999998 0 0.0013011799999999999 3.3 0.0013011 3.3 0.0013012 0 0.00130112 0 0.00130122 3.3 0.00130114 3.3 0.00130124 0 0.00130116 0 0.00130126 3.3 0.0013011799999999999 3.3 0.00130128 0 0.0013012 0 0.0013013 3.3 0.0013012199999999999 3.3 0.00130132 0 0.00130124 0 0.00130134 3.3 0.0013012599999999998 3.3 0.0013013599999999999 0 0.00130128 0 0.00130138 3.3 0.0013012999999999998 3.3 0.0013013999999999999 0 0.00130132 0 0.00130142 3.3 0.00130134 3.3 0.00130144 0 0.0013013599999999999 0 0.00130146 3.3 0.00130138 3.3 0.00130148 0 0.0013013999999999999 0 0.0013015 3.3 0.00130142 3.3 0.00130152 0 0.0013014399999999998 0 0.00130154 3.3 0.00130146 3.3 0.00130156 0 0.0013014799999999998 0 0.0013015799999999999 3.3 0.0013015 3.3 0.0013016 0 0.00130152 0 0.00130162 3.3 0.00130154 3.3 0.00130164 0 0.00130156 0 0.00130166 3.3 0.0013015799999999999 3.3 0.00130168 0 0.0013016 0 0.0013017 3.3 0.0013016199999999999 3.3 0.00130172 0 0.00130164 0 0.00130174 3.3 0.0013016599999999998 3.3 0.00130176 0 0.00130168 0 0.00130178 3.3 0.0013016999999999998 3.3 0.0013017999999999999 0 0.00130172 0 0.00130182 3.3 0.00130174 3.3 0.00130184 0 0.00130176 0 0.00130186 3.3 0.00130178 3.3 0.00130188 0 0.0013017999999999999 0 0.0013019 3.3 0.00130182 3.3 0.00130192 0 0.0013018399999999999 0 0.00130194 3.3 0.00130186 3.3 0.00130196 0 0.0013018799999999998 0 0.0013019799999999999 3.3 0.0013019 3.3 0.001302 0 0.0013019199999999998 0 0.0013020199999999999 3.3 0.00130194 3.3 0.00130204 0 0.00130196 0 0.00130206 3.3 0.0013019799999999999 3.3 0.00130208 0 0.001302 0 0.0013021 3.3 0.0013020199999999999 3.3 0.00130212 0 0.00130204 0 0.00130214 3.3 0.0013020599999999998 3.3 0.00130216 0 0.00130208 0 0.00130218 3.3 0.0013020999999999998 3.3 0.0013021999999999999 0 0.00130212 0 0.00130222 3.3 0.00130214 3.3 0.00130224 0 0.00130216 0 0.00130226 3.3 0.00130218 3.3 0.00130228 0 0.0013021999999999999 0 0.0013023 3.3 0.00130222 3.3 0.00130232 0 0.0013022399999999999 0 0.00130234 3.3 0.00130226 3.3 0.00130236 0 0.0013022799999999998 0 0.00130238 3.3 0.0013023 3.3 0.0013024 0 0.0013023199999999998 0 0.0013024199999999999 3.3 0.00130234 3.3 0.00130244 0 0.00130236 0 0.00130246 3.3 0.00130238 3.3 0.00130248 0 0.0013024 0 0.0013025 3.3 0.0013024199999999999 3.3 0.00130252 0 0.00130244 0 0.00130254 3.3 0.0013024599999999999 3.3 0.00130256 0 0.00130248 0 0.00130258 3.3 0.0013024999999999998 3.3 0.0013026 0 0.00130252 0 0.00130262 3.3 0.0013025399999999998 3.3 0.0013026399999999999 0 0.00130256 0 0.00130266 3.3 0.00130258 3.3 0.00130268 0 0.0013026 0 0.0013027 3.3 0.00130262 3.3 0.00130272 0 0.0013026399999999999 0 0.00130274 3.3 0.00130266 3.3 0.00130276 0 0.0013026799999999999 0 0.00130278 3.3 0.0013027 3.3 0.0013028 0 0.0013027199999999998 0 0.0013028199999999999 3.3 0.00130274 3.3 0.00130284 0 0.0013027599999999998 0 0.0013028599999999999 3.3 0.00130278 3.3 0.00130288 0 0.0013028 0 0.0013029 3.3 0.0013028199999999999 3.3 0.00130292 0 0.00130284 0 0.00130294 3.3 0.0013028599999999999 3.3 0.00130296 0 0.00130288 0 0.00130298 3.3 0.0013028999999999998 3.3 0.001303 0 0.00130292 0 0.00130302 3.3 0.0013029399999999998 3.3 0.0013030399999999999 0 0.00130296 0 0.00130306 3.3 0.00130298 3.3 0.00130308 0 0.001303 0 0.0013031 3.3 0.00130302 3.3 0.00130312 0 0.0013030399999999999 0 0.00130314 3.3 0.00130306 3.3 0.00130316 0 0.0013030799999999999 0 0.00130318 3.3 0.0013031 3.3 0.0013032 0 0.0013031199999999998 0 0.00130322 3.3 0.00130314 3.3 0.00130324 0 0.0013031599999999998 0 0.0013032599999999999 3.3 0.00130318 3.3 0.00130328 0 0.0013032 0 0.0013033 3.3 0.00130322 3.3 0.00130332 0 0.00130324 0 0.00130334 3.3 0.0013032599999999999 3.3 0.00130336 0 0.00130328 0 0.00130338 3.3 0.0013032999999999999 3.3 0.0013034 0 0.00130332 0 0.00130342 3.3 0.0013033399999999998 3.3 0.00130344 0 0.00130336 0 0.00130346 3.3 0.0013033799999999998 3.3 0.0013034799999999999 0 0.0013034 0 0.0013035 3.3 0.00130342 3.3 0.00130352 0 0.00130344 0 0.00130354 3.3 0.00130346 3.3 0.00130356 0 0.0013034799999999999 0 0.00130358 3.3 0.0013035 3.3 0.0013036 0 0.0013035199999999999 0 0.00130362 3.3 0.00130354 3.3 0.00130364 0 0.0013035599999999998 0 0.0013036599999999999 3.3 0.00130358 3.3 0.00130368 0 0.0013035999999999998 0 0.0013036999999999999 3.3 0.00130362 3.3 0.00130372 0 0.00130364 0 0.00130374 3.3 0.0013036599999999999 3.3 0.00130376 0 0.00130368 0 0.00130378 3.3 0.0013036999999999999 3.3 0.0013038 0 0.00130372 0 0.00130382 3.3 0.0013037399999999998 3.3 0.00130384 0 0.00130376 0 0.00130386 3.3 0.0013037799999999998 3.3 0.0013038799999999999 0 0.0013038 0 0.0013039 3.3 0.00130382 3.3 0.00130392 0 0.00130384 0 0.00130394 3.3 0.00130386 3.3 0.00130396 0 0.0013038799999999999 0 0.00130398 3.3 0.0013039 3.3 0.001304 0 0.0013039199999999999 0 0.00130402 3.3 0.00130394 3.3 0.00130404 0 0.0013039599999999998 0 0.00130406 3.3 0.00130398 3.3 0.00130408 0 0.0013039999999999998 0 0.0013040999999999999 3.3 0.00130402 3.3 0.00130412 0 0.00130404 0 0.00130414 3.3 0.00130406 3.3 0.00130416 0 0.00130408 0 0.00130418 3.3 0.0013040999999999999 3.3 0.0013042 0 0.00130412 0 0.00130422 3.3 0.0013041399999999999 3.3 0.00130424 0 0.00130416 0 0.00130426 3.3 0.0013041799999999998 3.3 0.00130428 0 0.0013042 0 0.0013043 3.3 0.0013042199999999998 3.3 0.0013043199999999999 0 0.00130424 0 0.00130434 3.3 0.00130426 3.3 0.00130436 0 0.00130428 0 0.00130438 3.3 0.0013043 3.3 0.0013044 0 0.0013043199999999999 0 0.00130442 3.3 0.00130434 3.3 0.00130444 0 0.0013043599999999999 0 0.00130446 3.3 0.00130438 3.3 0.00130448 0 0.0013043999999999998 0 0.0013044999999999999 3.3 0.00130442 3.3 0.00130452 0 0.0013044399999999998 0 0.0013045399999999999 3.3 0.00130446 3.3 0.00130456 0 0.00130448 0 0.00130458 3.3 0.0013044999999999999 3.3 0.0013046 0 0.00130452 0 0.00130462 3.3 0.0013045399999999999 3.3 0.00130464 0 0.00130456 0 0.00130466 3.3 0.0013045799999999998 3.3 0.00130468 0 0.0013046 0 0.0013047 3.3 0.0013046199999999998 3.3 0.0013047199999999999 0 0.00130464 0 0.00130474 3.3 0.00130466 3.3 0.00130476 0 0.00130468 0 0.00130478 3.3 0.0013047 3.3 0.0013048 0 0.0013047199999999999 0 0.00130482 3.3 0.00130474 3.3 0.00130484 0 0.0013047599999999999 0 0.00130486 3.3 0.00130478 3.3 0.00130488 0 0.0013047999999999998 0 0.0013049 3.3 0.00130482 3.3 0.00130492 0 0.0013048399999999998 0 0.0013049399999999999 3.3 0.00130486 3.3 0.00130496 0 0.00130488 0 0.00130498 3.3 0.0013049 3.3 0.001305 0 0.00130492 0 0.00130502 3.3 0.0013049399999999999 3.3 0.00130504 0 0.00130496 0 0.00130506 3.3 0.0013049799999999999 3.3 0.00130508 0 0.001305 0 0.0013051 3.3 0.0013050199999999998 3.3 0.0013051199999999999 0 0.00130504 0 0.00130514 3.3 0.0013050599999999998 3.3 0.0013051599999999999 0 0.00130508 0 0.00130518 3.3 0.0013051 3.3 0.0013052 0 0.0013051199999999999 0 0.00130522 3.3 0.00130514 3.3 0.00130524 0 0.0013051599999999999 0 0.00130526 3.3 0.00130518 3.3 0.00130528 0 0.0013051999999999998 0 0.0013053 3.3 0.00130522 3.3 0.00130532 0 0.0013052399999999998 0 0.0013053399999999999 3.3 0.00130526 3.3 0.00130536 0 0.00130528 0 0.00130538 3.3 0.0013053 3.3 0.0013054 0 0.00130532 0 0.00130542 3.3 0.0013053399999999999 3.3 0.00130544 0 0.00130536 0 0.00130546 3.3 0.0013053799999999999 3.3 0.00130548 0 0.0013054 0 0.0013055 3.3 0.0013054199999999998 3.3 0.00130552 0 0.00130544 0 0.00130554 3.3 0.0013054599999999998 3.3 0.0013055599999999999 0 0.00130548 0 0.00130558 3.3 0.0013055 3.3 0.0013056 0 0.00130552 0 0.00130562 3.3 0.00130554 3.3 0.00130564 0 0.0013055599999999999 0 0.00130566 3.3 0.00130558 3.3 0.00130568 0 0.0013055999999999999 0 0.0013057 3.3 0.00130562 3.3 0.00130572 0 0.0013056399999999998 0 0.00130574 3.3 0.00130566 3.3 0.00130576 0 0.0013056799999999998 0 0.0013057799999999999 3.3 0.0013057 3.3 0.0013058 0 0.00130572 0 0.00130582 3.3 0.00130574 3.3 0.00130584 0 0.00130576 0 0.00130586 3.3 0.0013057799999999999 3.3 0.00130588 0 0.0013058 0 0.0013059 3.3 0.0013058199999999999 3.3 0.00130592 0 0.00130584 0 0.00130594 3.3 0.0013058599999999998 3.3 0.0013059599999999999 0 0.00130588 0 0.00130598 3.3 0.0013058999999999998 3.3 0.0013059999999999999 0 0.00130592 0 0.00130602 3.3 0.00130594 3.3 0.00130604 0 0.0013059599999999999 0 0.00130606 3.3 0.00130598 3.3 0.00130608 0 0.0013059999999999999 0 0.0013061 3.3 0.00130602 3.3 0.00130612 0 0.0013060399999999998 0 0.00130614 3.3 0.00130606 3.3 0.00130616 0 0.0013060799999999998 0 0.0013061799999999999 3.3 0.0013061 3.3 0.0013062 0 0.00130612 0 0.00130622 3.3 0.00130614 3.3 0.00130624 0 0.00130616 0 0.00130626 3.3 0.0013061799999999999 3.3 0.00130628 0 0.0013062 0 0.0013063 3.3 0.0013062199999999999 3.3 0.00130632 0 0.00130624 0 0.00130634 3.3 0.0013062599999999998 3.3 0.00130636 0 0.00130628 0 0.00130638 3.3 0.0013062999999999998 3.3 0.0013063999999999999 0 0.00130632 0 0.00130642 3.3 0.00130634 3.3 0.00130644 0 0.00130636 0 0.00130646 3.3 0.00130638 3.3 0.00130648 0 0.0013063999999999999 0 0.0013065 3.3 0.00130642 3.3 0.00130652 0 0.0013064399999999999 0 0.00130654 3.3 0.00130646 3.3 0.00130656 0 0.0013064799999999998 0 0.00130658 3.3 0.0013065 3.3 0.0013066 0 0.0013065199999999998 0 0.0013066199999999999 3.3 0.00130654 3.3 0.00130664 0 0.00130656 0 0.00130666 3.3 0.00130658 3.3 0.00130668 0 0.0013066 0 0.0013067 3.3 0.0013066199999999999 3.3 0.00130672 0 0.00130664 0 0.00130674 3.3 0.0013066599999999999 3.3 0.00130676 0 0.00130668 0 0.00130678 3.3 0.0013066999999999998 3.3 0.0013067999999999999 0 0.00130672 0 0.00130682 3.3 0.0013067399999999998 3.3 0.0013068399999999999 0 0.00130676 0 0.00130686 3.3 0.00130678 3.3 0.00130688 0 0.0013067999999999999 0 0.0013069 3.3 0.00130682 3.3 0.00130692 0 0.0013068399999999999 0 0.00130694 3.3 0.00130686 3.3 0.00130696 0 0.0013068799999999998 0 0.00130698 3.3 0.0013069 3.3 0.001307 0 0.0013069199999999998 0 0.0013070199999999999 3.3 0.00130694 3.3 0.00130704 0 0.00130696 0 0.00130706 3.3 0.00130698 3.3 0.00130708 0 0.001307 0 0.0013071 3.3 0.0013070199999999999 3.3 0.00130712 0 0.00130704 0 0.00130714 3.3 0.0013070599999999999 3.3 0.00130716 0 0.00130708 0 0.00130718 3.3 0.0013070999999999998 3.3 0.0013072 0 0.00130712 0 0.00130722 3.3 0.0013071399999999998 3.3 0.0013072399999999999 0 0.00130716 0 0.00130726 3.3 0.00130718 3.3 0.00130728 0 0.0013072 0 0.0013073 3.3 0.00130722 3.3 0.00130732 0 0.0013072399999999999 0 0.00130734 3.3 0.00130726 3.3 0.00130736 0 0.0013072799999999999 0 0.00130738 3.3 0.0013073 3.3 0.0013074 0 0.0013073199999999998 0 0.00130742 3.3 0.00130734 3.3 0.00130744 0 0.0013073599999999998 0 0.0013074599999999999 3.3 0.00130738 3.3 0.00130748 0 0.0013074 0 0.0013075 3.3 0.00130742 3.3 0.00130752 0 0.00130744 0 0.00130754 3.3 0.0013074599999999999 3.3 0.00130756 0 0.00130748 0 0.00130758 3.3 0.0013074999999999999 3.3 0.0013076 0 0.00130752 0 0.00130762 3.3 0.0013075399999999998 3.3 0.0013076399999999999 0 0.00130756 0 0.00130766 3.3 0.0013075799999999998 3.3 0.0013076799999999999 0 0.0013076 0 0.0013077 3.3 0.00130762 3.3 0.00130772 0 0.0013076399999999999 0 0.00130774 3.3 0.00130766 3.3 0.00130776 0 0.0013076799999999999 0 0.00130778 3.3 0.0013077 3.3 0.0013078 0 0.0013077199999999998 0 0.00130782 3.3 0.00130774 3.3 0.00130784 0 0.0013077599999999998 0 0.0013078599999999999 3.3 0.00130778 3.3 0.00130788 0 0.0013078 0 0.0013079 3.3 0.00130782 3.3 0.00130792 0 0.00130784 0 0.00130794 3.3 0.0013078599999999999 3.3 0.00130796 0 0.00130788 0 0.00130798 3.3 0.0013078999999999999 3.3 0.001308 0 0.00130792 0 0.00130802 3.3 0.0013079399999999998 3.3 0.00130804 0 0.00130796 0 0.00130806 3.3 0.0013079799999999998 3.3 0.0013080799999999999 0 0.001308 0 0.0013081 3.3 0.00130802 3.3 0.00130812 0 0.00130804 0 0.00130814 3.3 0.00130806 3.3 0.00130816 0 0.0013080799999999999 0 0.00130818 3.3 0.0013081 3.3 0.0013082 0 0.0013081199999999999 0 0.00130822 3.3 0.00130814 3.3 0.00130824 0 0.0013081599999999998 0 0.00130826 3.3 0.00130818 3.3 0.00130828 0 0.0013081999999999998 0 0.0013082999999999999 3.3 0.00130822 3.3 0.00130832 0 0.00130824 0 0.00130834 3.3 0.00130826 3.3 0.00130836 0 0.00130828 0 0.00130838 3.3 0.0013082999999999999 3.3 0.0013084 0 0.00130832 0 0.00130842 3.3 0.0013083399999999999 3.3 0.00130844 0 0.00130836 0 0.00130846 3.3 0.0013083799999999998 3.3 0.0013084799999999999 0 0.0013084 0 0.0013085 3.3 0.0013084199999999998 3.3 0.0013085199999999999 0 0.00130844 0 0.00130854 3.3 0.00130846 3.3 0.00130856 0 0.0013084799999999999 0 0.00130858 3.3 0.0013085 3.3 0.0013086 0 0.0013085199999999999 0 0.00130862 3.3 0.00130854 3.3 0.00130864 0 0.0013085599999999998 0 0.00130866 3.3 0.00130858 3.3 0.00130868 0 0.0013085999999999998 0 0.0013086999999999999 3.3 0.00130862 3.3 0.00130872 0 0.00130864 0 0.00130874 3.3 0.00130866 3.3 0.00130876 0 0.00130868 0 0.00130878 3.3 0.0013086999999999999 3.3 0.0013088 0 0.00130872 0 0.00130882 3.3 0.0013087399999999999 3.3 0.00130884 0 0.00130876 0 0.00130886 3.3 0.0013087799999999998 3.3 0.00130888 0 0.0013088 0 0.0013089 3.3 0.0013088199999999998 3.3 0.0013089199999999999 0 0.00130884 0 0.00130894 3.3 0.00130886 3.3 0.00130896 0 0.00130888 0 0.00130898 3.3 0.0013089 3.3 0.001309 0 0.0013089199999999999 0 0.00130902 3.3 0.00130894 3.3 0.00130904 0 0.0013089599999999999 0 0.00130906 3.3 0.00130898 3.3 0.00130908 0 0.0013089999999999998 0 0.0013090999999999999 3.3 0.00130902 3.3 0.00130912 0 0.0013090399999999998 0 0.0013091399999999999 3.3 0.00130906 3.3 0.00130916 0 0.00130908 0 0.00130918 3.3 0.0013090999999999999 3.3 0.0013092 0 0.00130912 0 0.00130922 3.3 0.0013091399999999999 3.3 0.00130924 0 0.00130916 0 0.00130926 3.3 0.0013091799999999998 3.3 0.00130928 0 0.0013092 0 0.0013093 3.3 0.0013092199999999998 3.3 0.0013093199999999999 0 0.00130924 0 0.00130934 3.3 0.00130926 3.3 0.00130936 0 0.00130928 0 0.00130938 3.3 0.0013093 3.3 0.0013094 0 0.0013093199999999999 0 0.00130942 3.3 0.00130934 3.3 0.00130944 0 0.0013093599999999999 0 0.00130946 3.3 0.00130938 3.3 0.00130948 0 0.0013093999999999998 0 0.0013095 3.3 0.00130942 3.3 0.00130952 0 0.0013094399999999998 0 0.0013095399999999999 3.3 0.00130946 3.3 0.00130956 0 0.00130948 0 0.00130958 3.3 0.0013095 3.3 0.0013096 0 0.00130952 0 0.00130962 3.3 0.0013095399999999999 3.3 0.00130964 0 0.00130956 0 0.00130966 3.3 0.0013095799999999999 3.3 0.00130968 0 0.0013096 0 0.0013097 3.3 0.0013096199999999998 3.3 0.00130972 0 0.00130964 0 0.00130974 3.3 0.0013096599999999998 3.3 0.0013097599999999999 0 0.00130968 0 0.00130978 3.3 0.0013097 3.3 0.0013098 0 0.00130972 0 0.00130982 3.3 0.00130974 3.3 0.00130984 0 0.0013097599999999999 0 0.00130986 3.3 0.00130978 3.3 0.00130988 0 0.0013097999999999999 0 0.0013099 3.3 0.00130982 3.3 0.00130992 0 0.0013098399999999998 0 0.0013099399999999999 3.3 0.00130986 3.3 0.00130996 0 0.0013098799999999998 0 0.0013099799999999999 3.3 0.0013099 3.3 0.00131 0 0.00130992 0 0.00131002 3.3 0.0013099399999999999 3.3 0.00131004 0 0.00130996 0 0.00131006 3.3 0.0013099799999999999 3.3 0.00131008 0 0.00131 0 0.0013101 3.3 0.0013100199999999998 3.3 0.00131012 0 0.00131004 0 0.00131014 3.3 0.0013100599999999998 3.3 0.0013101599999999999 0 0.00131008 0 0.00131018 3.3 0.0013101 3.3 0.0013102 0 0.00131012 0 0.00131022 3.3 0.00131014 3.3 0.00131024 0 0.0013101599999999999 0 0.00131026 3.3 0.00131018 3.3 0.00131028 0 0.0013101999999999999 0 0.0013103 3.3 0.00131022 3.3 0.00131032 0 0.0013102399999999998 0 0.00131034 3.3 0.00131026 3.3 0.00131036 0 0.0013102799999999998 0 0.0013103799999999999 3.3 0.0013103 3.3 0.0013104 0 0.00131032 0 0.00131042 3.3 0.00131034 3.3 0.00131044 0 0.00131036 0 0.00131046 3.3 0.0013103799999999999 3.3 0.00131048 0 0.0013104 0 0.0013105 3.3 0.0013104199999999999 3.3 0.00131052 0 0.00131044 0 0.00131054 3.3 0.0013104599999999998 3.3 0.00131056 0 0.00131048 0 0.00131058 3.3 0.0013104999999999998 3.3 0.0013105999999999999 0 0.00131052 0 0.00131062 3.3 0.00131054 3.3 0.00131064 0 0.00131056 0 0.00131066 3.3 0.00131058 3.3 0.00131068 0 0.0013105999999999999 0 0.0013107 3.3 0.00131062 3.3 0.00131072 0 0.0013106399999999999 0 0.00131074 3.3 0.00131066 3.3 0.00131076 0 0.0013106799999999998 0 0.0013107799999999999 3.3 0.0013107 3.3 0.0013108 0 0.0013107199999999998 0 0.0013108199999999999 3.3 0.00131074 3.3 0.00131084 0 0.00131076 0 0.00131086 3.3 0.0013107799999999999 3.3 0.00131088 0 0.0013108 0 0.0013109 3.3 0.0013108199999999999 3.3 0.00131092 0 0.00131084 0 0.00131094 3.3 0.0013108599999999998 3.3 0.00131096 0 0.00131088 0 0.00131098 3.3 0.0013108999999999998 3.3 0.0013109999999999999 0 0.00131092 0 0.00131102 3.3 0.00131094 3.3 0.00131104 0 0.00131096 0 0.00131106 3.3 0.00131098 3.3 0.00131108 0 0.0013109999999999999 0 0.0013111 3.3 0.00131102 3.3 0.00131112 0 0.0013110399999999999 0 0.00131114 3.3 0.00131106 3.3 0.00131116 0 0.0013110799999999998 0 0.00131118 3.3 0.0013111 3.3 0.0013112 0 0.0013111199999999998 0 0.0013112199999999999 3.3 0.00131114 3.3 0.00131124 0 0.00131116 0 0.00131126 3.3 0.00131118 3.3 0.00131128 0 0.0013112 0 0.0013113 3.3 0.0013112199999999999 3.3 0.00131132 0 0.00131124 0 0.00131134 3.3 0.0013112599999999999 3.3 0.00131136 0 0.00131128 0 0.00131138 3.3 0.0013112999999999998 3.3 0.0013114 0 0.00131132 0 0.00131142 3.3 0.0013113399999999998 3.3 0.0013114399999999999 0 0.00131136 0 0.00131146 3.3 0.00131138 3.3 0.00131148 0 0.0013114 0 0.0013115 3.3 0.00131142 3.3 0.00131152 0 0.0013114399999999999 0 0.00131154 3.3 0.00131146 3.3 0.00131156 0 0.0013114799999999999 0 0.00131158 3.3 0.0013115 3.3 0.0013116 0 0.0013115199999999998 0 0.0013116199999999999 3.3 0.00131154 3.3 0.00131164 0 0.0013115599999999998 0 0.0013116599999999999 3.3 0.00131158 3.3 0.00131168 0 0.0013116 0 0.0013117 3.3 0.0013116199999999999 3.3 0.00131172 0 0.00131164 0 0.00131174 3.3 0.0013116599999999999 3.3 0.00131176 0 0.00131168 0 0.00131178 3.3 0.0013116999999999998 3.3 0.0013118 0 0.00131172 0 0.00131182 3.3 0.0013117399999999998 3.3 0.0013118399999999999 0 0.00131176 0 0.00131186 3.3 0.00131178 3.3 0.00131188 0 0.0013118 0 0.0013119 3.3 0.00131182 3.3 0.00131192 0 0.0013118399999999999 0 0.00131194 3.3 0.00131186 3.3 0.00131196 0 0.0013118799999999999 0 0.00131198 3.3 0.0013119 3.3 0.001312 0 0.0013119199999999998 0 0.00131202 3.3 0.00131194 3.3 0.00131204 0 0.0013119599999999998 0 0.0013120599999999999 3.3 0.00131198 3.3 0.00131208 0 0.001312 0 0.0013121 3.3 0.00131202 3.3 0.00131212 0 0.00131204 0 0.00131214 3.3 0.0013120599999999999 3.3 0.00131216 0 0.00131208 0 0.00131218 3.3 0.0013120999999999999 3.3 0.0013122 0 0.00131212 0 0.00131222 3.3 0.0013121399999999998 3.3 0.0013122399999999999 0 0.00131216 0 0.00131226 3.3 0.0013121799999999998 3.3 0.0013122799999999999 0 0.0013122 0 0.0013123 3.3 0.00131222 3.3 0.00131232 0 0.0013122399999999999 0 0.00131234 3.3 0.00131226 3.3 0.00131236 0 0.0013122799999999999 0 0.00131238 3.3 0.0013123 3.3 0.0013124 0 0.0013123199999999998 0 0.00131242 3.3 0.00131234 3.3 0.00131244 0 0.0013123599999999998 0 0.0013124599999999999 3.3 0.00131238 3.3 0.00131248 0 0.0013124 0 0.0013125 3.3 0.00131242 3.3 0.00131252 0 0.00131244 0 0.00131254 3.3 0.0013124599999999999 3.3 0.00131256 0 0.00131248 0 0.00131258 3.3 0.0013124999999999999 3.3 0.0013126 0 0.00131252 0 0.00131262 3.3 0.0013125399999999998 3.3 0.00131264 0 0.00131256 0 0.00131266 3.3 0.0013125799999999998 3.3 0.0013126799999999999 0 0.0013126 0 0.0013127 3.3 0.00131262 3.3 0.00131272 0 0.00131264 0 0.00131274 3.3 0.00131266 3.3 0.00131276 0 0.0013126799999999999 0 0.00131278 3.3 0.0013127 3.3 0.0013128 0 0.0013127199999999999 0 0.00131282 3.3 0.00131274 3.3 0.00131284 0 0.0013127599999999998 0 0.00131286 3.3 0.00131278 3.3 0.00131288 0 0.0013127999999999998 0 0.0013128999999999999 3.3 0.00131282 3.3 0.00131292 0 0.00131284 0 0.00131294 3.3 0.00131286 3.3 0.00131296 0 0.00131288 0 0.00131298 3.3 0.0013128999999999999 3.3 0.001313 0 0.00131292 0 0.00131302 3.3 0.0013129399999999999 3.3 0.00131304 0 0.00131296 0 0.00131306 3.3 0.0013129799999999998 3.3 0.0013130799999999999 0 0.001313 0 0.0013131 3.3 0.0013130199999999998 3.3 0.0013131199999999999 0 0.00131304 0 0.00131314 3.3 0.00131306 3.3 0.00131316 0 0.0013130799999999999 0 0.00131318 3.3 0.0013131 3.3 0.0013132 0 0.0013131199999999999 0 0.00131322 3.3 0.00131314 3.3 0.00131324 0 0.0013131599999999998 0 0.00131326 3.3 0.00131318 3.3 0.00131328 0 0.0013131999999999998 0 0.0013132999999999999 3.3 0.00131322 3.3 0.00131332 0 0.00131324 0 0.00131334 3.3 0.00131326 3.3 0.00131336 0 0.00131328 0 0.00131338 3.3 0.0013132999999999999 3.3 0.0013134 0 0.00131332 0 0.00131342 3.3 0.0013133399999999999 3.3 0.00131344 0 0.00131336 0 0.00131346 3.3 0.0013133799999999998 3.3 0.00131348 0 0.0013134 0 0.0013135 3.3 0.0013134199999999998 3.3 0.0013135199999999999 0 0.00131344 0 0.00131354 3.3 0.00131346 3.3 0.00131356 0 0.00131348 0 0.00131358 3.3 0.0013135 3.3 0.0013136 0 0.0013135199999999999 0 0.00131362 3.3 0.00131354 3.3 0.00131364 0 0.0013135599999999999 0 0.00131366 3.3 0.00131358 3.3 0.00131368 0 0.0013135999999999998 0 0.0013137 3.3 0.00131362 3.3 0.00131372 0 0.0013136399999999998 0 0.0013137399999999999 3.3 0.00131366 3.3 0.00131376 0 0.00131368 0 0.00131378 3.3 0.0013137 3.3 0.0013138 0 0.00131372 0 0.00131382 3.3 0.0013137399999999999 3.3 0.00131384 0 0.00131376 0 0.00131386 3.3 0.0013137799999999999 3.3 0.00131388 0 0.0013138 0 0.0013139 3.3 0.0013138199999999998 3.3 0.0013139199999999999 0 0.00131384 0 0.00131394 3.3 0.0013138599999999998 3.3 0.0013139599999999999 0 0.00131388 0 0.00131398 3.3 0.0013139 3.3 0.001314 0 0.0013139199999999999 0 0.00131402 3.3 0.00131394 3.3 0.00131404 0 0.0013139599999999999 0 0.00131406 3.3 0.00131398 3.3 0.00131408 0 0.0013139999999999998 0 0.0013141 3.3 0.00131402 3.3 0.00131412 0 0.0013140399999999998 0 0.0013141399999999999 3.3 0.00131406 3.3 0.00131416 0 0.00131408 0 0.00131418 3.3 0.0013141 3.3 0.0013142 0 0.00131412 0 0.00131422 3.3 0.0013141399999999999 3.3 0.00131424 0 0.00131416 0 0.00131426 3.3 0.0013141799999999999 3.3 0.00131428 0 0.0013142 0 0.0013143 3.3 0.0013142199999999998 3.3 0.00131432 0 0.00131424 0 0.00131434 3.3 0.0013142599999999998 3.3 0.0013143599999999999 0 0.00131428 0 0.00131438 3.3 0.0013143 3.3 0.0013144 0 0.00131432 0 0.00131442 3.3 0.00131434 3.3 0.00131444 0 0.0013143599999999999 0 0.00131446 3.3 0.00131438 3.3 0.00131448 0 0.0013143999999999999 0 0.0013145 3.3 0.00131442 3.3 0.00131452 0 0.0013144399999999998 0 0.00131454 3.3 0.00131446 3.3 0.00131456 0 0.0013144799999999998 0 0.0013145799999999999 3.3 0.0013145 3.3 0.0013146 0 0.00131452 0 0.00131462 3.3 0.00131454 3.3 0.00131464 0 0.00131456 0 0.00131466 3.3 0.0013145799999999999 3.3 0.00131468 0 0.0013146 0 0.0013147 3.3 0.0013146199999999999 3.3 0.00131472 0 0.00131464 0 0.00131474 3.3 0.0013146599999999998 3.3 0.0013147599999999999 0 0.00131468 0 0.00131478 3.3 0.0013146999999999998 3.3 0.0013147999999999999 0 0.00131472 0 0.00131482 3.3 0.00131474 3.3 0.00131484 0 0.0013147599999999999 0 0.00131486 3.3 0.00131478 3.3 0.00131488 0 0.0013147999999999999 0 0.0013149 3.3 0.00131482 3.3 0.00131492 0 0.0013148399999999998 0 0.00131494 3.3 0.00131486 3.3 0.00131496 0 0.0013148799999999998 0 0.0013149799999999999 3.3 0.0013149 3.3 0.001315 0 0.00131492 0 0.00131502 3.3 0.00131494 3.3 0.00131504 0 0.00131496 0 0.00131506 3.3 0.0013149799999999999 3.3 0.00131508 0 0.001315 0 0.0013151 3.3 0.0013150199999999999 3.3 0.00131512 0 0.00131504 0 0.00131514 3.3 0.0013150599999999998 3.3 0.00131516 0 0.00131508 0 0.00131518 3.3 0.0013150999999999998 3.3 0.0013151999999999999 0 0.00131512 0 0.00131522 3.3 0.00131514 3.3 0.00131524 0 0.00131516 0 0.00131526 3.3 0.00131518 3.3 0.00131528 0 0.0013151999999999999 0 0.0013153 3.3 0.00131522 3.3 0.00131532 0 0.0013152399999999999 0 0.00131534 3.3 0.00131526 3.3 0.00131536 0 0.0013152799999999998 0 0.0013153799999999999 3.3 0.0013153 3.3 0.0013154 0 0.0013153199999999998 0 0.0013154199999999999 3.3 0.00131534 3.3 0.00131544 0 0.00131536 0 0.00131546 3.3 0.0013153799999999999 3.3 0.00131548 0 0.0013154 0 0.0013155 3.3 0.0013154199999999999 3.3 0.00131552 0 0.00131544 0 0.00131554 3.3 0.0013154599999999998 3.3 0.00131556 0 0.00131548 0 0.00131558 3.3 0.0013154999999999998 3.3 0.0013155999999999999 0 0.00131552 0 0.00131562 3.3 0.0013155399999999998 3.3 0.0013156399999999999 0 0.00131556 0 0.00131566 3.3 0.00131558 3.3 0.00131568 0 0.0013155999999999999 0 0.0013157 3.3 0.00131562 3.3 0.00131572 0 0.0013156399999999999 0 0.00131574 3.3 0.00131566 3.3 0.00131576 0 0.0013156799999999998 0 0.00131578 3.3 0.0013157 3.3 0.0013158 0 0.0013157199999999998 0 0.0013158199999999999 3.3 0.00131574 3.3 0.00131584 0 0.00131576 0 0.00131586 3.3 0.00131578 3.3 0.00131588 0 0.0013158 0 0.0013159 3.3 0.0013158199999999999 3.3 0.00131592 0 0.00131584 0 0.00131594 3.3 0.0013158599999999999 3.3 0.00131596 0 0.00131588 0 0.00131598 3.3 0.0013158999999999998 3.3 0.001316 0 0.00131592 0 0.00131602 3.3 0.0013159399999999998 3.3 0.0013160399999999999 0 0.00131596 0 0.00131606 3.3 0.00131598 3.3 0.00131608 0 0.001316 0 0.0013161 3.3 0.00131602 3.3 0.00131612 0 0.0013160399999999999 0 0.00131614 3.3 0.00131606 3.3 0.00131616 0 0.0013160799999999999 0 0.00131618 3.3 0.0013161 3.3 0.0013162 0 0.0013161199999999998 0 0.0013162199999999999 3.3 0.00131614 3.3 0.00131624 0 0.0013161599999999998 0 0.0013162599999999999 3.3 0.00131618 3.3 0.00131628 0 0.0013162 0 0.0013163 3.3 0.0013162199999999999 3.3 0.00131632 0 0.00131624 0 0.00131634 3.3 0.0013162599999999999 3.3 0.00131636 0 0.00131628 0 0.00131638 3.3 0.0013162999999999998 3.3 0.0013164 0 0.00131632 0 0.00131642 3.3 0.0013163399999999998 3.3 0.0013164399999999999 0 0.00131636 0 0.00131646 3.3 0.00131638 3.3 0.00131648 0 0.0013164 0 0.0013165 3.3 0.00131642 3.3 0.00131652 0 0.0013164399999999999 0 0.00131654 3.3 0.00131646 3.3 0.00131656 0 0.0013164799999999999 0 0.00131658 3.3 0.0013165 3.3 0.0013166 0 0.0013165199999999998 0 0.00131662 3.3 0.00131654 3.3 0.00131664 0 0.0013165599999999998 0 0.0013166599999999999 3.3 0.00131658 3.3 0.00131668 0 0.0013166 0 0.0013167 3.3 0.00131662 3.3 0.00131672 0 0.00131664 0 0.00131674 3.3 0.0013166599999999999 3.3 0.00131676 0 0.00131668 0 0.00131678 3.3 0.0013166999999999999 3.3 0.0013168 0 0.00131672 0 0.00131682 3.3 0.0013167399999999998 3.3 0.00131684 0 0.00131676 0 0.00131686 3.3 0.0013167799999999998 3.3 0.0013168799999999999 0 0.0013168 0 0.0013169 3.3 0.00131682 3.3 0.00131692 0 0.00131684 0 0.00131694 3.3 0.00131686 3.3 0.00131696 0 0.0013168799999999999 0 0.00131698 3.3 0.0013169 3.3 0.001317 0 0.0013169199999999999 0 0.00131702 3.3 0.00131694 3.3 0.00131704 0 0.0013169599999999998 0 0.0013170599999999999 3.3 0.00131698 3.3 0.00131708 0 0.0013169999999999998 0 0.0013170999999999999 3.3 0.00131702 3.3 0.00131712 0 0.00131704 0 0.00131714 3.3 0.0013170599999999999 3.3 0.00131716 0 0.00131708 0 0.00131718 3.3 0.0013170999999999999 3.3 0.0013172 0 0.00131712 0 0.00131722 3.3 0.0013171399999999998 3.3 0.00131724 0 0.00131716 0 0.00131726 3.3 0.0013171799999999998 3.3 0.0013172799999999999 0 0.0013172 0 0.0013173 3.3 0.00131722 3.3 0.00131732 0 0.00131724 0 0.00131734 3.3 0.00131726 3.3 0.00131736 0 0.0013172799999999999 0 0.00131738 3.3 0.0013173 3.3 0.0013174 0 0.0013173199999999999 0 0.00131742 3.3 0.00131734 3.3 0.00131744 0 0.0013173599999999998 0 0.00131746 3.3 0.00131738 3.3 0.00131748 0 0.0013173999999999998 0 0.0013174999999999999 3.3 0.00131742 3.3 0.00131752 0 0.00131744 0 0.00131754 3.3 0.00131746 3.3 0.00131756 0 0.00131748 0 0.00131758 3.3 0.0013174999999999999 3.3 0.0013176 0 0.00131752 0 0.00131762 3.3 0.0013175399999999999 3.3 0.00131764 0 0.00131756 0 0.00131766 3.3 0.0013175799999999998 3.3 0.00131768 0 0.0013176 0 0.0013177 3.3 0.0013176199999999998 3.3 0.0013177199999999999 0 0.00131764 0 0.00131774 3.3 0.00131766 3.3 0.00131776 0 0.00131768 0 0.00131778 3.3 0.0013177 3.3 0.0013178 0 0.0013177199999999999 0 0.00131782 3.3 0.00131774 3.3 0.00131784 0 0.0013177599999999999 0 0.00131786 3.3 0.00131778 3.3 0.00131788 0 0.0013177999999999998 0 0.0013178999999999999 3.3 0.00131782 3.3 0.00131792 0 0.0013178399999999998 0 0.0013179399999999999 3.3 0.00131786 3.3 0.00131796 0 0.00131788 0 0.00131798 3.3 0.0013178999999999999 3.3 0.001318 0 0.00131792 0 0.00131802 3.3 0.0013179399999999999 3.3 0.00131804 0 0.00131796 0 0.00131806 3.3 0.0013179799999999998 3.3 0.00131808 0 0.001318 0 0.0013181 3.3 0.0013180199999999998 3.3 0.0013181199999999999 0 0.00131804 0 0.00131814 3.3 0.00131806 3.3 0.00131816 0 0.00131808 0 0.00131818 3.3 0.0013181 3.3 0.0013182 0 0.0013181199999999999 0 0.00131822 3.3 0.00131814 3.3 0.00131824 0 0.0013181599999999999 0 0.00131826 3.3 0.00131818 3.3 0.00131828 0 0.0013181999999999998 0 0.0013183 3.3 0.00131822 3.3 0.00131832 0 0.0013182399999999998 0 0.0013183399999999999 3.3 0.00131826 3.3 0.00131836 0 0.00131828 0 0.00131838 3.3 0.0013183 3.3 0.0013184 0 0.00131832 0 0.00131842 3.3 0.0013183399999999999 3.3 0.00131844 0 0.00131836 0 0.00131846 3.3 0.0013183799999999999 3.3 0.00131848 0 0.0013184 0 0.0013185 3.3 0.0013184199999999998 3.3 0.00131852 0 0.00131844 0 0.00131854 3.3 0.0013184599999999998 3.3 0.0013185599999999999 0 0.00131848 0 0.00131858 3.3 0.0013185 3.3 0.0013186 0 0.00131852 0 0.00131862 3.3 0.00131854 3.3 0.00131864 0 0.0013185599999999999 0 0.00131866 3.3 0.00131858 3.3 0.00131868 0 0.0013185999999999999 0 0.0013187 3.3 0.00131862 3.3 0.00131872 0 0.0013186399999999998 0 0.0013187399999999999 3.3 0.00131866 3.3 0.00131876 0 0.0013186799999999998 0 0.0013187799999999999 3.3 0.0013187 3.3 0.0013188 0 0.00131872 0 0.00131882 3.3 0.0013187399999999999 3.3 0.00131884 0 0.00131876 0 0.00131886 3.3 0.0013187799999999999 3.3 0.00131888 0 0.0013188 0 0.0013189 3.3 0.0013188199999999998 3.3 0.00131892 0 0.00131884 0 0.00131894 3.3 0.0013188599999999998 3.3 0.0013189599999999999 0 0.00131888 0 0.00131898 3.3 0.0013189 3.3 0.001319 0 0.00131892 0 0.00131902 3.3 0.00131894 3.3 0.00131904 0 0.0013189599999999999 0 0.00131906 3.3 0.00131898 3.3 0.00131908 0 0.0013189999999999999 0 0.0013191 3.3 0.00131902 3.3 0.00131912 0 0.0013190399999999998 0 0.00131914 3.3 0.00131906 3.3 0.00131916 0 0.0013190799999999998 0 0.0013191799999999999 3.3 0.0013191 3.3 0.0013192 0 0.00131912 0 0.00131922 3.3 0.00131914 3.3 0.00131924 0 0.00131916 0 0.00131926 3.3 0.0013191799999999999 3.3 0.00131928 0 0.0013192 0 0.0013193 3.3 0.0013192199999999999 3.3 0.00131932 0 0.00131924 0 0.00131934 3.3 0.0013192599999999998 3.3 0.0013193599999999999 0 0.00131928 0 0.00131938 3.3 0.0013192999999999998 3.3 0.0013193999999999999 0 0.00131932 0 0.00131942 3.3 0.00131934 3.3 0.00131944 0 0.0013193599999999999 0 0.00131946 3.3 0.00131938 3.3 0.00131948 0 0.0013193999999999999 0 0.0013195 3.3 0.00131942 3.3 0.00131952 0 0.0013194399999999998 0 0.00131954 3.3 0.00131946 3.3 0.00131956 0 0.0013194799999999998 0 0.0013195799999999999 3.3 0.0013195 3.3 0.0013196 0 0.00131952 0 0.00131962 3.3 0.00131954 3.3 0.00131964 0 0.00131956 0 0.00131966 3.3 0.0013195799999999999 3.3 0.00131968 0 0.0013196 0 0.0013197 3.3 0.0013196199999999999 3.3 0.00131972 0 0.00131964 0 0.00131974 3.3 0.0013196599999999998 3.3 0.00131976 0 0.00131968 0 0.00131978 3.3 0.0013196999999999998 3.3 0.0013197999999999999 0 0.00131972 0 0.00131982 3.3 0.00131974 3.3 0.00131984 0 0.00131976 0 0.00131986 3.3 0.00131978 3.3 0.00131988 0 0.0013197999999999999 0 0.0013199 3.3 0.00131982 3.3 0.00131992 0 0.0013198399999999999 0 0.00131994 3.3 0.00131986 3.3 0.00131996 0 0.0013198799999999998 0 0.00131998 3.3 0.0013199 3.3 0.00132 0 0.0013199199999999998 0 0.0013200199999999999 3.3 0.00131994 3.3 0.00132004 0 0.00131996 0 0.00132006 3.3 0.00131998 3.3 0.00132008 0 0.00132 0 0.0013201 3.3 0.0013200199999999999 3.3 0.00132012 0 0.00132004 0 0.00132014 3.3 0.0013200599999999999 3.3 0.00132016 0 0.00132008 0 0.00132018 3.3 0.0013200999999999998 3.3 0.0013201999999999999 0 0.00132012 0 0.00132022 3.3 0.0013201399999999998 3.3 0.0013202399999999999 0 0.00132016 0 0.00132026 3.3 0.00132018 3.3 0.00132028 0 0.0013201999999999999 0 0.0013203 3.3 0.00132022 3.3 0.00132032 0 0.0013202399999999999 0 0.00132034 3.3 0.00132026 3.3 0.00132036 0 0.0013202799999999998 0 0.00132038 3.3 0.0013203 3.3 0.0013204 0 0.0013203199999999998 0 0.0013204199999999999 3.3 0.00132034 3.3 0.00132044 0 0.00132036 0 0.00132046 3.3 0.00132038 3.3 0.00132048 0 0.0013204 0 0.0013205 3.3 0.0013204199999999999 3.3 0.00132052 0 0.00132044 0 0.00132054 3.3 0.0013204599999999999 3.3 0.00132056 0 0.00132048 0 0.00132058 3.3 0.0013204999999999998 3.3 0.0013206 0 0.00132052 0 0.00132062 3.3 0.0013205399999999998 3.3 0.0013206399999999999 0 0.00132056 0 0.00132066 3.3 0.00132058 3.3 0.00132068 0 0.0013206 0 0.0013207 3.3 0.00132062 3.3 0.00132072 0 0.0013206399999999999 0 0.00132074 3.3 0.00132066 3.3 0.00132076 0 0.0013206799999999999 0 0.00132078 3.3 0.0013207 3.3 0.0013208 0 0.0013207199999999998 0 0.00132082 3.3 0.00132074 3.3 0.00132084 0 0.0013207599999999998 0 0.0013208599999999999 3.3 0.00132078 3.3 0.00132088 0 0.0013208 0 0.0013209 3.3 0.00132082 3.3 0.00132092 0 0.00132084 0 0.00132094 3.3 0.0013208599999999999 3.3 0.00132096 0 0.00132088 0 0.00132098 3.3 0.0013208999999999999 3.3 0.001321 0 0.00132092 0 0.00132102 3.3 0.0013209399999999998 3.3 0.0013210399999999999 0 0.00132096 0 0.00132106 3.3 0.0013209799999999998 3.3 0.0013210799999999999 0 0.001321 0 0.0013211 3.3 0.00132102 3.3 0.00132112 0 0.0013210399999999999 0 0.00132114 3.3 0.00132106 3.3 0.00132116 0 0.0013210799999999999 0 0.00132118 3.3 0.0013211 3.3 0.0013212 0 0.0013211199999999998 0 0.00132122 3.3 0.00132114 3.3 0.00132124 0 0.0013211599999999998 0 0.0013212599999999999 3.3 0.00132118 3.3 0.00132128 0 0.0013212 0 0.0013213 3.3 0.00132122 3.3 0.00132132 0 0.00132124 0 0.00132134 3.3 0.0013212599999999999 3.3 0.00132136 0 0.00132128 0 0.00132138 3.3 0.0013212999999999999 3.3 0.0013214 0 0.00132132 0 0.00132142 3.3 0.0013213399999999998 3.3 0.00132144 0 0.00132136 0 0.00132146 3.3 0.0013213799999999998 3.3 0.0013214799999999999 0 0.0013214 0 0.0013215 3.3 0.00132142 3.3 0.00132152 0 0.00132144 0 0.00132154 3.3 0.00132146 3.3 0.00132156 0 0.0013214799999999999 0 0.00132158 3.3 0.0013215 3.3 0.0013216 0 0.0013215199999999999 0 0.00132162 3.3 0.00132154 3.3 0.00132164 0 0.0013215599999999998 0 0.00132166 3.3 0.00132158 3.3 0.00132168 0 0.0013215999999999998 0 0.0013216999999999999 3.3 0.00132162 3.3 0.00132172 0 0.00132164 0 0.00132174 3.3 0.00132166 3.3 0.00132176 0 0.00132168 0 0.00132178 3.3 0.0013216999999999999 3.3 0.0013218 0 0.00132172 0 0.00132182 3.3 0.0013217399999999999 3.3 0.00132184 0 0.00132176 0 0.00132186 3.3 0.0013217799999999998 3.3 0.0013218799999999999 0 0.0013218 0 0.0013219 3.3 0.0013218199999999998 3.3 0.0013219199999999999 0 0.00132184 0 0.00132194 3.3 0.00132186 3.3 0.00132196 0 0.0013218799999999999 0 0.00132198 3.3 0.0013219 3.3 0.001322 0 0.0013219199999999999 0 0.00132202 3.3 0.00132194 3.3 0.00132204 0 0.0013219599999999998 0 0.00132206 3.3 0.00132198 3.3 0.00132208 0 0.0013219999999999998 0 0.0013220999999999999 3.3 0.00132202 3.3 0.00132212 0 0.00132204 0 0.00132214 3.3 0.00132206 3.3 0.00132216 0 0.00132208 0 0.00132218 3.3 0.0013220999999999999 3.3 0.0013222 0 0.00132212 0 0.00132222 3.3 0.0013221399999999999 3.3 0.00132224 0 0.00132216 0 0.00132226 3.3 0.0013221799999999998 3.3 0.00132228 0 0.0013222 0 0.0013223 3.3 0.0013222199999999998 3.3 0.0013223199999999999 0 0.00132224 0 0.00132234 3.3 0.00132226 3.3 0.00132236 0 0.00132228 0 0.00132238 3.3 0.0013223 3.3 0.0013224 0 0.0013223199999999999 0 0.00132242 3.3 0.00132234 3.3 0.00132244 0 0.0013223599999999999 0 0.00132246 3.3 0.00132238 3.3 0.00132248 0 0.0013223999999999998 0 0.0013224999999999999 3.3 0.00132242 3.3 0.00132252 0 0.0013224399999999998 0 0.0013225399999999999 3.3 0.00132246 3.3 0.00132256 0 0.00132248 0 0.00132258 3.3 0.0013224999999999999 3.3 0.0013226 0 0.00132252 0 0.00132262 3.3 0.0013225399999999999 3.3 0.00132264 0 0.00132256 0 0.00132266 3.3 0.0013225799999999998 3.3 0.00132268 0 0.0013226 0 0.0013227 3.3 0.0013226199999999998 3.3 0.0013227199999999999 0 0.00132264 0 0.00132274 3.3 0.00132266 3.3 0.00132276 0 0.00132268 0 0.00132278 3.3 0.0013227 3.3 0.0013228 0 0.0013227199999999999 0 0.00132282 3.3 0.00132274 3.3 0.00132284 0 0.0013227599999999999 0 0.00132286 3.3 0.00132278 3.3 0.00132288 0 0.0013227999999999998 0 0.0013229 3.3 0.00132282 3.3 0.00132292 0 0.0013228399999999998 0 0.0013229399999999999 3.3 0.00132286 3.3 0.00132296 0 0.00132288 0 0.00132298 3.3 0.0013229 3.3 0.001323 0 0.00132292 0 0.00132302 3.3 0.0013229399999999999 3.3 0.00132304 0 0.00132296 0 0.00132306 3.3 0.0013229799999999999 3.3 0.00132308 0 0.001323 0 0.0013231 3.3 0.0013230199999999998 3.3 0.00132312 0 0.00132304 0 0.00132314 3.3 0.0013230599999999998 3.3 0.0013231599999999999 0 0.00132308 0 0.00132318 3.3 0.0013231 3.3 0.0013232 0 0.00132312 0 0.00132322 3.3 0.00132314 3.3 0.00132324 0 0.0013231599999999999 0 0.00132326 3.3 0.00132318 3.3 0.00132328 0 0.0013231999999999999 0 0.0013233 3.3 0.00132322 3.3 0.00132332 0 0.0013232399999999998 0 0.0013233399999999999 3.3 0.00132326 3.3 0.00132336 0 0.0013232799999999998 0 0.0013233799999999999 3.3 0.0013233 3.3 0.0013234 0 0.00132332 0 0.00132342 3.3 0.0013233399999999999 3.3 0.00132344 0 0.00132336 0 0.00132346 3.3 0.0013233799999999999 3.3 0.00132348 0 0.0013234 0 0.0013235 3.3 0.0013234199999999998 3.3 0.00132352 0 0.00132344 0 0.00132354 3.3 0.0013234599999999998 3.3 0.0013235599999999999 0 0.00132348 0 0.00132358 3.3 0.0013235 3.3 0.0013236 0 0.00132352 0 0.00132362 3.3 0.00132354 3.3 0.00132364 0 0.0013235599999999999 0 0.00132366 3.3 0.00132358 3.3 0.00132368 0 0.0013235999999999999 0 0.0013237 3.3 0.00132362 3.3 0.00132372 0 0.0013236399999999998 0 0.00132374 3.3 0.00132366 3.3 0.00132376 0 0.0013236799999999998 0 0.0013237799999999999 3.3 0.0013237 3.3 0.0013238 0 0.00132372 0 0.00132382 3.3 0.00132374 3.3 0.00132384 0 0.00132376 0 0.00132386 3.3 0.0013237799999999999 3.3 0.00132388 0 0.0013238 0 0.0013239 3.3 0.0013238199999999999 3.3 0.00132392 0 0.00132384 0 0.00132394 3.3 0.0013238599999999998 3.3 0.00132396 0 0.00132388 0 0.00132398 3.3 0.0013238999999999998 3.3 0.0013239999999999999 0 0.00132392 0 0.00132402 3.3 0.00132394 3.3 0.00132404 0 0.00132396 0 0.00132406 3.3 0.00132398 3.3 0.00132408 0 0.0013239999999999999 0 0.0013241 3.3 0.00132402 3.3 0.00132412 0 0.0013240399999999999 0 0.00132414 3.3 0.00132406 3.3 0.00132416 0 0.0013240799999999998 0 0.0013241799999999999 3.3 0.0013241 3.3 0.0013242 0 0.0013241199999999998 0 0.0013242199999999999 3.3 0.00132414 3.3 0.00132424 0 0.00132416 0 0.00132426 3.3 0.0013241799999999999 3.3 0.00132428 0 0.0013242 0 0.0013243 3.3 0.0013242199999999999 3.3 0.00132432 0 0.00132424 0 0.00132434 3.3 0.0013242599999999998 3.3 0.00132436 0 0.00132428 0 0.00132438 3.3 0.0013242999999999998 3.3 0.0013243999999999999 0 0.00132432 0 0.00132442 3.3 0.00132434 3.3 0.00132444 0 0.00132436 0 0.00132446 3.3 0.00132438 3.3 0.00132448 0 0.0013243999999999999 0 0.0013245 3.3 0.00132442 3.3 0.00132452 0 0.0013244399999999999 0 0.00132454 3.3 0.00132446 3.3 0.00132456 0 0.0013244799999999998 0 0.00132458 3.3 0.0013245 3.3 0.0013246 0 0.0013245199999999998 0 0.0013246199999999999 3.3 0.00132454 3.3 0.00132464 0 0.00132456 0 0.00132466 3.3 0.00132458 3.3 0.00132468 0 0.0013246 0 0.0013247 3.3 0.0013246199999999999 3.3 0.00132472 0 0.00132464 0 0.00132474 3.3 0.0013246599999999999 3.3 0.00132476 0 0.00132468 0 0.00132478 3.3 0.0013246999999999998 3.3 0.0013248 0 0.00132472 0 0.00132482 3.3 0.0013247399999999998 3.3 0.0013248399999999999 0 0.00132476 0 0.00132486 3.3 0.00132478 3.3 0.00132488 0 0.0013248 0 0.0013249 3.3 0.00132482 3.3 0.00132492 0 0.0013248399999999999 0 0.00132494 3.3 0.00132486 3.3 0.00132496 0 0.0013248799999999999 0 0.00132498 3.3 0.0013249 3.3 0.001325 0 0.0013249199999999998 0 0.0013250199999999999 3.3 0.00132494 3.3 0.00132504 0 0.0013249599999999998 0 0.0013250599999999999 3.3 0.00132498 3.3 0.00132508 0 0.001325 0 0.0013251 3.3 0.0013250199999999999 3.3 0.00132512 0 0.00132504 0 0.00132514 3.3 0.0013250599999999999 3.3 0.00132516 0 0.00132508 0 0.00132518 3.3 0.0013250999999999998 3.3 0.0013252 0 0.00132512 0 0.00132522 3.3 0.0013251399999999998 3.3 0.0013252399999999999 0 0.00132516 0 0.00132526 3.3 0.00132518 3.3 0.00132528 0 0.0013252 0 0.0013253 3.3 0.00132522 3.3 0.00132532 0 0.0013252399999999999 0 0.00132534 3.3 0.00132526 3.3 0.00132536 0 0.0013252799999999999 0 0.00132538 3.3 0.0013253 3.3 0.0013254 0 0.0013253199999999998 0 0.00132542 3.3 0.00132534 3.3 0.00132544 0 0.0013253599999999998 0 0.0013254599999999999 3.3 0.00132538 3.3 0.00132548 0 0.0013254 0 0.0013255 3.3 0.00132542 3.3 0.00132552 0 0.00132544 0 0.00132554 3.3 0.0013254599999999999 3.3 0.00132556 0 0.00132548 0 0.00132558 3.3 0.0013254999999999999 3.3 0.0013256 0 0.00132552 0 0.00132562 3.3 0.0013255399999999998 3.3 0.0013256399999999999 0 0.00132556 0 0.00132566 3.3 0.0013255799999999998 3.3 0.0013256799999999999 0 0.0013256 0 0.0013257 3.3 0.00132562 3.3 0.00132572 0 0.0013256399999999999 0 0.00132574 3.3 0.00132566 3.3 0.00132576 0 0.0013256799999999999 0 0.00132578 3.3 0.0013257 3.3 0.0013258 0 0.0013257199999999998 0 0.00132582 3.3 0.00132574 3.3 0.00132584 0 0.0013257599999999998 0 0.0013258599999999999 3.3 0.00132578 3.3 0.00132588 0 0.0013257999999999998 0 0.0013258999999999999 3.3 0.00132582 3.3 0.00132592 0 0.00132584 0 0.00132594 3.3 0.0013258599999999999 3.3 0.00132596 0 0.00132588 0 0.00132598 3.3 0.0013258999999999999 3.3 0.001326 0 0.00132592 0 0.00132602 3.3 0.0013259399999999998 3.3 0.00132604 0 0.00132596 0 0.00132606 3.3 0.0013259799999999998 3.3 0.0013260799999999999 0 0.001326 0 0.0013261 3.3 0.00132602 3.3 0.00132612 0 0.00132604 0 0.00132614 3.3 0.00132606 3.3 0.00132616 0 0.0013260799999999999 0 0.00132618 3.3 0.0013261 3.3 0.0013262 0 0.0013261199999999999 0 0.00132622 3.3 0.00132614 3.3 0.00132624 0 0.0013261599999999998 0 0.00132626 3.3 0.00132618 3.3 0.00132628 0 0.0013261999999999998 0 0.0013262999999999999 3.3 0.00132622 3.3 0.00132632 0 0.00132624 0 0.00132634 3.3 0.00132626 3.3 0.00132636 0 0.00132628 0 0.00132638 3.3 0.0013262999999999999 3.3 0.0013264 0 0.00132632 0 0.00132642 3.3 0.0013263399999999999 3.3 0.00132644 0 0.00132636 0 0.00132646 3.3 0.0013263799999999998 3.3 0.0013264799999999999 0 0.0013264 0 0.0013265 3.3 0.0013264199999999998 3.3 0.0013265199999999999 0 0.00132644 0 0.00132654 3.3 0.00132646 3.3 0.00132656 0 0.0013264799999999999 0 0.00132658 3.3 0.0013265 3.3 0.0013266 0 0.0013265199999999999 0 0.00132662 3.3 0.00132654 3.3 0.00132664 0 0.0013265599999999998 0 0.00132666 3.3 0.00132658 3.3 0.00132668 0 0.0013265999999999998 0 0.0013266999999999999 3.3 0.00132662 3.3 0.00132672 0 0.00132664 0 0.00132674 3.3 0.00132666 3.3 0.00132676 0 0.00132668 0 0.00132678 3.3 0.0013266999999999999 3.3 0.0013268 0 0.00132672 0 0.00132682 3.3 0.0013267399999999999 3.3 0.00132684 0 0.00132676 0 0.00132686 3.3 0.0013267799999999998 3.3 0.00132688 0 0.0013268 0 0.0013269 3.3 0.0013268199999999998 3.3 0.0013269199999999999 0 0.00132684 0 0.00132694 3.3 0.00132686 3.3 0.00132696 0 0.00132688 0 0.00132698 3.3 0.0013269 3.3 0.001327 0 0.0013269199999999999 0 0.00132702 3.3 0.00132694 3.3 0.00132704 0 0.0013269599999999999 0 0.00132706 3.3 0.00132698 3.3 0.00132708 0 0.0013269999999999998 0 0.0013271 3.3 0.00132702 3.3 0.00132712 0 0.0013270399999999998 0 0.0013271399999999999 3.3 0.00132706 3.3 0.00132716 0 0.00132708 0 0.00132718 3.3 0.0013271 3.3 0.0013272 0 0.00132712 0 0.00132722 3.3 0.0013271399999999999 3.3 0.00132724 0 0.00132716 0 0.00132726 3.3 0.0013271799999999999 3.3 0.00132728 0 0.0013272 0 0.0013273 3.3 0.0013272199999999998 3.3 0.0013273199999999999 0 0.00132724 0 0.00132734 3.3 0.0013272599999999998 3.3 0.0013273599999999999 0 0.00132728 0 0.00132738 3.3 0.0013273 3.3 0.0013274 0 0.0013273199999999999 0 0.00132742 3.3 0.00132734 3.3 0.00132744 0 0.0013273599999999999 0 0.00132746 3.3 0.00132738 3.3 0.00132748 0 0.0013273999999999998 0 0.0013275 3.3 0.00132742 3.3 0.00132752 0 0.0013274399999999998 0 0.0013275399999999999 3.3 0.00132746 3.3 0.00132756 0 0.00132748 0 0.00132758 3.3 0.0013275 3.3 0.0013276 0 0.00132752 0 0.00132762 3.3 0.0013275399999999999 3.3 0.00132764 0 0.00132756 0 0.00132766 3.3 0.0013275799999999999 3.3 0.00132768 0 0.0013276 0 0.0013277 3.3 0.0013276199999999998 3.3 0.00132772 0 0.00132764 0 0.00132774 3.3 0.0013276599999999998 3.3 0.0013277599999999999 0 0.00132768 0 0.00132778 3.3 0.0013277 3.3 0.0013278 0 0.00132772 0 0.00132782 3.3 0.00132774 3.3 0.00132784 0 0.0013277599999999999 0 0.00132786 3.3 0.00132778 3.3 0.00132788 0 0.0013277999999999999 0 0.0013279 3.3 0.00132782 3.3 0.00132792 0 0.0013278399999999998 0 0.00132794 3.3 0.00132786 3.3 0.00132796 0 0.0013278799999999998 0 0.0013279799999999999 3.3 0.0013279 3.3 0.001328 0 0.00132792 0 0.00132802 3.3 0.00132794 3.3 0.00132804 0 0.00132796 0 0.00132806 3.3 0.0013279799999999999 3.3 0.00132808 0 0.001328 0 0.0013281 3.3 0.0013280199999999999 3.3 0.00132812 0 0.00132804 0 0.00132814 3.3 0.0013280599999999998 3.3 0.0013281599999999999 0 0.00132808 0 0.00132818 3.3 0.0013280999999999998 3.3 0.0013281999999999999 0 0.00132812 0 0.00132822 3.3 0.00132814 3.3 0.00132824 0 0.0013281599999999999 0 0.00132826 3.3 0.00132818 3.3 0.00132828 0 0.0013281999999999999 0 0.0013283 3.3 0.00132822 3.3 0.00132832 0 0.0013282399999999998 0 0.00132834 3.3 0.00132826 3.3 0.00132836 0 0.0013282799999999998 0 0.0013283799999999999 3.3 0.0013283 3.3 0.0013284 0 0.00132832 0 0.00132842 3.3 0.00132834 3.3 0.00132844 0 0.00132836 0 0.00132846 3.3 0.0013283799999999999 3.3 0.00132848 0 0.0013284 0 0.0013285 3.3 0.0013284199999999999 3.3 0.00132852 0 0.00132844 0 0.00132854 3.3 0.0013284599999999998 3.3 0.00132856 0 0.00132848 0 0.00132858 3.3 0.0013284999999999998 3.3 0.0013285999999999999 0 0.00132852 0 0.00132862 3.3 0.00132854 3.3 0.00132864 0 0.00132856 0 0.00132866 3.3 0.00132858 3.3 0.00132868 0 0.0013285999999999999 0 0.0013287 3.3 0.00132862 3.3 0.00132872 0 0.0013286399999999999 0 0.00132874 3.3 0.00132866 3.3 0.00132876 0 0.0013286799999999998 0 0.00132878 3.3 0.0013287 3.3 0.0013288 0 0.0013287199999999998 0 0.0013288199999999999 3.3 0.00132874 3.3 0.00132884 0 0.00132876 0 0.00132886 3.3 0.00132878 3.3 0.00132888 0 0.0013288 0 0.0013289 3.3 0.0013288199999999999 3.3 0.00132892 0 0.00132884 0 0.00132894 3.3 0.0013288599999999999 3.3 0.00132896 0 0.00132888 0 0.00132898 3.3 0.0013288999999999998 3.3 0.0013289999999999999 0 0.00132892 0 0.00132902 3.3 0.0013289399999999998 3.3 0.0013290399999999999 0 0.00132896 0 0.00132906 3.3 0.00132898 3.3 0.00132908 0 0.0013289999999999999 0 0.0013291 3.3 0.00132902 3.3 0.00132912 0 0.0013290399999999999 0 0.00132914 3.3 0.00132906 3.3 0.00132916 0 0.0013290799999999998 0 0.00132918 3.3 0.0013291 3.3 0.0013292 0 0.0013291199999999998 0 0.0013292199999999999 3.3 0.00132914 3.3 0.00132924 0 0.00132916 0 0.00132926 3.3 0.00132918 3.3 0.00132928 0 0.0013292 0 0.0013293 3.3 0.0013292199999999999 3.3 0.00132932 0 0.00132924 0 0.00132934 3.3 0.0013292599999999999 3.3 0.00132936 0 0.00132928 0 0.00132938 3.3 0.0013292999999999998 3.3 0.0013294 0 0.00132932 0 0.00132942 3.3 0.0013293399999999998 3.3 0.0013294399999999999 0 0.00132936 0 0.00132946 3.3 0.00132938 3.3 0.00132948 0 0.0013294 0 0.0013295 3.3 0.00132942 3.3 0.00132952 0 0.0013294399999999999 0 0.00132954 3.3 0.00132946 3.3 0.00132956 0 0.0013294799999999999 0 0.00132958 3.3 0.0013295 3.3 0.0013296 0 0.0013295199999999998 0 0.0013296199999999999 3.3 0.00132954 3.3 0.00132964 0 0.0013295599999999998 0 0.0013296599999999999 3.3 0.00132958 3.3 0.00132968 0 0.0013296 0 0.0013297 3.3 0.0013296199999999999 3.3 0.00132972 0 0.00132964 0 0.00132974 3.3 0.0013296599999999999 3.3 0.00132976 0 0.00132968 0 0.00132978 3.3 0.0013296999999999998 3.3 0.0013298 0 0.00132972 0 0.00132982 3.3 0.0013297399999999998 3.3 0.0013298399999999999 0 0.00132976 0 0.00132986 3.3 0.00132978 3.3 0.00132988 0 0.0013298 0 0.0013299 3.3 0.00132982 3.3 0.00132992 0 0.0013298399999999999 0 0.00132994 3.3 0.00132986 3.3 0.00132996 0 0.0013298799999999999 0 0.00132998 3.3 0.0013299 3.3 0.00133 0 0.0013299199999999998 0 0.00133002 3.3 0.00132994 3.3 0.00133004 0 0.0013299599999999998 0 0.0013300599999999999 3.3 0.00132998 3.3 0.00133008 0 0.00133 0 0.0013301 3.3 0.00133002 3.3 0.00133012 0 0.00133004 0 0.00133014 3.3 0.0013300599999999999 3.3 0.00133016 0 0.00133008 0 0.00133018 3.3 0.0013300999999999999 3.3 0.0013302 0 0.00133012 0 0.00133022 3.3 0.0013301399999999998 3.3 0.00133024 0 0.00133016 0 0.00133026 3.3 0.0013301799999999998 3.3 0.0013302799999999999 0 0.0013302 0 0.0013303 3.3 0.00133022 3.3 0.00133032 0 0.00133024 0 0.00133034 3.3 0.00133026 3.3 0.00133036 0 0.0013302799999999999 0 0.00133038 3.3 0.0013303 3.3 0.0013304 0 0.0013303199999999999 0 0.00133042 3.3 0.00133034 3.3 0.00133044 0 0.0013303599999999998 0 0.0013304599999999999 3.3 0.00133038 3.3 0.00133048 0 0.0013303999999999998 0 0.0013304999999999999 3.3 0.00133042 3.3 0.00133052 0 0.00133044 0 0.00133054 3.3 0.0013304599999999999 3.3 0.00133056 0 0.00133048 0 0.00133058 3.3 0.0013304999999999999 3.3 0.0013306 0 0.00133052 0 0.00133062 3.3 0.0013305399999999998 3.3 0.00133064 0 0.00133056 0 0.00133066 3.3 0.0013305799999999998 3.3 0.0013306799999999999 0 0.0013306 0 0.0013307 3.3 0.00133062 3.3 0.00133072 0 0.00133064 0 0.00133074 3.3 0.00133066 3.3 0.00133076 0 0.0013306799999999999 0 0.00133078 3.3 0.0013307 3.3 0.0013308 0 0.0013307199999999999 0 0.00133082 3.3 0.00133074 3.3 0.00133084 0 0.0013307599999999998 0 0.00133086 3.3 0.00133078 3.3 0.00133088 0 0.0013307999999999998 0 0.0013308999999999999 3.3 0.00133082 3.3 0.00133092 0 0.00133084 0 0.00133094 3.3 0.00133086 3.3 0.00133096 0 0.00133088 0 0.00133098 3.3 0.0013308999999999999 3.3 0.001331 0 0.00133092 0 0.00133102 3.3 0.0013309399999999999 3.3 0.00133104 0 0.00133096 0 0.00133106 3.3 0.0013309799999999998 3.3 0.00133108 0 0.001331 0 0.0013311 3.3 0.0013310199999999998 3.3 0.0013311199999999999 0 0.00133104 0 0.00133114 3.3 0.00133106 3.3 0.00133116 0 0.00133108 0 0.00133118 3.3 0.0013311 3.3 0.0013312 0 0.0013311199999999999 0 0.00133122 3.3 0.00133114 3.3 0.00133124 0 0.0013311599999999999 0 0.00133126 3.3 0.00133118 3.3 0.00133128 0 0.0013311999999999998 0 0.0013312999999999999 3.3 0.00133122 3.3 0.00133132 0 0.0013312399999999998 0 0.0013313399999999999 3.3 0.00133126 3.3 0.00133136 0 0.00133128 0 0.00133138 3.3 0.0013312999999999999 3.3 0.0013314 0 0.00133132 0 0.00133142 3.3 0.0013313399999999999 3.3 0.00133144 0 0.00133136 0 0.00133146 3.3 0.0013313799999999998 3.3 0.00133148 0 0.0013314 0 0.0013315 3.3 0.0013314199999999998 3.3 0.0013315199999999999 0 0.00133144 0 0.00133154 3.3 0.00133146 3.3 0.00133156 0 0.00133148 0 0.00133158 3.3 0.0013315 3.3 0.0013316 0 0.0013315199999999999 0 0.00133162 3.3 0.00133154 3.3 0.00133164 0 0.0013315599999999999 0 0.00133166 3.3 0.00133158 3.3 0.00133168 0 0.0013315999999999998 0 0.0013317 3.3 0.00133162 3.3 0.00133172 0 0.0013316399999999998 0 0.0013317399999999999 3.3 0.00133166 3.3 0.00133176 0 0.00133168 0 0.00133178 3.3 0.0013317 3.3 0.0013318 0 0.00133172 0 0.00133182 3.3 0.0013317399999999999 3.3 0.00133184 0 0.00133176 0 0.00133186 3.3 0.0013317799999999999 3.3 0.00133188 0 0.0013318 0 0.0013319 3.3 0.0013318199999999998 3.3 0.00133192 0 0.00133184 0 0.00133194 3.3 0.0013318599999999998 3.3 0.0013319599999999999 0 0.00133188 0 0.00133198 3.3 0.0013319 3.3 0.001332 0 0.00133192 0 0.00133202 3.3 0.00133194 3.3 0.00133204 0 0.0013319599999999999 0 0.00133206 3.3 0.00133198 3.3 0.00133208 0 0.0013319999999999999 0 0.0013321 3.3 0.00133202 3.3 0.00133212 0 0.0013320399999999998 0 0.0013321399999999999 3.3 0.00133206 3.3 0.00133216 0 0.0013320799999999998 0 0.0013321799999999999 3.3 0.0013321 3.3 0.0013322 0 0.00133212 0 0.00133222 3.3 0.0013321399999999999 3.3 0.00133224 0 0.00133216 0 0.00133226 3.3 0.0013321799999999999 3.3 0.00133228 0 0.0013322 0 0.0013323 3.3 0.0013322199999999998 3.3 0.00133232 0 0.00133224 0 0.00133234 3.3 0.0013322599999999998 3.3 0.0013323599999999999 0 0.00133228 0 0.00133238 3.3 0.0013323 3.3 0.0013324 0 0.00133232 0 0.00133242 3.3 0.00133234 3.3 0.00133244 0 0.0013323599999999999 0 0.00133246 3.3 0.00133238 3.3 0.00133248 0 0.0013323999999999999 0 0.0013325 3.3 0.00133242 3.3 0.00133252 0 0.0013324399999999998 0 0.00133254 3.3 0.00133246 3.3 0.00133256 0 0.0013324799999999998 0 0.0013325799999999999 3.3 0.0013325 3.3 0.0013326 0 0.00133252 0 0.00133262 3.3 0.00133254 3.3 0.00133264 0 0.00133256 0 0.00133266 3.3 0.0013325799999999999 3.3 0.00133268 0 0.0013326 0 0.0013327 3.3 0.0013326199999999999 3.3 0.00133272 0 0.00133264 0 0.00133274 3.3 0.0013326599999999998 3.3 0.0013327599999999999 0 0.00133268 0 0.00133278 3.3 0.0013326999999999998 3.3 0.0013327999999999999 0 0.00133272 0 0.00133282 3.3 0.00133274 3.3 0.00133284 0 0.0013327599999999999 0 0.00133286 3.3 0.00133278 3.3 0.00133288 0 0.0013327999999999999 0 0.0013329 3.3 0.00133282 3.3 0.00133292 0 0.0013328399999999998 0 0.00133294 3.3 0.00133286 3.3 0.00133296 0 0.0013328799999999998 0 0.0013329799999999999 3.3 0.0013329 3.3 0.001333 0 0.00133292 0 0.00133302 3.3 0.00133294 3.3 0.00133304 0 0.00133296 0 0.00133306 3.3 0.0013329799999999999 3.3 0.00133308 0 0.001333 0 0.0013331 3.3 0.0013330199999999999 3.3 0.00133312 0 0.00133304 0 0.00133314 3.3 0.0013330599999999998 3.3 0.00133316 0 0.00133308 0 0.00133318 3.3 0.0013330999999999998 3.3 0.0013331999999999999 0 0.00133312 0 0.00133322 3.3 0.00133314 3.3 0.00133324 0 0.00133316 0 0.00133326 3.3 0.00133318 3.3 0.00133328 0 0.0013331999999999999 0 0.0013333 3.3 0.00133322 3.3 0.00133332 0 0.0013332399999999999 0 0.00133334 3.3 0.00133326 3.3 0.00133336 0 0.0013332799999999998 0 0.00133338 3.3 0.0013333 3.3 0.0013334 0 0.0013333199999999998 0 0.0013334199999999999 3.3 0.00133334 3.3 0.00133344 0 0.00133336 0 0.00133346 3.3 0.00133338 3.3 0.00133348 0 0.0013334 0 0.0013335 3.3 0.0013334199999999999 3.3 0.00133352 0 0.00133344 0 0.00133354 3.3 0.0013334599999999999 3.3 0.00133356 0 0.00133348 0 0.00133358 3.3 0.0013334999999999998 3.3 0.0013335999999999999 0 0.00133352 0 0.00133362 3.3 0.0013335399999999998 3.3 0.0013336399999999999 0 0.00133356 0 0.00133366 3.3 0.00133358 3.3 0.00133368 0 0.0013335999999999999 0 0.0013337 3.3 0.00133362 3.3 0.00133372 0 0.0013336399999999999 0 0.00133374 3.3 0.00133366 3.3 0.00133376 0 0.0013336799999999998 0 0.00133378 3.3 0.0013337 3.3 0.0013338 0 0.0013337199999999998 0 0.0013338199999999999 3.3 0.00133374 3.3 0.00133384 0 0.00133376 0 0.00133386 3.3 0.00133378 3.3 0.00133388 0 0.0013338 0 0.0013339 3.3 0.0013338199999999999 3.3 0.00133392 0 0.00133384 0 0.00133394 3.3 0.0013338599999999999 3.3 0.00133396 0 0.00133388 0 0.00133398 3.3 0.0013338999999999998 3.3 0.001334 0 0.00133392 0 0.00133402 3.3 0.0013339399999999998 3.3 0.0013340399999999999 0 0.00133396 0 0.00133406 3.3 0.00133398 3.3 0.00133408 0 0.001334 0 0.0013341 3.3 0.00133402 3.3 0.00133412 0 0.0013340399999999999 0 0.00133414 3.3 0.00133406 3.3 0.00133416 0 0.0013340799999999999 0 0.00133418 3.3 0.0013341 3.3 0.0013342 0 0.0013341199999999998 0 0.00133422 3.3 0.00133414 3.3 0.00133424 0 0.0013341599999999998 0 0.0013342599999999999 3.3 0.00133418 3.3 0.00133428 0 0.0013342 0 0.0013343 3.3 0.00133422 3.3 0.00133432 0 0.00133424 0 0.00133434 3.3 0.0013342599999999999 3.3 0.00133436 0 0.00133428 0 0.00133438 3.3 0.0013342999999999999 3.3 0.0013344 0 0.00133432 0 0.00133442 3.3 0.0013343399999999998 3.3 0.0013344399999999999 0 0.00133436 0 0.00133446 3.3 0.0013343799999999998 3.3 0.0013344799999999999 0 0.0013344 0 0.0013345 3.3 0.00133442 3.3 0.00133452 0 0.0013344399999999999 0 0.00133454 3.3 0.00133446 3.3 0.00133456 0 0.0013344799999999999 0 0.00133458 3.3 0.0013345 3.3 0.0013346 0 0.0013345199999999998 0 0.00133462 3.3 0.00133454 3.3 0.00133464 0 0.0013345599999999998 0 0.0013346599999999999 3.3 0.00133458 3.3 0.00133468 0 0.0013346 0 0.0013347 3.3 0.00133462 3.3 0.00133472 0 0.00133464 0 0.00133474 3.3 0.0013346599999999999 3.3 0.00133476 0 0.00133468 0 0.00133478 3.3 0.0013346999999999999 3.3 0.0013348 0 0.00133472 0 0.00133482 3.3 0.0013347399999999998 3.3 0.00133484 0 0.00133476 0 0.00133486 3.3 0.0013347799999999998 3.3 0.0013348799999999999 0 0.0013348 0 0.0013349 3.3 0.00133482 3.3 0.00133492 0 0.00133484 0 0.00133494 3.3 0.00133486 3.3 0.00133496 0 0.0013348799999999999 0 0.00133498 3.3 0.0013349 3.3 0.001335 0 0.0013349199999999999 0 0.00133502 3.3 0.00133494 3.3 0.00133504 0 0.0013349599999999998 0 0.00133506 3.3 0.00133498 3.3 0.00133508 0 0.0013349999999999998 0 0.0013350999999999999 3.3 0.00133502 3.3 0.00133512 0 0.00133504 0 0.00133514 3.3 0.00133506 3.3 0.00133516 0 0.00133508 0 0.00133518 3.3 0.0013350999999999999 3.3 0.0013352 0 0.00133512 0 0.00133522 3.3 0.0013351399999999999 3.3 0.00133524 0 0.00133516 0 0.00133526 3.3 0.0013351799999999998 3.3 0.0013352799999999999 0 0.0013352 0 0.0013353 3.3 0.0013352199999999998 3.3 0.0013353199999999999 0 0.00133524 0 0.00133534 3.3 0.00133526 3.3 0.00133536 0 0.0013352799999999999 0 0.00133538 3.3 0.0013353 3.3 0.0013354 0 0.0013353199999999999 0 0.00133542 3.3 0.00133534 3.3 0.00133544 0 0.0013353599999999998 0 0.00133546 3.3 0.00133538 3.3 0.00133548 0 0.0013353999999999998 0 0.0013354999999999999 3.3 0.00133542 3.3 0.00133552 0 0.00133544 0 0.00133554 3.3 0.00133546 3.3 0.00133556 0 0.00133548 0 0.00133558 3.3 0.0013354999999999999 3.3 0.0013356 0 0.00133552 0 0.00133562 3.3 0.0013355399999999999 3.3 0.00133564 0 0.00133556 0 0.00133566 3.3 0.0013355799999999998 3.3 0.00133568 0 0.0013356 0 0.0013357 3.3 0.0013356199999999998 3.3 0.0013357199999999999 0 0.00133564 0 0.00133574 3.3 0.00133566 3.3 0.00133576 0 0.00133568 0 0.00133578 3.3 0.0013357 3.3 0.0013358 0 0.0013357199999999999 0 0.00133582 3.3 0.00133574 3.3 0.00133584 0 0.0013357599999999999 0 0.00133586 3.3 0.00133578 3.3 0.00133588 0 0.0013357999999999998 0 0.0013358999999999999 3.3 0.00133582 3.3 0.00133592 0 0.0013358399999999998 0 0.0013359399999999999 3.3 0.00133586 3.3 0.00133596 0 0.00133588 0 0.00133598 3.3 0.0013358999999999999 3.3 0.001336 0 0.00133592 0 0.00133602 3.3 0.0013359399999999999 3.3 0.00133604 0 0.00133596 0 0.00133606 3.3 0.0013359799999999998 3.3 0.00133608 0 0.001336 0 0.0013361 3.3 0.0013360199999999998 3.3 0.0013361199999999999 0 0.00133604 0 0.00133614 3.3 0.0013360599999999998 3.3 0.0013361599999999999 0 0.00133608 0 0.00133618 3.3 0.0013361 3.3 0.0013362 0 0.0013361199999999999 0 0.00133622 3.3 0.00133614 3.3 0.00133624 0 0.0013361599999999999 0 0.00133626 3.3 0.00133618 3.3 0.00133628 0 0.0013361999999999998 0 0.0013363 3.3 0.00133622 3.3 0.00133632 0 0.0013362399999999998 0 0.0013363399999999999 3.3 0.00133626 3.3 0.00133636 0 0.00133628 0 0.00133638 3.3 0.0013363 3.3 0.0013364 0 0.00133632 0 0.00133642 3.3 0.0013363399999999999 3.3 0.00133644 0 0.00133636 0 0.00133646 3.3 0.0013363799999999999 3.3 0.00133648 0 0.0013364 0 0.0013365 3.3 0.0013364199999999998 3.3 0.00133652 0 0.00133644 0 0.00133654 3.3 0.0013364599999999998 3.3 0.0013365599999999999 0 0.00133648 0 0.00133658 3.3 0.0013365 3.3 0.0013366 0 0.00133652 0 0.00133662 3.3 0.00133654 3.3 0.00133664 0 0.0013365599999999999 0 0.00133666 3.3 0.00133658 3.3 0.00133668 0 0.0013365999999999999 0 0.0013367 3.3 0.00133662 3.3 0.00133672 0 0.0013366399999999998 0 0.0013367399999999999 3.3 0.00133666 3.3 0.00133676 0 0.0013366799999999998 0 0.0013367799999999999 3.3 0.0013367 3.3 0.0013368 0 0.00133672 0 0.00133682 3.3 0.0013367399999999999 3.3 0.00133684 0 0.00133676 0 0.00133686 3.3 0.0013367799999999999 3.3 0.00133688 0 0.0013368 0 0.0013369 3.3 0.0013368199999999998 3.3 0.00133692 0 0.00133684 0 0.00133694 3.3 0.0013368599999999998 3.3 0.0013369599999999999 0 0.00133688 0 0.00133698 3.3 0.0013369 3.3 0.001337 0 0.00133692 0 0.00133702 3.3 0.00133694 3.3 0.00133704 0 0.0013369599999999999 0 0.00133706 3.3 0.00133698 3.3 0.00133708 0 0.0013369999999999999 0 0.0013371 3.3 0.00133702 3.3 0.00133712 0 0.0013370399999999998 0 0.00133714 3.3 0.00133706 3.3 0.00133716 0 0.0013370799999999998 0 0.0013371799999999999 3.3 0.0013371 3.3 0.0013372 0 0.00133712 0 0.00133722 3.3 0.00133714 3.3 0.00133724 0 0.00133716 0 0.00133726 3.3 0.0013371799999999999 3.3 0.00133728 0 0.0013372 0 0.0013373 3.3 0.0013372199999999999 3.3 0.00133732 0 0.00133724 0 0.00133734 3.3 0.0013372599999999998 3.3 0.00133736 0 0.00133728 0 0.00133738 3.3 0.0013372999999999998 3.3 0.0013373999999999999 0 0.00133732 0 0.00133742 3.3 0.00133734 3.3 0.00133744 0 0.00133736 0 0.00133746 3.3 0.00133738 3.3 0.00133748 0 0.0013373999999999999 0 0.0013375 3.3 0.00133742 3.3 0.00133752 0 0.0013374399999999999 0 0.00133754 3.3 0.00133746 3.3 0.00133756 0 0.0013374799999999998 0 0.0013375799999999999 3.3 0.0013375 3.3 0.0013376 0 0.0013375199999999998 0 0.0013376199999999999 3.3 0.00133754 3.3 0.00133764 0 0.00133756 0 0.00133766 3.3 0.0013375799999999999 3.3 0.00133768 0 0.0013376 0 0.0013377 3.3 0.0013376199999999999 3.3 0.00133772 0 0.00133764 0 0.00133774 3.3 0.0013376599999999998 3.3 0.00133776 0 0.00133768 0 0.00133778 3.3 0.0013376999999999998 3.3 0.0013377999999999999 0 0.00133772 0 0.00133782 3.3 0.00133774 3.3 0.00133784 0 0.00133776 0 0.00133786 3.3 0.00133778 3.3 0.00133788 0 0.0013377999999999999 0 0.0013379 3.3 0.00133782 3.3 0.00133792 0 0.0013378399999999999 0 0.00133794 3.3 0.00133786 3.3 0.00133796 0 0.0013378799999999998 0 0.00133798 3.3 0.0013379 3.3 0.001338 0 0.0013379199999999998 0 0.0013380199999999999 3.3 0.00133794 3.3 0.00133804 0 0.00133796 0 0.00133806 3.3 0.00133798 3.3 0.00133808 0 0.001338 0 0.0013381 3.3 0.0013380199999999999 3.3 0.00133812 0 0.00133804 0 0.00133814 3.3 0.0013380599999999999 3.3 0.00133816 0 0.00133808 0 0.00133818 3.3 0.0013380999999999998 3.3 0.0013382 0 0.00133812 0 0.00133822 3.3 0.0013381399999999998 3.3 0.0013382399999999999 0 0.00133816 0 0.00133826 3.3 0.00133818 3.3 0.00133828 0 0.0013382 0 0.0013383 3.3 0.00133822 3.3 0.00133832 0 0.0013382399999999999 0 0.00133834 3.3 0.00133826 3.3 0.00133836 0 0.0013382799999999999 0 0.00133838 3.3 0.0013383 3.3 0.0013384 0 0.0013383199999999998 0 0.0013384199999999999 3.3 0.00133834 3.3 0.00133844 0 0.0013383599999999998 0 0.0013384599999999999 3.3 0.00133838 3.3 0.00133848 0 0.0013384 0 0.0013385 3.3 0.0013384199999999999 3.3 0.00133852 0 0.00133844 0 0.00133854 3.3 0.0013384599999999999 3.3 0.00133856 0 0.00133848 0 0.00133858 3.3 0.0013384999999999998 3.3 0.0013386 0 0.00133852 0 0.00133862 3.3 0.0013385399999999998 3.3 0.0013386399999999999 0 0.00133856 0 0.00133866 3.3 0.00133858 3.3 0.00133868 0 0.0013386 0 0.0013387 3.3 0.00133862 3.3 0.00133872 0 0.0013386399999999999 0 0.00133874 3.3 0.00133866 3.3 0.00133876 0 0.0013386799999999999 0 0.00133878 3.3 0.0013387 3.3 0.0013388 0 0.0013387199999999998 0 0.00133882 3.3 0.00133874 3.3 0.00133884 0 0.0013387599999999998 0 0.0013388599999999999 3.3 0.00133878 3.3 0.00133888 0 0.0013388 0 0.0013389 3.3 0.00133882 3.3 0.00133892 0 0.00133884 0 0.00133894 3.3 0.0013388599999999999 3.3 0.00133896 0 0.00133888 0 0.00133898 3.3 0.0013388999999999999 3.3 0.001339 0 0.00133892 0 0.00133902 3.3 0.0013389399999999998 3.3 0.00133904 0 0.00133896 0 0.00133906 3.3 0.0013389799999999998 3.3 0.0013390799999999999 0 0.001339 0 0.0013391 3.3 0.00133902 3.3 0.00133912 0 0.00133904 0 0.00133914 3.3 0.00133906 3.3 0.00133916 0 0.0013390799999999999 0 0.00133918 3.3 0.0013391 3.3 0.0013392 0 0.0013391199999999999 0 0.00133922 3.3 0.00133914 3.3 0.00133924 0 0.0013391599999999998 0 0.0013392599999999999 3.3 0.00133918 3.3 0.00133928 0 0.0013391999999999998 0 0.0013392999999999999 3.3 0.00133922 3.3 0.00133932 0 0.00133924 0 0.00133934 3.3 0.0013392599999999999 3.3 0.00133936 0 0.00133928 0 0.00133938 3.3 0.0013392999999999999 3.3 0.0013394 0 0.00133932 0 0.00133942 3.3 0.0013393399999999998 3.3 0.00133944 0 0.00133936 0 0.00133946 3.3 0.0013393799999999998 3.3 0.0013394799999999999 0 0.0013394 0 0.0013395 3.3 0.00133942 3.3 0.00133952 0 0.00133944 0 0.00133954 3.3 0.00133946 3.3 0.00133956 0 0.0013394799999999999 0 0.00133958 3.3 0.0013395 3.3 0.0013396 0 0.0013395199999999999 0 0.00133962 3.3 0.00133954 3.3 0.00133964 0 0.0013395599999999998 0 0.00133966 3.3 0.00133958 3.3 0.00133968 0 0.0013395999999999998 0 0.0013396999999999999 3.3 0.00133962 3.3 0.00133972 0 0.00133964 0 0.00133974 3.3 0.00133966 3.3 0.00133976 0 0.00133968 0 0.00133978 3.3 0.0013396999999999999 3.3 0.0013398 0 0.00133972 0 0.00133982 3.3 0.0013397399999999999 3.3 0.00133984 0 0.00133976 0 0.00133986 3.3 0.0013397799999999998 3.3 0.0013398799999999999 0 0.0013398 0 0.0013399 3.3 0.0013398199999999998 3.3 0.0013399199999999999 0 0.00133984 0 0.00133994 3.3 0.00133986 3.3 0.00133996 0 0.0013398799999999999 0 0.00133998 3.3 0.0013399 3.3 0.00134 0 0.0013399199999999999 0 0.00134002 3.3 0.00133994 3.3 0.00134004 0 0.0013399599999999998 0 0.00134006 3.3 0.00133998 3.3 0.00134008 0 0.0013399999999999998 0 0.0013400999999999999 3.3 0.00134002 3.3 0.00134012 0 0.00134004 0 0.00134014 3.3 0.00134006 3.3 0.00134016 0 0.00134008 0 0.00134018 3.3 0.0013400999999999999 3.3 0.0013402 0 0.00134012 0 0.00134022 3.3 0.0013401399999999999 3.3 0.00134024 0 0.00134016 0 0.00134026 3.3 0.0013401799999999998 3.3 0.00134028 0 0.0013402 0 0.0013403 3.3 0.0013402199999999998 3.3 0.0013403199999999999 0 0.00134024 0 0.00134034 3.3 0.00134026 3.3 0.00134036 0 0.00134028 0 0.00134038 3.3 0.0013403 3.3 0.0013404 0 0.0013403199999999999 0 0.00134042 3.3 0.00134034 3.3 0.00134044 0 0.0013403599999999999 0 0.00134046 3.3 0.00134038 3.3 0.00134048 0 0.0013403999999999998 0 0.0013405 3.3 0.00134042 3.3 0.00134052 0 0.0013404399999999998 0 0.0013405399999999999 3.3 0.00134046 3.3 0.00134056 0 0.00134048 0 0.00134058 3.3 0.0013405 3.3 0.0013406 0 0.00134052 0 0.00134062 3.3 0.0013405399999999999 3.3 0.00134064 0 0.00134056 0 0.00134066 3.3 0.0013405799999999999 3.3 0.00134068 0 0.0013406 0 0.0013407 3.3 0.0013406199999999998 3.3 0.0013407199999999999 0 0.00134064 0 0.00134074 3.3 0.0013406599999999998 3.3 0.0013407599999999999 0 0.00134068 0 0.00134078 3.3 0.0013407 3.3 0.0013408 0 0.0013407199999999999 0 0.00134082 3.3 0.00134074 3.3 0.00134084 0 0.0013407599999999999 0 0.00134086 3.3 0.00134078 3.3 0.00134088 0 0.0013407999999999998 0 0.0013409 3.3 0.00134082 3.3 0.00134092 0 0.0013408399999999998 0 0.0013409399999999999 3.3 0.00134086 3.3 0.00134096 0 0.00134088 0 0.00134098 3.3 0.0013409 3.3 0.001341 0 0.00134092 0 0.00134102 3.3 0.0013409399999999999 3.3 0.00134104 0 0.00134096 0 0.00134106 3.3 0.0013409799999999999 3.3 0.00134108 0 0.001341 0 0.0013411 3.3 0.0013410199999999998 3.3 0.00134112 0 0.00134104 0 0.00134114 3.3 0.0013410599999999998 3.3 0.0013411599999999999 0 0.00134108 0 0.00134118 3.3 0.0013411 3.3 0.0013412 0 0.00134112 0 0.00134122 3.3 0.00134114 3.3 0.00134124 0 0.0013411599999999999 0 0.00134126 3.3 0.00134118 3.3 0.00134128 0 0.0013411999999999999 0 0.0013413 3.3 0.00134122 3.3 0.00134132 0 0.0013412399999999998 0 0.00134134 3.3 0.00134126 3.3 0.00134136 0 0.0013412799999999998 0 0.0013413799999999999 3.3 0.0013413 3.3 0.0013414 0 0.00134132 0 0.00134142 3.3 0.00134134 3.3 0.00134144 0 0.00134136 0 0.00134146 3.3 0.0013413799999999999 3.3 0.00134148 0 0.0013414 0 0.0013415 3.3 0.0013414199999999999 3.3 0.00134152 0 0.00134144 0 0.00134154 3.3 0.0013414599999999998 3.3 0.0013415599999999999 0 0.00134148 0 0.00134158 3.3 0.0013414999999999998 3.3 0.0013415999999999999 0 0.00134152 0 0.00134162 3.3 0.00134154 3.3 0.00134164 0 0.0013415599999999999 0 0.00134166 3.3 0.00134158 3.3 0.00134168 0 0.0013415999999999999 0 0.0013417 3.3 0.00134162 3.3 0.00134172 0 0.0013416399999999998 0 0.00134174 3.3 0.00134166 3.3 0.00134176 0 0.0013416799999999998 0 0.0013417799999999999 3.3 0.0013417 3.3 0.0013418 0 0.00134172 0 0.00134182 3.3 0.00134174 3.3 0.00134184 0 0.00134176 0 0.00134186 3.3 0.0013417799999999999 3.3 0.00134188 0 0.0013418 0 0.0013419 3.3 0.0013418199999999999 3.3 0.00134192 0 0.00134184 0 0.00134194 3.3 0.0013418599999999998 3.3 0.00134196 0 0.00134188 0 0.00134198 3.3 0.0013418999999999998 3.3 0.0013419999999999999 0 0.00134192 0 0.00134202 3.3 0.00134194 3.3 0.00134204 0 0.00134196 0 0.00134206 3.3 0.00134198 3.3 0.00134208 0 0.0013419999999999999 0 0.0013421 3.3 0.00134202 3.3 0.00134212 0 0.0013420399999999999 0 0.00134214 3.3 0.00134206 3.3 0.00134216 0 0.0013420799999999998 0 0.00134218 3.3 0.0013421 3.3 0.0013422 0 0.0013421199999999998 0 0.0013422199999999999 3.3 0.00134214 3.3 0.00134224 0 0.00134216 0 0.00134226 3.3 0.00134218 3.3 0.00134228 0 0.0013422 0 0.0013423 3.3 0.0013422199999999999 3.3 0.00134232 0 0.00134224 0 0.00134234 3.3 0.0013422599999999999 3.3 0.00134236 0 0.00134228 0 0.00134238 3.3 0.0013422999999999998 3.3 0.0013423999999999999 0 0.00134232 0 0.00134242 3.3 0.0013423399999999998 3.3 0.0013424399999999999 0 0.00134236 0 0.00134246 3.3 0.00134238 3.3 0.00134248 0 0.0013423999999999999 0 0.0013425 3.3 0.00134242 3.3 0.00134252 0 0.0013424399999999999 0 0.00134254 3.3 0.00134246 3.3 0.00134256 0 0.0013424799999999998 0 0.00134258 3.3 0.0013425 3.3 0.0013426 0 0.0013425199999999998 0 0.0013426199999999999 3.3 0.00134254 3.3 0.00134264 0 0.00134256 0 0.00134266 3.3 0.00134258 3.3 0.00134268 0 0.0013426 0 0.0013427 3.3 0.0013426199999999999 3.3 0.00134272 0 0.00134264 0 0.00134274 3.3 0.0013426599999999999 3.3 0.00134276 0 0.00134268 0 0.00134278 3.3 0.0013426999999999998 3.3 0.0013428 0 0.00134272 0 0.00134282 3.3 0.0013427399999999998 3.3 0.0013428399999999999 0 0.00134276 0 0.00134286 3.3 0.00134278 3.3 0.00134288 0 0.0013428 0 0.0013429 3.3 0.00134282 3.3 0.00134292 0 0.0013428399999999999 0 0.00134294 3.3 0.00134286 3.3 0.00134296 0 0.0013428799999999999 0 0.00134298 3.3 0.0013429 3.3 0.001343 0 0.0013429199999999998 0 0.0013430199999999999 3.3 0.00134294 3.3 0.00134304 0 0.0013429599999999998 0 0.0013430599999999999 3.3 0.00134298 3.3 0.00134308 0 0.001343 0 0.0013431 3.3 0.0013430199999999999 3.3 0.00134312 0 0.00134304 0 0.00134314 3.3 0.0013430599999999999 3.3 0.00134316 0 0.00134308 0 0.00134318 3.3 0.0013430999999999998 3.3 0.0013432 0 0.00134312 0 0.00134322 3.3 0.0013431399999999998 3.3 0.0013432399999999999 0 0.00134316 0 0.00134326 3.3 0.0013431799999999998 3.3 0.0013432799999999999 0 0.0013432 0 0.0013433 3.3 0.00134322 3.3 0.00134332 0 0.0013432399999999999 0 0.00134334 3.3 0.00134326 3.3 0.00134336 0 0.0013432799999999999 0 0.00134338 3.3 0.0013433 3.3 0.0013434 0 0.0013433199999999998 0 0.00134342 3.3 0.00134334 3.3 0.00134344 0 0.0013433599999999998 0 0.0013434599999999999 3.3 0.00134338 3.3 0.00134348 0 0.0013434 0 0.0013435 3.3 0.00134342 3.3 0.00134352 0 0.00134344 0 0.00134354 3.3 0.0013434599999999999 3.3 0.00134356 0 0.00134348 0 0.00134358 3.3 0.0013434999999999999 3.3 0.0013436 0 0.00134352 0 0.00134362 3.3 0.0013435399999999998 3.3 0.00134364 0 0.00134356 0 0.00134366 3.3 0.0013435799999999998 3.3 0.0013436799999999999 0 0.0013436 0 0.0013437 3.3 0.00134362 3.3 0.00134372 0 0.00134364 0 0.00134374 3.3 0.00134366 3.3 0.00134376 0 0.0013436799999999999 0 0.00134378 3.3 0.0013437 3.3 0.0013438 0 0.0013437199999999999 0 0.00134382 3.3 0.00134374 3.3 0.00134384 0 0.0013437599999999998 0 0.0013438599999999999 3.3 0.00134378 3.3 0.00134388 0 0.0013437999999999998 0 0.0013438999999999999 3.3 0.00134382 3.3 0.00134392 0 0.00134384 0 0.00134394 3.3 0.0013438599999999999 3.3 0.00134396 0 0.00134388 0 0.00134398 3.3 0.0013438999999999999 3.3 0.001344 0 0.00134392 0 0.00134402 3.3 0.0013439399999999998 3.3 0.00134404 0 0.00134396 0 0.00134406 3.3 0.0013439799999999998 3.3 0.0013440799999999999 0 0.001344 0 0.0013441 3.3 0.00134402 3.3 0.00134412 0 0.00134404 0 0.00134414 3.3 0.00134406 3.3 0.00134416 0 0.0013440799999999999 0 0.00134418 3.3 0.0013441 3.3 0.0013442 0 0.0013441199999999999 0 0.00134422 3.3 0.00134414 3.3 0.00134424 0 0.0013441599999999998 0 0.00134426 3.3 0.00134418 3.3 0.00134428 0 0.0013441999999999998 0 0.0013442999999999999 3.3 0.00134422 3.3 0.00134432 0 0.00134424 0 0.00134434 3.3 0.00134426 3.3 0.00134436 0 0.00134428 0 0.00134438 3.3 0.0013442999999999999 3.3 0.0013444 0 0.00134432 0 0.00134442 3.3 0.0013443399999999999 3.3 0.00134444 0 0.00134436 0 0.00134446 3.3 0.0013443799999999998 3.3 0.00134448 0 0.0013444 0 0.0013445 3.3 0.0013444199999999998 3.3 0.0013445199999999999 0 0.00134444 0 0.00134454 3.3 0.00134446 3.3 0.00134456 0 0.00134448 0 0.00134458 3.3 0.0013445 3.3 0.0013446 0 0.0013445199999999999 0 0.00134462 3.3 0.00134454 3.3 0.00134464 0 0.0013445599999999999 0 0.00134466 3.3 0.00134458 3.3 0.00134468 0 0.0013445999999999998 0 0.0013446999999999999 3.3 0.00134462 3.3 0.00134472 0 0.0013446399999999998 0 0.0013447399999999999 3.3 0.00134466 3.3 0.00134476 0 0.00134468 0 0.00134478 3.3 0.0013446999999999999 3.3 0.0013448 0 0.00134472 0 0.00134482 3.3 0.0013447399999999999 3.3 0.00134484 0 0.00134476 0 0.00134486 3.3 0.0013447799999999998 3.3 0.00134488 0 0.0013448 0 0.0013449 3.3 0.0013448199999999998 3.3 0.0013449199999999999 0 0.00134484 0 0.00134494 3.3 0.00134486 3.3 0.00134496 0 0.00134488 0 0.00134498 3.3 0.0013449 3.3 0.001345 0 0.0013449199999999999 0 0.00134502 3.3 0.00134494 3.3 0.00134504 0 0.0013449599999999999 0 0.00134506 3.3 0.00134498 3.3 0.00134508 0 0.0013449999999999998 0 0.0013451 3.3 0.00134502 3.3 0.00134512 0 0.0013450399999999998 0 0.0013451399999999999 3.3 0.00134506 3.3 0.00134516 0 0.00134508 0 0.00134518 3.3 0.0013451 3.3 0.0013452 0 0.00134512 0 0.00134522 3.3 0.0013451399999999999 3.3 0.00134524 0 0.00134516 0 0.00134526 3.3 0.0013451799999999999 3.3 0.00134528 0 0.0013452 0 0.0013453 3.3 0.0013452199999999998 3.3 0.00134532 0 0.00134524 0 0.00134534 3.3 0.0013452599999999998 3.3 0.0013453599999999999 0 0.00134528 0 0.00134538 3.3 0.0013453 3.3 0.0013454 0 0.00134532 0 0.00134542 3.3 0.00134534 3.3 0.00134544 0 0.0013453599999999999 0 0.00134546 3.3 0.00134538 3.3 0.00134548 0 0.0013453999999999999 0 0.0013455 3.3 0.00134542 3.3 0.00134552 0 0.0013454399999999998 0 0.0013455399999999999 3.3 0.00134546 3.3 0.00134556 0 0.0013454799999999998 0 0.0013455799999999999 3.3 0.0013455 3.3 0.0013456 0 0.00134552 0 0.00134562 3.3 0.0013455399999999999 3.3 0.00134564 0 0.00134556 0 0.00134566 3.3 0.0013455799999999999 3.3 0.00134568 0 0.0013456 0 0.0013457 3.3 0.0013456199999999998 3.3 0.00134572 0 0.00134564 0 0.00134574 3.3 0.0013456599999999998 3.3 0.0013457599999999999 0 0.00134568 0 0.00134578 3.3 0.0013457 3.3 0.0013458 0 0.00134572 0 0.00134582 3.3 0.00134574 3.3 0.00134584 0 0.0013457599999999999 0 0.00134586 3.3 0.00134578 3.3 0.00134588 0 0.0013457999999999999 0 0.0013459 3.3 0.00134582 3.3 0.00134592 0 0.0013458399999999998 0 0.00134594 3.3 0.00134586 3.3 0.00134596 0 0.0013458799999999998 0 0.0013459799999999999 3.3 0.0013459 3.3 0.001346 0 0.00134592 0 0.00134602 3.3 0.00134594 3.3 0.00134604 0 0.00134596 0 0.00134606 3.3 0.0013459799999999999 3.3 0.00134608 0 0.001346 0 0.0013461 3.3 0.0013460199999999999 3.3 0.00134612 0 0.00134604 0 0.00134614 3.3 0.0013460599999999998 3.3 0.0013461599999999999 0 0.00134608 0 0.00134618 3.3 0.0013460999999999998 3.3 0.0013461999999999999 0 0.00134612 0 0.00134622 3.3 0.00134614 3.3 0.00134624 0 0.0013461599999999999 0 0.00134626 3.3 0.00134618 3.3 0.00134628 0 0.0013461999999999999 0 0.0013463 3.3 0.00134622 3.3 0.00134632 0 0.0013462399999999998 0 0.00134634 3.3 0.00134626 3.3 0.00134636 0 0.0013462799999999998 0 0.0013463799999999999 3.3 0.0013463 3.3 0.0013464 0 0.0013463199999999998 0 0.0013464199999999999 3.3 0.00134634 3.3 0.00134644 0 0.00134636 0 0.00134646 3.3 0.0013463799999999999 3.3 0.00134648 0 0.0013464 0 0.0013465 3.3 0.0013464199999999999 3.3 0.00134652 0 0.00134644 0 0.00134654 3.3 0.0013464599999999998 3.3 0.00134656 0 0.00134648 0 0.00134658 3.3 0.0013464999999999998 3.3 0.0013465999999999999 0 0.00134652 0 0.00134662 3.3 0.00134654 3.3 0.00134664 0 0.00134656 0 0.00134666 3.3 0.00134658 3.3 0.00134668 0 0.0013465999999999999 0 0.0013467 3.3 0.00134662 3.3 0.00134672 0 0.0013466399999999999 0 0.00134674 3.3 0.00134666 3.3 0.00134676 0 0.0013466799999999998 0 0.00134678 3.3 0.0013467 3.3 0.0013468 0 0.0013467199999999998 0 0.0013468199999999999 3.3 0.00134674 3.3 0.00134684 0 0.00134676 0 0.00134686 3.3 0.00134678 3.3 0.00134688 0 0.0013468 0 0.0013469 3.3 0.0013468199999999999 3.3 0.00134692 0 0.00134684 0 0.00134694 3.3 0.0013468599999999999 3.3 0.00134696 0 0.00134688 0 0.00134698 3.3 0.0013468999999999998 3.3 0.0013469999999999999 0 0.00134692 0 0.00134702 3.3 0.0013469399999999998 3.3 0.0013470399999999999 0 0.00134696 0 0.00134706 3.3 0.00134698 3.3 0.00134708 0 0.0013469999999999999 0 0.0013471 3.3 0.00134702 3.3 0.00134712 0 0.0013470399999999999 0 0.00134714 3.3 0.00134706 3.3 0.00134716 0 0.0013470799999999998 0 0.00134718 3.3 0.0013471 3.3 0.0013472 0 0.0013471199999999998 0 0.0013472199999999999 3.3 0.00134714 3.3 0.00134724 0 0.00134716 0 0.00134726 3.3 0.00134718 3.3 0.00134728 0 0.0013472 0 0.0013473 3.3 0.0013472199999999999 3.3 0.00134732 0 0.00134724 0 0.00134734 3.3 0.0013472599999999999 3.3 0.00134736 0 0.00134728 0 0.00134738 3.3 0.0013472999999999998 3.3 0.0013474 0 0.00134732 0 0.00134742 3.3 0.0013473399999999998 3.3 0.0013474399999999999 0 0.00134736 0 0.00134746 3.3 0.00134738 3.3 0.00134748 0 0.0013474 0 0.0013475 3.3 0.00134742 3.3 0.00134752 0 0.0013474399999999999 0 0.00134754 3.3 0.00134746 3.3 0.00134756 0 0.0013474799999999999 0 0.00134758 3.3 0.0013475 3.3 0.0013476 0 0.0013475199999999998 0 0.00134762 3.3 0.00134754 3.3 0.00134764 0 0.0013475599999999998 0 0.0013476599999999999 3.3 0.00134758 3.3 0.00134768 0 0.0013476 0 0.0013477 3.3 0.00134762 3.3 0.00134772 0 0.00134764 0 0.00134774 3.3 0.0013476599999999999 3.3 0.00134776 0 0.00134768 0 0.00134778 3.3 0.0013476999999999999 3.3 0.0013478 0 0.00134772 0 0.00134782 3.3 0.0013477399999999998 3.3 0.0013478399999999999 0 0.00134776 0 0.00134786 3.3 0.0013477799999999998 3.3 0.0013478799999999999 0 0.0013478 0 0.0013479 3.3 0.00134782 3.3 0.00134792 0 0.0013478399999999999 0 0.00134794 3.3 0.00134786 3.3 0.00134796 0 0.0013478799999999999 0 0.00134798 3.3 0.0013479 3.3 0.001348 0 0.0013479199999999998 0 0.00134802 3.3 0.00134794 3.3 0.00134804 0 0.0013479599999999998 0 0.0013480599999999999 3.3 0.00134798 3.3 0.00134808 0 0.001348 0 0.0013481 3.3 0.00134802 3.3 0.00134812 0 0.00134804 0 0.00134814 3.3 0.0013480599999999999 3.3 0.00134816 0 0.00134808 0 0.00134818 3.3 0.0013480999999999999 3.3 0.0013482 0 0.00134812 0 0.00134822 3.3 0.0013481399999999998 3.3 0.00134824 0 0.00134816 0 0.00134826 3.3 0.0013481799999999998 3.3 0.0013482799999999999 0 0.0013482 0 0.0013483 3.3 0.00134822 3.3 0.00134832 0 0.00134824 0 0.00134834 3.3 0.00134826 3.3 0.00134836 0 0.0013482799999999999 0 0.00134838 3.3 0.0013483 3.3 0.0013484 0 0.0013483199999999999 0 0.00134842 3.3 0.00134834 3.3 0.00134844 0 0.0013483599999999998 0 0.00134846 3.3 0.00134838 3.3 0.00134848 0 0.0013483999999999998 0 0.0013484999999999999 3.3 0.00134842 3.3 0.00134852 0 0.00134844 0 0.00134854 3.3 0.00134846 3.3 0.00134856 0 0.00134848 0 0.00134858 3.3 0.0013484999999999999 3.3 0.0013486 0 0.00134852 0 0.00134862 3.3 0.0013485399999999999 3.3 0.00134864 0 0.00134856 0 0.00134866 3.3 0.0013485799999999998 3.3 0.0013486799999999999 0 0.0013486 0 0.0013487 3.3 0.0013486199999999998 3.3 0.0013487199999999999 0 0.00134864 0 0.00134874 3.3 0.00134866 3.3 0.00134876 0 0.0013486799999999999 0 0.00134878 3.3 0.0013487 3.3 0.0013488 0 0.0013487199999999999 0 0.00134882 3.3 0.00134874 3.3 0.00134884 0 0.0013487599999999998 0 0.00134886 3.3 0.00134878 3.3 0.00134888 0 0.0013487999999999998 0 0.0013488999999999999 3.3 0.00134882 3.3 0.00134892 0 0.00134884 0 0.00134894 3.3 0.00134886 3.3 0.00134896 0 0.00134888 0 0.00134898 3.3 0.0013488999999999999 3.3 0.001349 0 0.00134892 0 0.00134902 3.3 0.0013489399999999999 3.3 0.00134904 0 0.00134896 0 0.00134906 3.3 0.0013489799999999998 3.3 0.00134908 0 0.001349 0 0.0013491 3.3 0.0013490199999999998 3.3 0.0013491199999999999 0 0.00134904 0 0.00134914 3.3 0.00134906 3.3 0.00134916 0 0.00134908 0 0.00134918 3.3 0.0013491 3.3 0.0013492 0 0.0013491199999999999 0 0.00134922 3.3 0.00134914 3.3 0.00134924 0 0.0013491599999999999 0 0.00134926 3.3 0.00134918 3.3 0.00134928 0 0.0013491999999999998 0 0.0013493 3.3 0.00134922 3.3 0.00134932 0 0.0013492399999999998 0 0.0013493399999999999 3.3 0.00134926 3.3 0.00134936 0 0.00134928 0 0.00134938 3.3 0.0013493 3.3 0.0013494 0 0.00134932 0 0.00134942 3.3 0.0013493399999999999 3.3 0.00134944 0 0.00134936 0 0.00134946 3.3 0.0013493799999999999 3.3 0.00134948 0 0.0013494 0 0.0013495 3.3 0.0013494199999999998 3.3 0.0013495199999999999 0 0.00134944 0 0.00134954 3.3 0.0013494599999999998 3.3 0.0013495599999999999 0 0.00134948 0 0.00134958 3.3 0.0013495 3.3 0.0013496 0 0.0013495199999999999 0 0.00134962 3.3 0.00134954 3.3 0.00134964 0 0.0013495599999999999 0 0.00134966 3.3 0.00134958 3.3 0.00134968 0 0.0013495999999999998 0 0.0013497 3.3 0.00134962 3.3 0.00134972 0 0.0013496399999999998 0 0.0013497399999999999 3.3 0.00134966 3.3 0.00134976 0 0.00134968 0 0.00134978 3.3 0.0013497 3.3 0.0013498 0 0.00134972 0 0.00134982 3.3 0.0013497399999999999 3.3 0.00134984 0 0.00134976 0 0.00134986 3.3 0.0013497799999999999 3.3 0.00134988 0 0.0013498 0 0.0013499 3.3 0.0013498199999999998 3.3 0.00134992 0 0.00134984 0 0.00134994 3.3 0.0013498599999999998 3.3 0.0013499599999999999 0 0.00134988 0 0.00134998 3.3 0.0013499 3.3 0.00135 0 0.00134992 0 0.00135002 3.3 0.00134994 3.3 0.00135004 0 0.0013499599999999999 0 0.00135006 3.3 0.00134998 3.3 0.00135008 0 0.0013499999999999999 0 0.0013501 3.3 0.00135002 3.3 0.00135012 0 0.0013500399999999998 0 0.0013501399999999999 3.3 0.00135006 3.3 0.00135016 0 0.0013500799999999998 0 0.0013501799999999999 3.3 0.0013501 3.3 0.0013502 0 0.00135012 0 0.00135022 3.3 0.0013501399999999999 3.3 0.00135024 0 0.00135016 0 0.00135026 3.3 0.0013501799999999999 3.3 0.00135028 0 0.0013502 0 0.0013503 3.3 0.0013502199999999998 3.3 0.00135032 0 0.00135024 0 0.00135034 3.3 0.0013502599999999998 3.3 0.0013503599999999999 0 0.00135028 0 0.00135038 3.3 0.0013503 3.3 0.0013504 0 0.00135032 0 0.00135042 3.3 0.00135034 3.3 0.00135044 0 0.0013503599999999999 0 0.00135046 3.3 0.00135038 3.3 0.00135048 0 0.0013503999999999999 0 0.0013505 3.3 0.00135042 3.3 0.00135052 0 0.0013504399999999998 0 0.00135054 3.3 0.00135046 3.3 0.00135056 0 0.0013504799999999998 0 0.0013505799999999999 3.3 0.0013505 3.3 0.0013506 0 0.00135052 0 0.00135062 3.3 0.00135054 3.3 0.00135064 0 0.00135056 0 0.00135066 3.3 0.0013505799999999999 3.3 0.00135068 0 0.0013506 0 0.0013507 3.3 0.0013506199999999999 3.3 0.00135072 0 0.00135064 0 0.00135074 3.3 0.0013506599999999998 3.3 0.00135076 0 0.00135068 0 0.00135078 3.3 0.0013506999999999998 3.3 0.0013507999999999999 0 0.00135072 0 0.00135082 3.3 0.00135074 3.3 0.00135084 0 0.00135076 0 0.00135086 3.3 0.00135078 3.3 0.00135088 0 0.0013507999999999999 0 0.0013509 3.3 0.00135082 3.3 0.00135092 0 0.0013508399999999999 0 0.00135094 3.3 0.00135086 3.3 0.00135096 0 0.0013508799999999998 0 0.0013509799999999999 3.3 0.0013509 3.3 0.001351 0 0.0013509199999999998 0 0.0013510199999999999 3.3 0.00135094 3.3 0.00135104 0 0.00135096 0 0.00135106 3.3 0.0013509799999999999 3.3 0.00135108 0 0.001351 0 0.0013511 3.3 0.0013510199999999999 3.3 0.00135112 0 0.00135104 0 0.00135114 3.3 0.0013510599999999998 3.3 0.00135116 0 0.00135108 0 0.00135118 3.3 0.0013510999999999998 3.3 0.0013511999999999999 0 0.00135112 0 0.00135122 3.3 0.00135114 3.3 0.00135124 0 0.00135116 0 0.00135126 3.3 0.00135118 3.3 0.00135128 0 0.0013511999999999999 0 0.0013513 3.3 0.00135122 3.3 0.00135132 0 0.0013512399999999999 0 0.00135134 3.3 0.00135126 3.3 0.00135136 0 0.0013512799999999998 0 0.00135138 3.3 0.0013513 3.3 0.0013514 0 0.0013513199999999998 0 0.0013514199999999999 3.3 0.00135134 3.3 0.00135144 0 0.00135136 0 0.00135146 3.3 0.00135138 3.3 0.00135148 0 0.0013514 0 0.0013515 3.3 0.0013514199999999999 3.3 0.00135152 0 0.00135144 0 0.00135154 3.3 0.0013514599999999999 3.3 0.00135156 0 0.00135148 0 0.00135158 3.3 0.0013514999999999998 3.3 0.0013516 0 0.00135152 0 0.00135162 3.3 0.0013515399999999998 3.3 0.0013516399999999999 0 0.00135156 0 0.00135166 3.3 0.00135158 3.3 0.00135168 0 0.0013516 0 0.0013517 3.3 0.00135162 3.3 0.00135172 0 0.0013516399999999999 0 0.00135174 3.3 0.00135166 3.3 0.00135176 0 0.0013516799999999999 0 0.00135178 3.3 0.0013517 3.3 0.0013518 0 0.0013517199999999998 0 0.0013518199999999999 3.3 0.00135174 3.3 0.00135184 0 0.0013517599999999998 0 0.0013518599999999999 3.3 0.00135178 3.3 0.00135188 0 0.0013518 0 0.0013519 3.3 0.0013518199999999999 3.3 0.00135192 0 0.00135184 0 0.00135194 3.3 0.0013518599999999999 3.3 0.00135196 0 0.00135188 0 0.00135198 3.3 0.0013518999999999998 3.3 0.001352 0 0.00135192 0 0.00135202 3.3 0.0013519399999999998 3.3 0.0013520399999999999 0 0.00135196 0 0.00135206 3.3 0.00135198 3.3 0.00135208 0 0.001352 0 0.0013521 3.3 0.00135202 3.3 0.00135212 0 0.0013520399999999999 0 0.00135214 3.3 0.00135206 3.3 0.00135216 0 0.0013520799999999999 0 0.00135218 3.3 0.0013521 3.3 0.0013522 0 0.0013521199999999998 0 0.00135222 3.3 0.00135214 3.3 0.00135224 0 0.0013521599999999998 0 0.0013522599999999999 3.3 0.00135218 3.3 0.00135228 0 0.0013522 0 0.0013523 3.3 0.00135222 3.3 0.00135232 0 0.00135224 0 0.00135234 3.3 0.0013522599999999999 3.3 0.00135236 0 0.00135228 0 0.00135238 3.3 0.0013522999999999999 3.3 0.0013524 0 0.00135232 0 0.00135242 3.3 0.0013523399999999998 3.3 0.00135244 0 0.00135236 0 0.00135246 3.3 0.0013523799999999998 3.3 0.0013524799999999999 0 0.0013524 0 0.0013525 3.3 0.00135242 3.3 0.00135252 0 0.00135244 0 0.00135254 3.3 0.00135246 3.3 0.00135256 0 0.0013524799999999999 0 0.00135258 3.3 0.0013525 3.3 0.0013526 0 0.0013525199999999999 0 0.00135262 3.3 0.00135254 3.3 0.00135264 0 0.0013525599999999998 0 0.0013526599999999999 3.3 0.00135258 3.3 0.00135268 0 0.0013525999999999998 0 0.0013526999999999999 3.3 0.00135262 3.3 0.00135272 0 0.00135264 0 0.00135274 3.3 0.0013526599999999999 3.3 0.00135276 0 0.00135268 0 0.00135278 3.3 0.0013526999999999999 3.3 0.0013528 0 0.00135272 0 0.00135282 3.3 0.0013527399999999998 3.3 0.00135284 0 0.00135276 0 0.00135286 3.3 0.0013527799999999998 3.3 0.0013528799999999999 0 0.0013528 0 0.0013529 3.3 0.00135282 3.3 0.00135292 0 0.00135284 0 0.00135294 3.3 0.00135286 3.3 0.00135296 0 0.0013528799999999999 0 0.00135298 3.3 0.0013529 3.3 0.001353 0 0.0013529199999999999 0 0.00135302 3.3 0.00135294 3.3 0.00135304 0 0.0013529599999999998 0 0.00135306 3.3 0.00135298 3.3 0.00135308 0 0.0013529999999999998 0 0.0013530999999999999 3.3 0.00135302 3.3 0.00135312 0 0.00135304 0 0.00135314 3.3 0.00135306 3.3 0.00135316 0 0.00135308 0 0.00135318 3.3 0.0013530999999999999 3.3 0.0013532 0 0.00135312 0 0.00135322 3.3 0.0013531399999999999 3.3 0.00135324 0 0.00135316 0 0.00135326 3.3 0.0013531799999999998 3.3 0.0013532799999999999 0 0.0013532 0 0.0013533 3.3 0.0013532199999999998 3.3 0.0013533199999999999 0 0.00135324 0 0.00135334 3.3 0.00135326 3.3 0.00135336 0 0.0013532799999999999 0 0.00135338 3.3 0.0013533 3.3 0.0013534 0 0.0013533199999999999 0 0.00135342 3.3 0.00135334 3.3 0.00135344 0 0.0013533599999999998 0 0.00135346 3.3 0.00135338 3.3 0.00135348 0 0.0013533999999999998 0 0.0013534999999999999 3.3 0.00135342 3.3 0.00135352 0 0.0013534399999999998 0 0.0013535399999999999 3.3 0.00135346 3.3 0.00135356 0 0.00135348 0 0.00135358 3.3 0.0013534999999999999 3.3 0.0013536 0 0.00135352 0 0.00135362 3.3 0.0013535399999999999 3.3 0.00135364 0 0.00135356 0 0.00135366 3.3 0.0013535799999999998 3.3 0.00135368 0 0.0013536 0 0.0013537 3.3 0.0013536199999999998 3.3 0.0013537199999999999 0 0.00135364 0 0.00135374 3.3 0.00135366 3.3 0.00135376 0 0.00135368 0 0.00135378 3.3 0.0013537 3.3 0.0013538 0 0.0013537199999999999 0 0.00135382 3.3 0.00135374 3.3 0.00135384 0 0.0013537599999999999 0 0.00135386 3.3 0.00135378 3.3 0.00135388 0 0.0013537999999999998 0 0.0013539 3.3 0.00135382 3.3 0.00135392 0 0.0013538399999999998 0 0.0013539399999999999 3.3 0.00135386 3.3 0.00135396 0 0.00135388 0 0.00135398 3.3 0.0013539 3.3 0.001354 0 0.00135392 0 0.00135402 3.3 0.0013539399999999999 3.3 0.00135404 0 0.00135396 0 0.00135406 3.3 0.0013539799999999999 3.3 0.00135408 0 0.001354 0 0.0013541 3.3 0.0013540199999999998 3.3 0.0013541199999999999 0 0.00135404 0 0.00135414 3.3 0.0013540599999999998 3.3 0.0013541599999999999 0 0.00135408 0 0.00135418 3.3 0.0013541 3.3 0.0013542 0 0.0013541199999999999 0 0.00135422 3.3 0.00135414 3.3 0.00135424 0 0.0013541599999999999 0 0.00135426 3.3 0.00135418 3.3 0.00135428 0 0.0013541999999999998 0 0.0013543 3.3 0.00135422 3.3 0.00135432 0 0.0013542399999999998 0 0.0013543399999999999 3.3 0.00135426 3.3 0.00135436 0 0.00135428 0 0.00135438 3.3 0.0013543 3.3 0.0013544 0 0.00135432 0 0.00135442 3.3 0.0013543399999999999 3.3 0.00135444 0 0.00135436 0 0.00135446 3.3 0.0013543799999999999 3.3 0.00135448 0 0.0013544 0 0.0013545 3.3 0.0013544199999999998 3.3 0.00135452 0 0.00135444 0 0.00135454 3.3 0.0013544599999999998 3.3 0.0013545599999999999 0 0.00135448 0 0.00135458 3.3 0.0013545 3.3 0.0013546 0 0.00135452 0 0.00135462 3.3 0.00135454 3.3 0.00135464 0 0.0013545599999999999 0 0.00135466 3.3 0.00135458 3.3 0.00135468 0 0.0013545999999999999 0 0.0013547 3.3 0.00135462 3.3 0.00135472 0 0.0013546399999999998 0 0.00135474 3.3 0.00135466 3.3 0.00135476 0 0.0013546799999999998 0 0.0013547799999999999 3.3 0.0013547 3.3 0.0013548 0 0.00135472 0 0.00135482 3.3 0.00135474 3.3 0.00135484 0 0.00135476 0 0.00135486 3.3 0.0013547799999999999 3.3 0.00135488 0 0.0013548 0 0.0013549 3.3 0.0013548199999999999 3.3 0.00135492 0 0.00135484 0 0.00135494 3.3 0.0013548599999999998 3.3 0.0013549599999999999 0 0.00135488 0 0.00135498 3.3 0.0013548999999999998 3.3 0.0013549999999999999 0 0.00135492 0 0.00135502 3.3 0.00135494 3.3 0.00135504 0 0.0013549599999999999 0 0.00135506 3.3 0.00135498 3.3 0.00135508 0 0.0013549999999999999 0 0.0013551 3.3 0.00135502 3.3 0.00135512 0 0.0013550399999999998 0 0.00135514 3.3 0.00135506 3.3 0.00135516 0 0.0013550799999999998 0 0.0013551799999999999 3.3 0.0013551 3.3 0.0013552 0 0.00135512 0 0.00135522 3.3 0.00135514 3.3 0.00135524 0 0.00135516 0 0.00135526 3.3 0.0013551799999999999 3.3 0.00135528 0 0.0013552 0 0.0013553 3.3 0.0013552199999999999 3.3 0.00135532 0 0.00135524 0 0.00135534 3.3 0.0013552599999999998 3.3 0.00135536 0 0.00135528 0 0.00135538 3.3 0.0013552999999999998 3.3 0.0013553999999999999 0 0.00135532 0 0.00135542 3.3 0.00135534 3.3 0.00135544 0 0.00135536 0 0.00135546 3.3 0.00135538 3.3 0.00135548 0 0.0013553999999999999 0 0.0013555 3.3 0.00135542 3.3 0.00135552 0 0.0013554399999999999 0 0.00135554 3.3 0.00135546 3.3 0.00135556 0 0.0013554799999999998 0 0.00135558 3.3 0.0013555 3.3 0.0013556 0 0.0013555199999999998 0 0.0013556199999999999 3.3 0.00135554 3.3 0.00135564 0 0.00135556 0 0.00135566 3.3 0.00135558 3.3 0.00135568 0 0.0013556 0 0.0013557 3.3 0.0013556199999999999 3.3 0.00135572 0 0.00135564 0 0.00135574 3.3 0.0013556599999999999 3.3 0.00135576 0 0.00135568 0 0.00135578 3.3 0.0013556999999999998 3.3 0.0013557999999999999 0 0.00135572 0 0.00135582 3.3 0.0013557399999999998 3.3 0.0013558399999999999 0 0.00135576 0 0.00135586 3.3 0.00135578 3.3 0.00135588 0 0.0013557999999999999 0 0.0013559 3.3 0.00135582 3.3 0.00135592 0 0.0013558399999999999 0 0.00135594 3.3 0.00135586 3.3 0.00135596 0 0.0013558799999999998 0 0.00135598 3.3 0.0013559 3.3 0.001356 0 0.0013559199999999998 0 0.0013560199999999999 3.3 0.00135594 3.3 0.00135604 0 0.00135596 0 0.00135606 3.3 0.00135598 3.3 0.00135608 0 0.001356 0 0.0013561 3.3 0.0013560199999999999 3.3 0.00135612 0 0.00135604 0 0.00135614 3.3 0.0013560599999999999 3.3 0.00135616 0 0.00135608 0 0.00135618 3.3 0.0013560999999999998 3.3 0.0013562 0 0.00135612 0 0.00135622 3.3 0.0013561399999999998 3.3 0.0013562399999999999 0 0.00135616 0 0.00135626 3.3 0.00135618 3.3 0.00135628 0 0.0013562 0 0.0013563 3.3 0.00135622 3.3 0.00135632 0 0.0013562399999999999 0 0.00135634 3.3 0.00135626 3.3 0.00135636 0 0.0013562799999999999 0 0.00135638 3.3 0.0013563 3.3 0.0013564 0 0.0013563199999999998 0 0.0013564199999999999 3.3 0.00135634 3.3 0.00135644 0 0.0013563599999999998 0 0.0013564599999999999 3.3 0.00135638 3.3 0.00135648 0 0.0013564 0 0.0013565 3.3 0.0013564199999999999 3.3 0.00135652 0 0.00135644 0 0.00135654 3.3 0.0013564599999999999 3.3 0.00135656 0 0.00135648 0 0.00135658 3.3 0.0013564999999999998 3.3 0.0013566 0 0.00135652 0 0.00135662 3.3 0.0013565399999999998 3.3 0.0013566399999999999 0 0.00135656 0 0.00135666 3.3 0.0013565799999999998 3.3 0.0013566799999999999 0 0.0013566 0 0.0013567 3.3 0.00135662 3.3 0.00135672 0 0.0013566399999999999 0 0.00135674 3.3 0.00135666 3.3 0.00135676 0 0.0013566799999999999 0 0.00135678 3.3 0.0013567 3.3 0.0013568 0 0.0013567199999999998 0 0.00135682 3.3 0.00135674 3.3 0.00135684 0 0.0013567599999999998 0 0.0013568599999999999 3.3 0.00135678 3.3 0.00135688 0 0.0013568 0 0.0013569 3.3 0.00135682 3.3 0.00135692 0 0.00135684 0 0.00135694 3.3 0.0013568599999999999 3.3 0.00135696 0 0.00135688 0 0.00135698 3.3 0.0013568999999999999 3.3 0.001357 0 0.00135692 0 0.00135702 3.3 0.0013569399999999998 3.3 0.00135704 0 0.00135696 0 0.00135706 3.3 0.0013569799999999998 3.3 0.0013570799999999999 0 0.001357 0 0.0013571 3.3 0.00135702 3.3 0.00135712 0 0.00135704 0 0.00135714 3.3 0.00135706 3.3 0.00135716 0 0.0013570799999999999 0 0.00135718 3.3 0.0013571 3.3 0.0013572 0 0.0013571199999999999 0 0.00135722 3.3 0.00135714 3.3 0.00135724 0 0.0013571599999999998 0 0.0013572599999999999 3.3 0.00135718 3.3 0.00135728 0 0.0013571999999999998 0 0.0013572999999999999 3.3 0.00135722 3.3 0.00135732 0 0.00135724 0 0.00135734 3.3 0.0013572599999999999 3.3 0.00135736 0 0.00135728 0 0.00135738 3.3 0.0013572999999999999 3.3 0.0013574 0 0.00135732 0 0.00135742 3.3 0.0013573399999999998 3.3 0.00135744 0 0.00135736 0 0.00135746 3.3 0.0013573799999999998 3.3 0.0013574799999999999 0 0.0013574 0 0.0013575 3.3 0.00135742 3.3 0.00135752 0 0.00135744 0 0.00135754 3.3 0.00135746 3.3 0.00135756 0 0.0013574799999999999 0 0.00135758 3.3 0.0013575 3.3 0.0013576 0 0.0013575199999999999 0 0.00135762 3.3 0.00135754 3.3 0.00135764 0 0.0013575599999999998 0 0.00135766 3.3 0.00135758 3.3 0.00135768 0 0.0013575999999999998 0 0.0013576999999999999 3.3 0.00135762 3.3 0.00135772 0 0.00135764 0 0.00135774 3.3 0.00135766 3.3 0.00135776 0 0.00135768 0 0.00135778 3.3 0.0013576999999999999 3.3 0.0013578 0 0.00135772 0 0.00135782 3.3 0.0013577399999999999 3.3 0.00135784 0 0.00135776 0 0.00135786 3.3 0.0013577799999999998 3.3 0.00135788 0 0.0013578 0 0.0013579 3.3 0.0013578199999999998 3.3 0.0013579199999999999 0 0.00135784 0 0.00135794 3.3 0.00135786 3.3 0.00135796 0 0.00135788 0 0.00135798 3.3 0.0013579 3.3 0.001358 0 0.0013579199999999999 0 0.00135802 3.3 0.00135794 3.3 0.00135804 0 0.0013579599999999999 0 0.00135806 3.3 0.00135798 3.3 0.00135808 0 0.0013579999999999998 0 0.0013580999999999999 3.3 0.00135802 3.3 0.00135812 0 0.0013580399999999998 0 0.0013581399999999999 3.3 0.00135806 3.3 0.00135816 0 0.00135808 0 0.00135818 3.3 0.0013580999999999999 3.3 0.0013582 0 0.00135812 0 0.00135822 3.3 0.0013581399999999999 3.3 0.00135824 0 0.00135816 0 0.00135826 3.3 0.0013581799999999998 3.3 0.00135828 0 0.0013582 0 0.0013583 3.3 0.0013582199999999998 3.3 0.0013583199999999999 0 0.00135824 0 0.00135834 3.3 0.00135826 3.3 0.00135836 0 0.00135828 0 0.00135838 3.3 0.0013583 3.3 0.0013584 0 0.0013583199999999999 0 0.00135842 3.3 0.00135834 3.3 0.00135844 0 0.0013583599999999999 0 0.00135846 3.3 0.00135838 3.3 0.00135848 0 0.0013583999999999998 0 0.0013585 3.3 0.00135842 3.3 0.00135852 0 0.0013584399999999998 0 0.0013585399999999999 3.3 0.00135846 3.3 0.00135856 0 0.00135848 0 0.00135858 3.3 0.0013585 3.3 0.0013586 0 0.00135852 0 0.00135862 3.3 0.0013585399999999999 3.3 0.00135864 0 0.00135856 0 0.00135866 3.3 0.0013585799999999999 3.3 0.00135868 0 0.0013586 0 0.0013587 3.3 0.0013586199999999998 3.3 0.00135872 0 0.00135864 0 0.00135874 3.3 0.0013586599999999998 3.3 0.0013587599999999999 0 0.00135868 0 0.00135878 3.3 0.0013587 3.3 0.0013588 0 0.00135872 0 0.00135882 3.3 0.00135874 3.3 0.00135884 0 0.0013587599999999999 0 0.00135886 3.3 0.00135878 3.3 0.00135888 0 0.0013587999999999999 0 0.0013589 3.3 0.00135882 3.3 0.00135892 0 0.0013588399999999998 0 0.0013589399999999999 3.3 0.00135886 3.3 0.00135896 0 0.0013588799999999998 0 0.0013589799999999999 3.3 0.0013589 3.3 0.001359 0 0.00135892 0 0.00135902 3.3 0.0013589399999999999 3.3 0.00135904 0 0.00135896 0 0.00135906 3.3 0.0013589799999999999 3.3 0.00135908 0 0.001359 0 0.0013591 3.3 0.0013590199999999998 3.3 0.00135912 0 0.00135904 0 0.00135914 3.3 0.0013590599999999998 3.3 0.0013591599999999999 0 0.00135908 0 0.00135918 3.3 0.0013591 3.3 0.0013592 0 0.00135912 0 0.00135922 3.3 0.00135914 3.3 0.00135924 0 0.0013591599999999999 0 0.00135926 3.3 0.00135918 3.3 0.00135928 0 0.0013591999999999999 0 0.0013593 3.3 0.00135922 3.3 0.00135932 0 0.0013592399999999998 0 0.00135934 3.3 0.00135926 3.3 0.00135936 0 0.0013592799999999998 0 0.0013593799999999999 3.3 0.0013593 3.3 0.0013594 0 0.00135932 0 0.00135942 3.3 0.00135934 3.3 0.00135944 0 0.00135936 0 0.00135946 3.3 0.0013593799999999999 3.3 0.00135948 0 0.0013594 0 0.0013595 3.3 0.0013594199999999999 3.3 0.00135952 0 0.00135944 0 0.00135954 3.3 0.0013594599999999998 3.3 0.00135956 0 0.00135948 0 0.00135958 3.3 0.0013594999999999998 3.3 0.0013595999999999999 0 0.00135952 0 0.00135962 3.3 0.00135954 3.3 0.00135964 0 0.00135956 0 0.00135966 3.3 0.00135958 3.3 0.00135968 0 0.0013595999999999999 0 0.0013597 3.3 0.00135962 3.3 0.00135972 0 0.0013596399999999999 0 0.00135974 3.3 0.00135966 3.3 0.00135976 0 0.0013596799999999998 0 0.0013597799999999999 3.3 0.0013597 3.3 0.0013598 0 0.0013597199999999998 0 0.0013598199999999999 3.3 0.00135974 3.3 0.00135984 0 0.00135976 0 0.00135986 3.3 0.0013597799999999999 3.3 0.00135988 0 0.0013598 0 0.0013599 3.3 0.0013598199999999999 3.3 0.00135992 0 0.00135984 0 0.00135994 3.3 0.0013598599999999998 3.3 0.00135996 0 0.00135988 0 0.00135998 3.3 0.0013598999999999998 3.3 0.0013599999999999999 0 0.00135992 0 0.00136002 3.3 0.00135994 3.3 0.00136004 0 0.00135996 0 0.00136006 3.3 0.00135998 3.3 0.00136008 0 0.0013599999999999999 0 0.0013601 3.3 0.00136002 3.3 0.00136012 0 0.0013600399999999999 0 0.00136014 3.3 0.00136006 3.3 0.00136016 0 0.0013600799999999998 0 0.00136018 3.3 0.0013601 3.3 0.0013602 0 0.0013601199999999998 0 0.0013602199999999999 3.3 0.00136014 3.3 0.00136024 0 0.00136016 0 0.00136026 3.3 0.00136018 3.3 0.00136028 0 0.0013602 0 0.0013603 3.3 0.0013602199999999999 3.3 0.00136032 0 0.00136024 0 0.00136034 3.3 0.0013602599999999999 3.3 0.00136036 0 0.00136028 0 0.00136038 3.3 0.0013602999999999998 3.3 0.0013603999999999999 0 0.00136032 0 0.00136042 3.3 0.0013603399999999998 3.3 0.0013604399999999999 0 0.00136036 0 0.00136046 3.3 0.00136038 3.3 0.00136048 0 0.0013603999999999999 0 0.0013605 3.3 0.00136042 3.3 0.00136052 0 0.0013604399999999999 0 0.00136054 3.3 0.00136046 3.3 0.00136056 0 0.0013604799999999998 0 0.00136058 3.3 0.0013605 3.3 0.0013606 0 0.0013605199999999998 0 0.0013606199999999999 3.3 0.00136054 3.3 0.00136064 0 0.0013605599999999998 0 0.0013606599999999999 3.3 0.00136058 3.3 0.00136068 0 0.0013606 0 0.0013607 3.3 0.0013606199999999999 3.3 0.00136072 0 0.00136064 0 0.00136074 3.3 0.0013606599999999999 3.3 0.00136076 0 0.00136068 0 0.00136078 3.3 0.0013606999999999998 3.3 0.0013608 0 0.00136072 0 0.00136082 3.3 0.0013607399999999998 3.3 0.0013608399999999999 0 0.00136076 0 0.00136086 3.3 0.00136078 3.3 0.00136088 0 0.0013608 0 0.0013609 3.3 0.00136082 3.3 0.00136092 0 0.0013608399999999999 0 0.00136094 3.3 0.00136086 3.3 0.00136096 0 0.0013608799999999999 0 0.00136098 3.3 0.0013609 3.3 0.001361 0 0.0013609199999999998 0 0.00136102 3.3 0.00136094 3.3 0.00136104 0 0.0013609599999999998 0 0.0013610599999999999 3.3 0.00136098 3.3 0.00136108 0 0.001361 0 0.0013611 3.3 0.00136102 3.3 0.00136112 0 0.00136104 0 0.00136114 3.3 0.0013610599999999999 3.3 0.00136116 0 0.00136108 0 0.00136118 3.3 0.0013610999999999999 3.3 0.0013612 0 0.00136112 0 0.00136122 3.3 0.0013611399999999998 3.3 0.0013612399999999999 0 0.00136116 0 0.00136126 3.3 0.0013611799999999998 3.3 0.0013612799999999999 0 0.0013612 0 0.0013613 3.3 0.00136122 3.3 0.00136132 0 0.0013612399999999999 0 0.00136134 3.3 0.00136126 3.3 0.00136136 0 0.0013612799999999999 0 0.00136138 3.3 0.0013613 3.3 0.0013614 0 0.0013613199999999998 0 0.00136142 3.3 0.00136134 3.3 0.00136144 0 0.0013613599999999998 0 0.0013614599999999999 3.3 0.00136138 3.3 0.00136148 0 0.0013614 0 0.0013615 3.3 0.00136142 3.3 0.00136152 0 0.00136144 0 0.00136154 3.3 0.0013614599999999999 3.3 0.00136156 0 0.00136148 0 0.00136158 3.3 0.0013614999999999999 3.3 0.0013616 0 0.00136152 0 0.00136162 3.3 0.0013615399999999998 3.3 0.00136164 0 0.00136156 0 0.00136166 3.3 0.0013615799999999998 3.3 0.0013616799999999999 0 0.0013616 0 0.0013617 3.3 0.00136162 3.3 0.00136172 0 0.00136164 0 0.00136174 3.3 0.00136166 3.3 0.00136176 0 0.0013616799999999999 0 0.00136178 3.3 0.0013617 3.3 0.0013618 0 0.0013617199999999999 0 0.00136182 3.3 0.00136174 3.3 0.00136184 0 0.0013617599999999998 0 0.00136186 3.3 0.00136178 3.3 0.00136188 0 0.0013617999999999998 0 0.0013618999999999999 3.3 0.00136182 3.3 0.00136192 0 0.00136184 0 0.00136194 3.3 0.00136186 3.3 0.00136196 0 0.00136188 0 0.00136198 3.3 0.0013618999999999999 3.3 0.001362 0 0.00136192 0 0.00136202 3.3 0.0013619399999999999 3.3 0.00136204 0 0.00136196 0 0.00136206 3.3 0.0013619799999999998 3.3 0.0013620799999999999 0 0.001362 0 0.0013621 3.3 0.0013620199999999998 3.3 0.0013621199999999999 0 0.00136204 0 0.00136214 3.3 0.00136206 3.3 0.00136216 0 0.0013620799999999999 0 0.00136218 3.3 0.0013621 3.3 0.0013622 0 0.0013621199999999999 0 0.00136222 3.3 0.00136214 3.3 0.00136224 0 0.0013621599999999998 0 0.00136226 3.3 0.00136218 3.3 0.00136228 0 0.0013621999999999998 0 0.0013622999999999999 3.3 0.00136222 3.3 0.00136232 0 0.00136224 0 0.00136234 3.3 0.00136226 3.3 0.00136236 0 0.00136228 0 0.00136238 3.3 0.0013622999999999999 3.3 0.0013624 0 0.00136232 0 0.00136242 3.3 0.0013623399999999999 3.3 0.00136244 0 0.00136236 0 0.00136246 3.3 0.0013623799999999998 3.3 0.00136248 0 0.0013624 0 0.0013625 3.3 0.0013624199999999998 3.3 0.0013625199999999999 0 0.00136244 0 0.00136254 3.3 0.00136246 3.3 0.00136256 0 0.00136248 0 0.00136258 3.3 0.0013625 3.3 0.0013626 0 0.0013625199999999999 0 0.00136262 3.3 0.00136254 3.3 0.00136264 0 0.0013625599999999999 0 0.00136266 3.3 0.00136258 3.3 0.00136268 0 0.0013625999999999998 0 0.0013627 3.3 0.00136262 3.3 0.00136272 0 0.0013626399999999998 0 0.0013627399999999999 3.3 0.00136266 3.3 0.00136276 0 0.00136268 0 0.00136278 3.3 0.0013627 3.3 0.0013628 0 0.00136272 0 0.00136282 3.3 0.0013627399999999999 3.3 0.00136284 0 0.00136276 0 0.00136286 3.3 0.0013627799999999999 3.3 0.00136288 0 0.0013628 0 0.0013629 3.3 0.0013628199999999998 3.3 0.0013629199999999999 0 0.00136284 0 0.00136294 3.3 0.0013628599999999998 3.3 0.0013629599999999999 0 0.00136288 0 0.00136298 3.3 0.0013629 3.3 0.001363 0 0.0013629199999999999 0 0.00136302 3.3 0.00136294 3.3 0.00136304 0 0.0013629599999999999 0 0.00136306 3.3 0.00136298 3.3 0.00136308 0 0.0013629999999999998 0 0.0013631 3.3 0.00136302 3.3 0.00136312 0 0.0013630399999999998 0 0.0013631399999999999 3.3 0.00136306 3.3 0.00136316 0 0.00136308 0 0.00136318 3.3 0.0013631 3.3 0.0013632 0 0.00136312 0 0.00136322 3.3 0.0013631399999999999 3.3 0.00136324 0 0.00136316 0 0.00136326 3.3 0.0013631799999999999 3.3 0.00136328 0 0.0013632 0 0.0013633 3.3 0.0013632199999999998 3.3 0.00136332 0 0.00136324 0 0.00136334 3.3 0.0013632599999999998 3.3 0.0013633599999999999 0 0.00136328 0 0.00136338 3.3 0.0013633 3.3 0.0013634 0 0.00136332 0 0.00136342 3.3 0.00136334 3.3 0.00136344 0 0.0013633599999999999 0 0.00136346 3.3 0.00136338 3.3 0.00136348 0 0.0013633999999999999 0 0.0013635 3.3 0.00136342 3.3 0.00136352 0 0.0013634399999999998 0 0.0013635399999999999 3.3 0.00136346 3.3 0.00136356 0 0.0013634799999999998 0 0.0013635799999999999 3.3 0.0013635 3.3 0.0013636 0 0.00136352 0 0.00136362 3.3 0.0013635399999999999 3.3 0.00136364 0 0.00136356 0 0.00136366 3.3 0.0013635799999999999 3.3 0.00136368 0 0.0013636 0 0.0013637 3.3 0.0013636199999999998 3.3 0.00136372 0 0.00136364 0 0.00136374 3.3 0.0013636599999999998 3.3 0.0013637599999999999 0 0.00136368 0 0.00136378 3.3 0.0013636999999999998 3.3 0.0013637999999999999 0 0.00136372 0 0.00136382 3.3 0.00136374 3.3 0.00136384 0 0.0013637599999999999 0 0.00136386 3.3 0.00136378 3.3 0.00136388 0 0.0013637999999999999 0 0.0013639 3.3 0.00136382 3.3 0.00136392 0 0.0013638399999999998 0 0.00136394 3.3 0.00136386 3.3 0.00136396 0 0.0013638799999999998 0 0.0013639799999999999 3.3 0.0013639 3.3 0.001364 0 0.00136392 0 0.00136402 3.3 0.00136394 3.3 0.00136404 0 0.00136396 0 0.00136406 3.3 0.0013639799999999999 3.3 0.00136408 0 0.001364 0 0.0013641 3.3 0.0013640199999999999 3.3 0.00136412 0 0.00136404 0 0.00136414 3.3 0.0013640599999999998 3.3 0.00136416 0 0.00136408 0 0.00136418 3.3 0.0013640999999999998 3.3 0.0013641999999999999 0 0.00136412 0 0.00136422 3.3 0.00136414 3.3 0.00136424 0 0.00136416 0 0.00136426 3.3 0.00136418 3.3 0.00136428 0 0.0013641999999999999 0 0.0013643 3.3 0.00136422 3.3 0.00136432 0 0.0013642399999999999 0 0.00136434 3.3 0.00136426 3.3 0.00136436 0 0.0013642799999999998 0 0.0013643799999999999 3.3 0.0013643 3.3 0.0013644 0 0.0013643199999999998 0 0.0013644199999999999 3.3 0.00136434 3.3 0.00136444 0 0.00136436 0 0.00136446 3.3 0.0013643799999999999 3.3 0.00136448 0 0.0013644 0 0.0013645 3.3 0.0013644199999999999 3.3 0.00136452 0 0.00136444 0 0.00136454 3.3 0.0013644599999999998 3.3 0.00136456 0 0.00136448 0 0.00136458 3.3 0.0013644999999999998 3.3 0.0013645999999999999 0 0.00136452 0 0.00136462 3.3 0.00136454 3.3 0.00136464 0 0.00136456 0 0.00136466 3.3 0.00136458 3.3 0.00136468 0 0.0013645999999999999 0 0.0013647 3.3 0.00136462 3.3 0.00136472 0 0.0013646399999999999 0 0.00136474 3.3 0.00136466 3.3 0.00136476 0 0.0013646799999999998 0 0.00136478 3.3 0.0013647 3.3 0.0013648 0 0.0013647199999999998 0 0.0013648199999999999 3.3 0.00136474 3.3 0.00136484 0 0.00136476 0 0.00136486 3.3 0.00136478 3.3 0.00136488 0 0.0013648 0 0.0013649 3.3 0.0013648199999999999 3.3 0.00136492 0 0.00136484 0 0.00136494 3.3 0.0013648599999999999 3.3 0.00136496 0 0.00136488 0 0.00136498 3.3 0.0013648999999999998 3.3 0.001365 0 0.00136492 0 0.00136502 3.3 0.0013649399999999998 3.3 0.0013650399999999999 0 0.00136496 0 0.00136506 3.3 0.00136498 3.3 0.00136508 0 0.001365 0 0.0013651 3.3 0.00136502 3.3 0.00136512 0 0.0013650399999999999 0 0.00136514 3.3 0.00136506 3.3 0.00136516 0 0.0013650799999999999 0 0.00136518 3.3 0.0013651 3.3 0.0013652 0 0.0013651199999999998 0 0.0013652199999999999 3.3 0.00136514 3.3 0.00136524 0 0.0013651599999999998 0 0.0013652599999999999 3.3 0.00136518 3.3 0.00136528 0 0.0013652 0 0.0013653 3.3 0.0013652199999999999 3.3 0.00136532 0 0.00136524 0 0.00136534 3.3 0.0013652599999999999 3.3 0.00136536 0 0.00136528 0 0.00136538 3.3 0.0013652999999999998 3.3 0.0013654 0 0.00136532 0 0.00136542 3.3 0.0013653399999999998 3.3 0.0013654399999999999 0 0.00136536 0 0.00136546 3.3 0.00136538 3.3 0.00136548 0 0.0013654 0 0.0013655 3.3 0.00136542 3.3 0.00136552 0 0.0013654399999999999 0 0.00136554 3.3 0.00136546 3.3 0.00136556 0 0.0013654799999999999 0 0.00136558 3.3 0.0013655 3.3 0.0013656 0 0.0013655199999999998 0 0.00136562 3.3 0.00136554 3.3 0.00136564 0 0.0013655599999999998 0 0.0013656599999999999 3.3 0.00136558 3.3 0.00136568 0 0.0013656 0 0.0013657 3.3 0.00136562 3.3 0.00136572 0 0.00136564 0 0.00136574 3.3 0.0013656599999999999 3.3 0.00136576 0 0.00136568 0 0.00136578 3.3 0.0013656999999999999 3.3 0.0013658 0 0.00136572 0 0.00136582 3.3 0.0013657399999999998 3.3 0.00136584 0 0.00136576 0 0.00136586 3.3 0.0013657799999999998 3.3 0.0013658799999999999 0 0.0013658 0 0.0013659 3.3 0.00136582 3.3 0.00136592 0 0.00136584 0 0.00136594 3.3 0.00136586 3.3 0.00136596 0 0.0013658799999999999 0 0.00136598 3.3 0.0013659 3.3 0.001366 0 0.0013659199999999999 0 0.00136602 3.3 0.00136594 3.3 0.00136604 0 0.0013659599999999998 0 0.0013660599999999999 3.3 0.00136598 3.3 0.00136608 0 0.0013659999999999998 0 0.0013660999999999999 3.3 0.00136602 3.3 0.00136612 0 0.00136604 0 0.00136614 3.3 0.0013660599999999999 3.3 0.00136616 0 0.00136608 0 0.00136618 3.3 0.0013660999999999999 3.3 0.0013662 0 0.00136612 0 0.00136622 3.3 0.0013661399999999998 3.3 0.00136624 0 0.00136616 0 0.00136626 3.3 0.0013661799999999998 3.3 0.0013662799999999999 0 0.0013662 0 0.0013663 3.3 0.00136622 3.3 0.00136632 0 0.00136624 0 0.00136634 3.3 0.00136626 3.3 0.00136636 0 0.0013662799999999999 0 0.00136638 3.3 0.0013663 3.3 0.0013664 0 0.0013663199999999999 0 0.00136642 3.3 0.00136634 3.3 0.00136644 0 0.0013663599999999998 0 0.00136646 3.3 0.00136638 3.3 0.00136648 0 0.0013663999999999998 0 0.0013664999999999999 3.3 0.00136642 3.3 0.00136652 0 0.00136644 0 0.00136654 3.3 0.00136646 3.3 0.00136656 0 0.00136648 0 0.00136658 3.3 0.0013664999999999999 3.3 0.0013666 0 0.00136652 0 0.00136662 3.3 0.0013665399999999999 3.3 0.00136664 0 0.00136656 0 0.00136666 3.3 0.0013665799999999998 3.3 0.0013666799999999999 0 0.0013666 0 0.0013667 3.3 0.0013666199999999998 3.3 0.0013667199999999999 0 0.00136664 0 0.00136674 3.3 0.00136666 3.3 0.00136676 0 0.0013666799999999999 0 0.00136678 3.3 0.0013667 3.3 0.0013668 0 0.0013667199999999999 0 0.00136682 3.3 0.00136674 3.3 0.00136684 0 0.0013667599999999999 0 0.00136686 3.3 0.00136678 3.3 0.00136688 0 0.0013667999999999998 0 0.0013668999999999999 3.3 0.00136682 3.3 0.00136692 0 0.0013668399999999998 0 0.0013669399999999999 3.3 0.00136686 3.3 0.00136696 0 0.00136688 0 0.00136698 3.3 0.0013668999999999999 3.3 0.001367 0 0.00136692 0 0.00136702 3.3 0.0013669399999999999 3.3 0.00136704 0 0.00136696 0 0.00136706 3.3 0.0013669799999999998 3.3 0.00136708 0 0.001367 0 0.0013671 3.3 0.0013670199999999998 3.3 0.0013671199999999999 0 0.00136704 0 0.00136714 3.3 0.00136706 3.3 0.00136716 0 0.00136708 0 0.00136718 3.3 0.0013671 3.3 0.0013672 0 0.0013671199999999999 0 0.00136722 3.3 0.00136714 3.3 0.00136724 0 0.0013671599999999999 0 0.00136726 3.3 0.00136718 3.3 0.00136728 0 0.0013671999999999998 0 0.0013673 3.3 0.00136722 3.3 0.00136732 0 0.0013672399999999998 0 0.0013673399999999999 3.3 0.00136726 3.3 0.00136736 0 0.00136728 0 0.00136738 3.3 0.0013673 3.3 0.0013674 0 0.00136732 0 0.00136742 3.3 0.0013673399999999999 3.3 0.00136744 0 0.00136736 0 0.00136746 3.3 0.0013673799999999999 3.3 0.00136748 0 0.0013674 0 0.0013675 3.3 0.0013674199999999998 3.3 0.0013675199999999999 0 0.00136744 0 0.00136754 3.3 0.0013674599999999998 3.3 0.0013675599999999999 0 0.00136748 0 0.00136758 3.3 0.0013675 3.3 0.0013676 0 0.0013675199999999999 0 0.00136762 3.3 0.00136754 3.3 0.00136764 0 0.0013675599999999999 0 0.00136766 3.3 0.00136758 3.3 0.00136768 0 0.0013675999999999998 0 0.0013677 3.3 0.00136762 3.3 0.00136772 0 0.0013676399999999998 0 0.0013677399999999999 3.3 0.00136766 3.3 0.00136776 0 0.00136768 0 0.00136778 3.3 0.0013677 3.3 0.0013678 0 0.00136772 0 0.00136782 3.3 0.0013677399999999999 3.3 0.00136784 0 0.00136776 0 0.00136786 3.3 0.0013677799999999999 3.3 0.00136788 0 0.0013678 0 0.0013679 3.3 0.0013678199999999998 3.3 0.00136792 0 0.00136784 0 0.00136794 3.3 0.0013678599999999998 3.3 0.0013679599999999999 0 0.00136788 0 0.00136798 3.3 0.0013679 3.3 0.001368 0 0.00136792 0 0.00136802 3.3 0.00136794 3.3 0.00136804 0 0.0013679599999999999 0 0.00136806 3.3 0.00136798 3.3 0.00136808 0 0.0013679999999999999 0 0.0013681 3.3 0.00136802 3.3 0.00136812 0 0.0013680399999999998 0 0.00136814 3.3 0.00136806 3.3 0.00136816 0 0.0013680799999999998 0 0.0013681799999999999 3.3 0.0013681 3.3 0.0013682 0 0.00136812 0 0.00136822 3.3 0.00136814 3.3 0.00136824 0 0.00136816 0 0.00136826 3.3 0.0013681799999999999 3.3 0.00136828 0 0.0013682 0 0.0013683 3.3 0.0013682199999999999 3.3 0.00136832 0 0.00136824 0 0.00136834 3.3 0.0013682599999999998 3.3 0.0013683599999999999 0 0.00136828 0 0.00136838 3.3 0.0013682999999999998 3.3 0.0013683999999999999 0 0.00136832 0 0.00136842 3.3 0.00136834 3.3 0.00136844 0 0.0013683599999999999 0 0.00136846 3.3 0.00136838 3.3 0.00136848 0 0.0013683999999999999 0 0.0013685 3.3 0.00136842 3.3 0.00136852 0 0.0013684399999999998 0 0.00136854 3.3 0.00136846 3.3 0.00136856 0 0.0013684799999999998 0 0.0013685799999999999 3.3 0.0013685 3.3 0.0013686 0 0.00136852 0 0.00136862 3.3 0.00136854 3.3 0.00136864 0 0.00136856 0 0.00136866 3.3 0.0013685799999999999 3.3 0.00136868 0 0.0013686 0 0.0013687 3.3 0.0013686199999999999 3.3 0.00136872 0 0.00136864 0 0.00136874 3.3 0.0013686599999999998 3.3 0.00136876 0 0.00136868 0 0.00136878 3.3 0.0013686999999999998 3.3 0.0013687999999999999 0 0.00136872 0 0.00136882 3.3 0.00136874 3.3 0.00136884 0 0.00136876 0 0.00136886 3.3 0.00136878 3.3 0.00136888 0 0.0013687999999999999 0 0.0013689 3.3 0.00136882 3.3 0.00136892 0 0.0013688399999999999 0 0.00136894 3.3 0.00136886 3.3 0.00136896 0 0.0013688799999999998 0 0.00136898 3.3 0.0013689 3.3 0.001369 0 0.0013689199999999998 0 0.0013690199999999999 3.3 0.00136894 3.3 0.00136904 0 0.00136896 0 0.00136906 3.3 0.00136898 3.3 0.00136908 0 0.001369 0 0.0013691 3.3 0.0013690199999999999 3.3 0.00136912 0 0.00136904 0 0.00136914 3.3 0.0013690599999999999 3.3 0.00136916 0 0.00136908 0 0.00136918 3.3 0.0013690999999999998 3.3 0.0013691999999999999 0 0.00136912 0 0.00136922 3.3 0.0013691399999999998 3.3 0.0013692399999999999 0 0.00136916 0 0.00136926 3.3 0.00136918 3.3 0.00136928 0 0.0013691999999999999 0 0.0013693 3.3 0.00136922 3.3 0.00136932 0 0.0013692399999999999 0 0.00136934 3.3 0.00136926 3.3 0.00136936 0 0.0013692799999999998 0 0.00136938 3.3 0.0013693 3.3 0.0013694 0 0.0013693199999999998 0 0.0013694199999999999 3.3 0.00136934 3.3 0.00136944 0 0.00136936 0 0.00136946 3.3 0.00136938 3.3 0.00136948 0 0.0013694 0 0.0013695 3.3 0.0013694199999999999 3.3 0.00136952 0 0.00136944 0 0.00136954 3.3 0.0013694599999999999 3.3 0.00136956 0 0.00136948 0 0.00136958 3.3 0.0013694999999999998 3.3 0.0013696 0 0.00136952 0 0.00136962 3.3 0.0013695399999999998 3.3 0.0013696399999999999 0 0.00136956 0 0.00136966 3.3 0.00136958 3.3 0.00136968 0 0.0013696 0 0.0013697 3.3 0.00136962 3.3 0.00136972 0 0.0013696399999999999 0 0.00136974 3.3 0.00136966 3.3 0.00136976 0 0.0013696799999999999 0 0.00136978 3.3 0.0013697 3.3 0.0013698 0 0.0013697199999999998 0 0.00136982 3.3 0.00136974 3.3 0.00136984 0 0.0013697599999999998 0 0.0013698599999999999 3.3 0.00136978 3.3 0.00136988 0 0.0013698 0 0.0013699 3.3 0.00136982 3.3 0.00136992 0 0.00136984 0 0.00136994 3.3 0.0013698599999999999 3.3 0.00136996 0 0.00136988 0 0.00136998 3.3 0.0013698999999999999 3.3 0.00137 0 0.00136992 0 0.00137002 3.3 0.0013699399999999998 3.3 0.0013700399999999999 0 0.00136996 0 0.00137006 3.3 0.0013699799999999998 3.3 0.0013700799999999999 0 0.00137 0 0.0013701 3.3 0.00137002 3.3 0.00137012 0 0.0013700399999999999 0 0.00137014 3.3 0.00137006 3.3 0.00137016 0 0.0013700799999999999 0 0.00137018 3.3 0.0013701 3.3 0.0013702 0 0.0013701199999999998 0 0.00137022 3.3 0.00137014 3.3 0.00137024 0 0.0013701599999999998 0 0.0013702599999999999 3.3 0.00137018 3.3 0.00137028 0 0.0013702 0 0.0013703 3.3 0.00137022 3.3 0.00137032 0 0.00137024 0 0.00137034 3.3 0.0013702599999999999 3.3 0.00137036 0 0.00137028 0 0.00137038 3.3 0.0013702999999999999 3.3 0.0013704 0 0.00137032 0 0.00137042 3.3 0.0013703399999999998 3.3 0.00137044 0 0.00137036 0 0.00137046 3.3 0.0013703799999999998 3.3 0.0013704799999999999 0 0.0013704 0 0.0013705 3.3 0.00137042 3.3 0.00137052 0 0.00137044 0 0.00137054 3.3 0.00137046 3.3 0.00137056 0 0.0013704799999999999 0 0.00137058 3.3 0.0013705 3.3 0.0013706 0 0.0013705199999999999 0 0.00137062 3.3 0.00137054 3.3 0.00137064 0 0.0013705599999999998 0 0.0013706599999999999 3.3 0.00137058 3.3 0.00137068 0 0.0013705999999999998 0 0.0013706999999999999 3.3 0.00137062 3.3 0.00137072 0 0.00137064 0 0.00137074 3.3 0.0013706599999999999 3.3 0.00137076 0 0.00137068 0 0.00137078 3.3 0.0013706999999999999 3.3 0.0013708 0 0.00137072 0 0.00137082 3.3 0.0013707399999999998 3.3 0.00137084 0 0.00137076 0 0.00137086 3.3 0.0013707799999999998 3.3 0.0013708799999999999 0 0.0013708 0 0.0013709 3.3 0.0013708199999999998 3.3 0.0013709199999999999 0 0.00137084 0 0.00137094 3.3 0.00137086 3.3 0.00137096 0 0.0013708799999999999 0 0.00137098 3.3 0.0013709 3.3 0.001371 0 0.0013709199999999999 0 0.00137102 3.3 0.00137094 3.3 0.00137104 0 0.0013709599999999998 0 0.00137106 3.3 0.00137098 3.3 0.00137108 0 0.0013709999999999998 0 0.0013710999999999999 3.3 0.00137102 3.3 0.00137112 0 0.00137104 0 0.00137114 3.3 0.00137106 3.3 0.00137116 0 0.00137108 0 0.00137118 3.3 0.0013710999999999999 3.3 0.0013712 0 0.00137112 0 0.00137122 3.3 0.0013711399999999999 3.3 0.00137124 0 0.00137116 0 0.00137126 3.3 0.0013711799999999998 3.3 0.00137128 0 0.0013712 0 0.0013713 3.3 0.0013712199999999998 3.3 0.0013713199999999999 0 0.00137124 0 0.00137134 3.3 0.00137126 3.3 0.00137136 0 0.00137128 0 0.00137138 3.3 0.0013713 3.3 0.0013714 0 0.0013713199999999999 0 0.00137142 3.3 0.00137134 3.3 0.00137144 0 0.0013713599999999999 0 0.00137146 3.3 0.00137138 3.3 0.00137148 0 0.0013713999999999998 0 0.0013714999999999999 3.3 0.00137142 3.3 0.00137152 0 0.0013714399999999998 0 0.0013715399999999999 3.3 0.00137146 3.3 0.00137156 0 0.00137148 0 0.00137158 3.3 0.0013714999999999999 3.3 0.0013716 0 0.00137152 0 0.00137162 3.3 0.0013715399999999999 3.3 0.00137164 0 0.00137156 0 0.00137166 3.3 0.0013715799999999998 3.3 0.00137168 0 0.0013716 0 0.0013717 3.3 0.0013716199999999998 3.3 0.0013717199999999999 0 0.00137164 0 0.00137174 3.3 0.00137166 3.3 0.00137176 0 0.00137168 0 0.00137178 3.3 0.0013717 3.3 0.0013718 0 0.0013717199999999999 0 0.00137182 3.3 0.00137174 3.3 0.00137184 0 0.0013717599999999999 0 0.00137186 3.3 0.00137178 3.3 0.00137188 0 0.0013717999999999998 0 0.0013719 3.3 0.00137182 3.3 0.00137192 0 0.0013718399999999998 0 0.0013719399999999999 3.3 0.00137186 3.3 0.00137196 0 0.00137188 0 0.00137198 3.3 0.0013719 3.3 0.001372 0 0.00137192 0 0.00137202 3.3 0.0013719399999999999 3.3 0.00137204 0 0.00137196 0 0.00137206 3.3 0.0013719799999999999 3.3 0.00137208 0 0.001372 0 0.0013721 3.3 0.0013720199999999998 3.3 0.00137212 0 0.00137204 0 0.00137214 3.3 0.0013720599999999998 3.3 0.0013721599999999999 0 0.00137208 0 0.00137218 3.3 0.0013721 3.3 0.0013722 0 0.00137212 0 0.00137222 3.3 0.00137214 3.3 0.00137224 0 0.0013721599999999999 0 0.00137226 3.3 0.00137218 3.3 0.00137228 0 0.0013721999999999999 0 0.0013723 3.3 0.00137222 3.3 0.00137232 0 0.0013722399999999998 0 0.0013723399999999999 3.3 0.00137226 3.3 0.00137236 0 0.0013722799999999998 0 0.0013723799999999999 3.3 0.0013723 3.3 0.0013724 0 0.00137232 0 0.00137242 3.3 0.0013723399999999999 3.3 0.00137244 0 0.00137236 0 0.00137246 3.3 0.0013723799999999999 3.3 0.00137248 0 0.0013724 0 0.0013725 3.3 0.0013724199999999998 3.3 0.00137252 0 0.00137244 0 0.00137254 3.3 0.0013724599999999998 3.3 0.0013725599999999999 0 0.00137248 0 0.00137258 3.3 0.0013725 3.3 0.0013726 0 0.00137252 0 0.00137262 3.3 0.00137254 3.3 0.00137264 0 0.0013725599999999999 0 0.00137266 3.3 0.00137258 3.3 0.00137268 0 0.0013725999999999999 0 0.0013727 3.3 0.00137262 3.3 0.00137272 0 0.0013726399999999998 0 0.00137274 3.3 0.00137266 3.3 0.00137276 0 0.0013726799999999998 0 0.0013727799999999999 3.3 0.0013727 3.3 0.0013728 0 0.00137272 0 0.00137282 3.3 0.00137274 3.3 0.00137284 0 0.00137276 0 0.00137286 3.3 0.0013727799999999999 3.3 0.00137288 0 0.0013728 0 0.0013729 3.3 0.0013728199999999999 3.3 0.00137292 0 0.00137284 0 0.00137294 3.3 0.0013728599999999998 3.3 0.00137296 0 0.00137288 0 0.00137298 3.3 0.0013728999999999998 3.3 0.0013729999999999999 0 0.00137292 0 0.00137302 3.3 0.00137294 3.3 0.00137304 0 0.00137296 0 0.00137306 3.3 0.00137298 3.3 0.00137308 0 0.0013729999999999999 0 0.0013731 3.3 0.00137302 3.3 0.00137312 0 0.0013730399999999999 0 0.00137314 3.3 0.00137306 3.3 0.00137316 0 0.0013730799999999998 0 0.0013731799999999999 3.3 0.0013731 3.3 0.0013732 0 0.0013731199999999998 0 0.0013732199999999999 3.3 0.00137314 3.3 0.00137324 0 0.00137316 0 0.00137326 3.3 0.0013731799999999999 3.3 0.00137328 0 0.0013732 0 0.0013733 3.3 0.0013732199999999999 3.3 0.00137332 0 0.00137324 0 0.00137334 3.3 0.0013732599999999998 3.3 0.00137336 0 0.00137328 0 0.00137338 3.3 0.0013732999999999998 3.3 0.0013733999999999999 0 0.00137332 0 0.00137342 3.3 0.00137334 3.3 0.00137344 0 0.00137336 0 0.00137346 3.3 0.00137338 3.3 0.00137348 0 0.0013733999999999999 0 0.0013735 3.3 0.00137342 3.3 0.00137352 0 0.0013734399999999999 0 0.00137354 3.3 0.00137346 3.3 0.00137356 0 0.0013734799999999998 0 0.00137358 3.3 0.0013735 3.3 0.0013736 0 0.0013735199999999998 0 0.0013736199999999999 3.3 0.00137354 3.3 0.00137364 0 0.00137356 0 0.00137366 3.3 0.00137358 3.3 0.00137368 0 0.0013736 0 0.0013737 3.3 0.0013736199999999999 3.3 0.00137372 0 0.00137364 0 0.00137374 3.3 0.0013736599999999999 3.3 0.00137376 0 0.00137368 0 0.00137378 3.3 0.0013736999999999998 3.3 0.0013737999999999999 0 0.00137372 0 0.00137382 3.3 0.0013737399999999998 3.3 0.0013738399999999999 0 0.00137376 0 0.00137386 3.3 0.00137378 3.3 0.00137388 0 0.0013737999999999999 0 0.0013739 3.3 0.00137382 3.3 0.00137392 0 0.0013738399999999999 0 0.00137394 3.3 0.00137386 3.3 0.00137396 0 0.0013738799999999998 0 0.00137398 3.3 0.0013739 3.3 0.001374 0 0.0013739199999999998 0 0.0013740199999999999 3.3 0.00137394 3.3 0.00137404 0 0.0013739599999999998 0 0.0013740599999999999 3.3 0.00137398 3.3 0.00137408 0 0.001374 0 0.0013741 3.3 0.0013740199999999999 3.3 0.00137412 0 0.00137404 0 0.00137414 3.3 0.0013740599999999999 3.3 0.00137416 0 0.00137408 0 0.00137418 3.3 0.0013740999999999998 3.3 0.0013742 0 0.00137412 0 0.00137422 3.3 0.0013741399999999998 3.3 0.0013742399999999999 0 0.00137416 0 0.00137426 3.3 0.00137418 3.3 0.00137428 0 0.0013742 0 0.0013743 3.3 0.00137422 3.3 0.00137432 0 0.0013742399999999999 0 0.00137434 3.3 0.00137426 3.3 0.00137436 0 0.0013742799999999999 0 0.00137438 3.3 0.0013743 3.3 0.0013744 0 0.0013743199999999998 0 0.00137442 3.3 0.00137434 3.3 0.00137444 0 0.0013743599999999998 0 0.0013744599999999999 3.3 0.00137438 3.3 0.00137448 0 0.0013744 0 0.0013745 3.3 0.00137442 3.3 0.00137452 0 0.00137444 0 0.00137454 3.3 0.0013744599999999999 3.3 0.00137456 0 0.00137448 0 0.00137458 3.3 0.0013744999999999999 3.3 0.0013746 0 0.00137452 0 0.00137462 3.3 0.0013745399999999998 3.3 0.0013746399999999999 0 0.00137456 0 0.00137466 3.3 0.0013745799999999998 3.3 0.0013746799999999999 0 0.0013746 0 0.0013747 3.3 0.00137462 3.3 0.00137472 0 0.0013746399999999999 0 0.00137474 3.3 0.00137466 3.3 0.00137476 0 0.0013746799999999999 0 0.00137478 3.3 0.0013747 3.3 0.0013748 0 0.0013747199999999998 0 0.00137482 3.3 0.00137474 3.3 0.00137484 0 0.0013747599999999998 0 0.0013748599999999999 3.3 0.00137478 3.3 0.00137488 0 0.0013748 0 0.0013749 3.3 0.00137482 3.3 0.00137492 0 0.00137484 0 0.00137494 3.3 0.0013748599999999999 3.3 0.00137496 0 0.00137488 0 0.00137498 3.3 0.0013748999999999999 3.3 0.001375 0 0.00137492 0 0.00137502 3.3 0.0013749399999999998 3.3 0.00137504 0 0.00137496 0 0.00137506 3.3 0.0013749799999999998 3.3 0.0013750799999999999 0 0.001375 0 0.0013751 3.3 0.00137502 3.3 0.00137512 0 0.00137504 0 0.00137514 3.3 0.00137506 3.3 0.00137516 0 0.0013750799999999999 0 0.00137518 3.3 0.0013751 3.3 0.0013752 0 0.0013751199999999999 0 0.00137522 3.3 0.00137514 3.3 0.00137524 0 0.0013751599999999998 0 0.00137526 3.3 0.00137518 3.3 0.00137528 0 0.0013751999999999998 0 0.0013752999999999999 3.3 0.00137522 3.3 0.00137532 0 0.00137524 0 0.00137534 3.3 0.00137526 3.3 0.00137536 0 0.00137528 0 0.00137538 3.3 0.0013752999999999999 3.3 0.0013754 0 0.00137532 0 0.00137542 3.3 0.0013753399999999999 3.3 0.00137544 0 0.00137536 0 0.00137546 3.3 0.0013753799999999998 3.3 0.0013754799999999999 0 0.0013754 0 0.0013755 3.3 0.0013754199999999998 3.3 0.0013755199999999999 0 0.00137544 0 0.00137554 3.3 0.00137546 3.3 0.00137556 0 0.0013754799999999999 0 0.00137558 3.3 0.0013755 3.3 0.0013756 0 0.0013755199999999999 0 0.00137562 3.3 0.00137554 3.3 0.00137564 0 0.0013755599999999998 0 0.00137566 3.3 0.00137558 3.3 0.00137568 0 0.0013755999999999998 0 0.0013756999999999999 3.3 0.00137562 3.3 0.00137572 0 0.00137564 0 0.00137574 3.3 0.00137566 3.3 0.00137576 0 0.00137568 0 0.00137578 3.3 0.0013756999999999999 3.3 0.0013758 0 0.00137572 0 0.00137582 3.3 0.0013757399999999999 3.3 0.00137584 0 0.00137576 0 0.00137586 3.3 0.0013757799999999998 3.3 0.00137588 0 0.0013758 0 0.0013759 3.3 0.0013758199999999998 3.3 0.0013759199999999999 0 0.00137584 0 0.00137594 3.3 0.00137586 3.3 0.00137596 0 0.00137588 0 0.00137598 3.3 0.0013759 3.3 0.001376 0 0.0013759199999999999 0 0.00137602 3.3 0.00137594 3.3 0.00137604 0 0.0013759599999999999 0 0.00137606 3.3 0.00137598 3.3 0.00137608 0 0.0013759999999999998 0 0.0013761 3.3 0.00137602 3.3 0.00137612 0 0.0013760399999999998 0 0.0013761399999999999 3.3 0.00137606 3.3 0.00137616 0 0.00137608 0 0.00137618 3.3 0.0013761 3.3 0.0013762 0 0.00137612 0 0.00137622 3.3 0.0013761399999999999 3.3 0.00137624 0 0.00137616 0 0.00137626 3.3 0.0013761799999999999 3.3 0.00137628 0 0.0013762 0 0.0013763 3.3 0.0013762199999999998 3.3 0.0013763199999999999 0 0.00137624 0 0.00137634 3.3 0.0013762599999999998 3.3 0.0013763599999999999 0 0.00137628 0 0.00137638 3.3 0.0013763 3.3 0.0013764 0 0.0013763199999999999 0 0.00137642 3.3 0.00137634 3.3 0.00137644 0 0.0013763599999999999 0 0.00137646 3.3 0.00137638 3.3 0.00137648 0 0.0013763999999999998 0 0.0013765 3.3 0.00137642 3.3 0.00137652 0 0.0013764399999999998 0 0.0013765399999999999 3.3 0.00137646 3.3 0.00137656 0 0.00137648 0 0.00137658 3.3 0.0013765 3.3 0.0013766 0 0.00137652 0 0.00137662 3.3 0.0013765399999999999 3.3 0.00137664 0 0.00137656 0 0.00137666 3.3 0.0013765799999999999 3.3 0.00137668 0 0.0013766 0 0.0013767 3.3 0.0013766199999999998 3.3 0.00137672 0 0.00137664 0 0.00137674 3.3 0.0013766599999999998 3.3 0.0013767599999999999 0 0.00137668 0 0.00137678 3.3 0.0013767 3.3 0.0013768 0 0.00137672 0 0.00137682 3.3 0.00137674 3.3 0.00137684 0 0.0013767599999999999 0 0.00137686 3.3 0.00137678 3.3 0.00137688 0 0.0013767999999999999 0 0.0013769 3.3 0.00137682 3.3 0.00137692 0 0.0013768399999999998 0 0.0013769399999999999 3.3 0.00137686 3.3 0.00137696 0 0.0013768799999999998 0 0.0013769799999999999 3.3 0.0013769 3.3 0.001377 0 0.00137692 0 0.00137702 3.3 0.0013769399999999999 3.3 0.00137704 0 0.00137696 0 0.00137706 3.3 0.0013769799999999999 3.3 0.00137708 0 0.001377 0 0.0013771 3.3 0.0013770199999999999 3.3 0.00137712 0 0.00137704 0 0.00137714 3.3 0.0013770599999999998 3.3 0.0013771599999999999 0 0.00137708 0 0.00137718 3.3 0.0013770999999999998 3.3 0.0013771999999999999 0 0.00137712 0 0.00137722 3.3 0.00137714 3.3 0.00137724 0 0.0013771599999999999 0 0.00137726 3.3 0.00137718 3.3 0.00137728 0 0.0013771999999999999 0 0.0013773 3.3 0.00137722 3.3 0.00137732 0 0.0013772399999999998 0 0.00137734 3.3 0.00137726 3.3 0.00137736 0 0.0013772799999999998 0 0.0013773799999999999 3.3 0.0013773 3.3 0.0013774 0 0.00137732 0 0.00137742 3.3 0.00137734 3.3 0.00137744 0 0.00137736 0 0.00137746 3.3 0.0013773799999999999 3.3 0.00137748 0 0.0013774 0 0.0013775 3.3 0.0013774199999999999 3.3 0.00137752 0 0.00137744 0 0.00137754 3.3 0.0013774599999999998 3.3 0.00137756 0 0.00137748 0 0.00137758 3.3 0.0013774999999999998 3.3 0.0013775999999999999 0 0.00137752 0 0.00137762 3.3 0.00137754 3.3 0.00137764 0 0.00137756 0 0.00137766 3.3 0.00137758 3.3 0.00137768 0 0.0013775999999999999 0 0.0013777 3.3 0.00137762 3.3 0.00137772 0 0.0013776399999999999 0 0.00137774 3.3 0.00137766 3.3 0.00137776 0 0.0013776799999999998 0 0.0013777799999999999 3.3 0.0013777 3.3 0.0013778 0 0.0013777199999999998 0 0.0013778199999999999 3.3 0.00137774 3.3 0.00137784 0 0.00137776 0 0.00137786 3.3 0.0013777799999999999 3.3 0.00137788 0 0.0013778 0 0.0013779 3.3 0.0013778199999999999 3.3 0.00137792 0 0.00137784 0 0.00137794 3.3 0.0013778599999999998 3.3 0.00137796 0 0.00137788 0 0.00137798 3.3 0.0013778999999999998 3.3 0.0013779999999999999 0 0.00137792 0 0.00137802 3.3 0.0013779399999999998 3.3 0.0013780399999999999 0 0.00137796 0 0.00137806 3.3 0.00137798 3.3 0.00137808 0 0.0013779999999999999 0 0.0013781 3.3 0.00137802 3.3 0.00137812 0 0.0013780399999999999 0 0.00137814 3.3 0.00137806 3.3 0.00137816 0 0.0013780799999999998 0 0.00137818 3.3 0.0013781 3.3 0.0013782 0 0.0013781199999999998 0 0.0013782199999999999 3.3 0.00137814 3.3 0.00137824 0 0.00137816 0 0.00137826 3.3 0.00137818 3.3 0.00137828 0 0.0013782 0 0.0013783 3.3 0.0013782199999999999 3.3 0.00137832 0 0.00137824 0 0.00137834 3.3 0.0013782599999999999 3.3 0.00137836 0 0.00137828 0 0.00137838 3.3 0.0013782999999999998 3.3 0.0013784 0 0.00137832 0 0.00137842 3.3 0.0013783399999999998 3.3 0.0013784399999999999 0 0.00137836 0 0.00137846 3.3 0.00137838 3.3 0.00137848 0 0.0013784 0 0.0013785 3.3 0.00137842 3.3 0.00137852 0 0.0013784399999999999 0 0.00137854 3.3 0.00137846 3.3 0.00137856 0 0.0013784799999999999 0 0.00137858 3.3 0.0013785 3.3 0.0013786 0 0.0013785199999999998 0 0.0013786199999999999 3.3 0.00137854 3.3 0.00137864 0 0.0013785599999999998 0 0.0013786599999999999 3.3 0.00137858 3.3 0.00137868 0 0.0013786 0 0.0013787 3.3 0.0013786199999999999 3.3 0.00137872 0 0.00137864 0 0.00137874 3.3 0.0013786599999999999 3.3 0.00137876 0 0.00137868 0 0.00137878 3.3 0.0013786999999999998 3.3 0.0013788 0 0.00137872 0 0.00137882 3.3 0.0013787399999999998 3.3 0.0013788399999999999 0 0.00137876 0 0.00137886 3.3 0.00137878 3.3 0.00137888 0 0.0013788 0 0.0013789 3.3 0.00137882 3.3 0.00137892 0 0.0013788399999999999 0 0.00137894 3.3 0.00137886 3.3 0.00137896 0 0.0013788799999999999 0 0.00137898 3.3 0.0013789 3.3 0.001379 0 0.0013789199999999998 0 0.00137902 3.3 0.00137894 3.3 0.00137904 0 0.0013789599999999998 0 0.0013790599999999999 3.3 0.00137898 3.3 0.00137908 0 0.001379 0 0.0013791 3.3 0.00137902 3.3 0.00137912 0 0.00137904 0 0.00137914 3.3 0.0013790599999999999 3.3 0.00137916 0 0.00137908 0 0.00137918 3.3 0.0013790999999999999 3.3 0.0013792 0 0.00137912 0 0.00137922 3.3 0.0013791399999999998 3.3 0.00137924 0 0.00137916 0 0.00137926 3.3 0.0013791799999999998 3.3 0.0013792799999999999 0 0.0013792 0 0.0013793 3.3 0.00137922 3.3 0.00137932 0 0.00137924 0 0.00137934 3.3 0.00137926 3.3 0.00137936 0 0.0013792799999999999 0 0.00137938 3.3 0.0013793 3.3 0.0013794 0 0.0013793199999999999 0 0.00137942 3.3 0.00137934 3.3 0.00137944 0 0.0013793599999999998 0 0.0013794599999999999 3.3 0.00137938 3.3 0.00137948 0 0.0013793999999999998 0 0.0013794999999999999 3.3 0.00137942 3.3 0.00137952 0 0.00137944 0 0.00137954 3.3 0.0013794599999999999 3.3 0.00137956 0 0.00137948 0 0.00137958 3.3 0.0013794999999999999 3.3 0.0013796 0 0.00137952 0 0.00137962 3.3 0.0013795399999999998 3.3 0.00137964 0 0.00137956 0 0.00137966 3.3 0.0013795799999999998 3.3 0.0013796799999999999 0 0.0013796 0 0.0013797 3.3 0.00137962 3.3 0.00137972 0 0.00137964 0 0.00137974 3.3 0.00137966 3.3 0.00137976 0 0.0013796799999999999 0 0.00137978 3.3 0.0013797 3.3 0.0013798 0 0.0013797199999999999 0 0.00137982 3.3 0.00137974 3.3 0.00137984 0 0.0013797599999999998 0 0.00137986 3.3 0.00137978 3.3 0.00137988 0 0.0013797999999999998 0 0.0013798999999999999 3.3 0.00137982 3.3 0.00137992 0 0.00137984 0 0.00137994 3.3 0.00137986 3.3 0.00137996 0 0.00137988 0 0.00137998 3.3 0.0013798999999999999 3.3 0.00138 0 0.00137992 0 0.00138002 3.3 0.0013799399999999999 3.3 0.00138004 0 0.00137996 0 0.00138006 3.3 0.0013799799999999998 3.3 0.00138008 0 0.00138 0 0.0013801 3.3 0.0013800199999999998 3.3 0.0013801199999999999 0 0.00138004 0 0.00138014 3.3 0.00138006 3.3 0.00138016 0 0.00138008 0 0.00138018 3.3 0.0013801 3.3 0.0013802 0 0.0013801199999999999 0 0.00138022 3.3 0.00138014 3.3 0.00138024 0 0.0013801599999999999 0 0.00138026 3.3 0.00138018 3.3 0.00138028 0 0.0013801999999999998 0 0.0013802999999999999 3.3 0.00138022 3.3 0.00138032 0 0.0013802399999999998 0 0.0013803399999999999 3.3 0.00138026 3.3 0.00138036 0 0.00138028 0 0.00138038 3.3 0.0013802999999999999 3.3 0.0013804 0 0.00138032 0 0.00138042 3.3 0.0013803399999999999 3.3 0.00138044 0 0.00138036 0 0.00138046 3.3 0.0013803799999999998 3.3 0.00138048 0 0.0013804 0 0.0013805 3.3 0.0013804199999999998 3.3 0.0013805199999999999 0 0.00138044 0 0.00138054 3.3 0.00138046 3.3 0.00138056 0 0.00138048 0 0.00138058 3.3 0.0013805 3.3 0.0013806 0 0.0013805199999999999 0 0.00138062 3.3 0.00138054 3.3 0.00138064 0 0.0013805599999999999 0 0.00138066 3.3 0.00138058 3.3 0.00138068 0 0.0013805999999999998 0 0.0013807 3.3 0.00138062 3.3 0.00138072 0 0.0013806399999999998 0 0.0013807399999999999 3.3 0.00138066 3.3 0.00138076 0 0.00138068 0 0.00138078 3.3 0.0013807 3.3 0.0013808 0 0.00138072 0 0.00138082 3.3 0.0013807399999999999 3.3 0.00138084 0 0.00138076 0 0.00138086 3.3 0.0013807799999999999 3.3 0.00138088 0 0.0013808 0 0.0013809 3.3 0.0013808199999999998 3.3 0.0013809199999999999 0 0.00138084 0 0.00138094 3.3 0.0013808599999999998 3.3 0.0013809599999999999 0 0.00138088 0 0.00138098 3.3 0.0013809 3.3 0.001381 0 0.0013809199999999999 0 0.00138102 3.3 0.00138094 3.3 0.00138104 0 0.0013809599999999999 0 0.00138106 3.3 0.00138098 3.3 0.00138108 0 0.0013809999999999998 0 0.0013811 3.3 0.00138102 3.3 0.00138112 0 0.0013810399999999998 0 0.0013811399999999999 3.3 0.00138106 3.3 0.00138116 0 0.0013810799999999998 0 0.0013811799999999999 3.3 0.0013811 3.3 0.0013812 0 0.00138112 0 0.00138122 3.3 0.0013811399999999999 3.3 0.00138124 0 0.00138116 0 0.00138126 3.3 0.0013811799999999999 3.3 0.00138128 0 0.0013812 0 0.0013813 3.3 0.0013812199999999998 3.3 0.00138132 0 0.00138124 0 0.00138134 3.3 0.0013812599999999998 3.3 0.0013813599999999999 0 0.00138128 0 0.00138138 3.3 0.0013813 3.3 0.0013814 0 0.00138132 0 0.00138142 3.3 0.00138134 3.3 0.00138144 0 0.0013813599999999999 0 0.00138146 3.3 0.00138138 3.3 0.00138148 0 0.0013813999999999999 0 0.0013815 3.3 0.00138142 3.3 0.00138152 0 0.0013814399999999998 0 0.00138154 3.3 0.00138146 3.3 0.00138156 0 0.0013814799999999998 0 0.0013815799999999999 3.3 0.0013815 3.3 0.0013816 0 0.00138152 0 0.00138162 3.3 0.00138154 3.3 0.00138164 0 0.00138156 0 0.00138166 3.3 0.0013815799999999999 3.3 0.00138168 0 0.0013816 0 0.0013817 3.3 0.0013816199999999999 3.3 0.00138172 0 0.00138164 0 0.00138174 3.3 0.0013816599999999998 3.3 0.0013817599999999999 0 0.00138168 0 0.00138178 3.3 0.0013816999999999998 3.3 0.0013817999999999999 0 0.00138172 0 0.00138182 3.3 0.00138174 3.3 0.00138184 0 0.0013817599999999999 0 0.00138186 3.3 0.00138178 3.3 0.00138188 0 0.0013817999999999999 0 0.0013819 3.3 0.00138182 3.3 0.00138192 0 0.0013818399999999998 0 0.00138194 3.3 0.00138186 3.3 0.00138196 0 0.0013818799999999998 0 0.0013819799999999999 3.3 0.0013819 3.3 0.001382 0 0.00138192 0 0.00138202 3.3 0.00138194 3.3 0.00138204 0 0.00138196 0 0.00138206 3.3 0.0013819799999999999 3.3 0.00138208 0 0.001382 0 0.0013821 3.3 0.0013820199999999999 3.3 0.00138212 0 0.00138204 0 0.00138214 3.3 0.0013820599999999998 3.3 0.00138216 0 0.00138208 0 0.00138218 3.3 0.0013820999999999998 3.3 0.0013821999999999999 0 0.00138212 0 0.00138222 3.3 0.00138214 3.3 0.00138224 0 0.00138216 0 0.00138226 3.3 0.00138218 3.3 0.00138228 0 0.0013821999999999999 0 0.0013823 3.3 0.00138222 3.3 0.00138232 0 0.0013822399999999999 0 0.00138234 3.3 0.00138226 3.3 0.00138236 0 0.0013822799999999998 0 0.00138238 3.3 0.0013823 3.3 0.0013824 0 0.0013823199999999998 0 0.0013824199999999999 3.3 0.00138234 3.3 0.00138244 0 0.00138236 0 0.00138246 3.3 0.00138238 3.3 0.00138248 0 0.0013824 0 0.0013825 3.3 0.0013824199999999999 3.3 0.00138252 0 0.00138244 0 0.00138254 3.3 0.0013824599999999999 3.3 0.00138256 0 0.00138248 0 0.00138258 3.3 0.0013824999999999998 3.3 0.0013825999999999999 0 0.00138252 0 0.00138262 3.3 0.0013825399999999998 3.3 0.0013826399999999999 0 0.00138256 0 0.00138266 3.3 0.00138258 3.3 0.00138268 0 0.0013825999999999999 0 0.0013827 3.3 0.00138262 3.3 0.00138272 0 0.0013826399999999999 0 0.00138274 3.3 0.00138266 3.3 0.00138276 0 0.0013826799999999998 0 0.00138278 3.3 0.0013827 3.3 0.0013828 0 0.0013827199999999998 0 0.0013828199999999999 3.3 0.00138274 3.3 0.00138284 0 0.00138276 0 0.00138286 3.3 0.00138278 3.3 0.00138288 0 0.0013828 0 0.0013829 3.3 0.0013828199999999999 3.3 0.00138292 0 0.00138284 0 0.00138294 3.3 0.0013828599999999999 3.3 0.00138296 0 0.00138288 0 0.00138298 3.3 0.0013828999999999998 3.3 0.001383 0 0.00138292 0 0.00138302 3.3 0.0013829399999999998 3.3 0.0013830399999999999 0 0.00138296 0 0.00138306 3.3 0.00138298 3.3 0.00138308 0 0.001383 0 0.0013831 3.3 0.00138302 3.3 0.00138312 0 0.0013830399999999999 0 0.00138314 3.3 0.00138306 3.3 0.00138316 0 0.0013830799999999999 0 0.00138318 3.3 0.0013831 3.3 0.0013832 0 0.0013831199999999998 0 0.00138322 3.3 0.00138314 3.3 0.00138324 0 0.0013831599999999998 0 0.0013832599999999999 3.3 0.00138318 3.3 0.00138328 0 0.0013832 0 0.0013833 3.3 0.00138322 3.3 0.00138332 0 0.00138324 0 0.00138334 3.3 0.0013832599999999999 3.3 0.00138336 0 0.00138328 0 0.00138338 3.3 0.0013832999999999999 3.3 0.0013834 0 0.00138332 0 0.00138342 3.3 0.0013833399999999998 3.3 0.0013834399999999999 0 0.00138336 0 0.00138346 3.3 0.0013833799999999998 3.3 0.0013834799999999999 0 0.0013834 0 0.0013835 3.3 0.00138342 3.3 0.00138352 0 0.0013834399999999999 0 0.00138354 3.3 0.00138346 3.3 0.00138356 0 0.0013834799999999999 0 0.00138358 3.3 0.0013835 3.3 0.0013836 0 0.0013835199999999998 0 0.00138362 3.3 0.00138354 3.3 0.00138364 0 0.0013835599999999998 0 0.0013836599999999999 3.3 0.00138358 3.3 0.00138368 0 0.0013836 0 0.0013837 3.3 0.00138362 3.3 0.00138372 0 0.00138364 0 0.00138374 3.3 0.0013836599999999999 3.3 0.00138376 0 0.00138368 0 0.00138378 3.3 0.0013836999999999999 3.3 0.0013838 0 0.00138372 0 0.00138382 3.3 0.0013837399999999998 3.3 0.00138384 0 0.00138376 0 0.00138386 3.3 0.0013837799999999998 3.3 0.0013838799999999999 0 0.0013838 0 0.0013839 3.3 0.00138382 3.3 0.00138392 0 0.00138384 0 0.00138394 3.3 0.00138386 3.3 0.00138396 0 0.0013838799999999999 0 0.00138398 3.3 0.0013839 3.3 0.001384 0 0.0013839199999999999 0 0.00138402 3.3 0.00138394 3.3 0.00138404 0 0.0013839599999999998 0 0.0013840599999999999 3.3 0.00138398 3.3 0.00138408 0 0.0013839999999999998 0 0.0013840999999999999 3.3 0.00138402 3.3 0.00138412 0 0.00138404 0 0.00138414 3.3 0.0013840599999999999 3.3 0.00138416 0 0.00138408 0 0.00138418 3.3 0.0013840999999999999 3.3 0.0013842 0 0.00138412 0 0.00138422 3.3 0.0013841399999999998 3.3 0.00138424 0 0.00138416 0 0.00138426 3.3 0.0013841799999999998 3.3 0.0013842799999999999 0 0.0013842 0 0.0013843 3.3 0.0013842199999999998 3.3 0.0013843199999999999 0 0.00138424 0 0.00138434 3.3 0.00138426 3.3 0.00138436 0 0.0013842799999999999 0 0.00138438 3.3 0.0013843 3.3 0.0013844 0 0.0013843199999999999 0 0.00138442 3.3 0.00138434 3.3 0.00138444 0 0.0013843599999999998 0 0.00138446 3.3 0.00138438 3.3 0.00138448 0 0.0013843999999999998 0 0.0013844999999999999 3.3 0.00138442 3.3 0.00138452 0 0.00138444 0 0.00138454 3.3 0.00138446 3.3 0.00138456 0 0.00138448 0 0.00138458 3.3 0.0013844999999999999 3.3 0.0013846 0 0.00138452 0 0.00138462 3.3 0.0013845399999999999 3.3 0.00138464 0 0.00138456 0 0.00138466 3.3 0.0013845799999999998 3.3 0.00138468 0 0.0013846 0 0.0013847 3.3 0.0013846199999999998 3.3 0.0013847199999999999 0 0.00138464 0 0.00138474 3.3 0.00138466 3.3 0.00138476 0 0.00138468 0 0.00138478 3.3 0.0013847 3.3 0.0013848 0 0.0013847199999999999 0 0.00138482 3.3 0.00138474 3.3 0.00138484 0 0.0013847599999999999 0 0.00138486 3.3 0.00138478 3.3 0.00138488 0 0.0013847999999999998 0 0.0013848999999999999 3.3 0.00138482 3.3 0.00138492 0 0.0013848399999999998 0 0.0013849399999999999 3.3 0.00138486 3.3 0.00138496 0 0.00138488 0 0.00138498 3.3 0.0013848999999999999 3.3 0.001385 0 0.00138492 0 0.00138502 3.3 0.0013849399999999999 3.3 0.00138504 0 0.00138496 0 0.00138506 3.3 0.0013849799999999998 3.3 0.00138508 0 0.001385 0 0.0013851 3.3 0.0013850199999999998 3.3 0.0013851199999999999 0 0.00138504 0 0.00138514 3.3 0.00138506 3.3 0.00138516 0 0.00138508 0 0.00138518 3.3 0.0013851 3.3 0.0013852 0 0.0013851199999999999 0 0.00138522 3.3 0.00138514 3.3 0.00138524 0 0.0013851599999999999 0 0.00138526 3.3 0.00138518 3.3 0.00138528 0 0.0013851999999999998 0 0.0013853 3.3 0.00138522 3.3 0.00138532 0 0.0013852399999999998 0 0.0013853399999999999 3.3 0.00138526 3.3 0.00138536 0 0.00138528 0 0.00138538 3.3 0.0013853 3.3 0.0013854 0 0.00138532 0 0.00138542 3.3 0.0013853399999999999 3.3 0.00138544 0 0.00138536 0 0.00138546 3.3 0.0013853799999999999 3.3 0.00138548 0 0.0013854 0 0.0013855 3.3 0.0013854199999999998 3.3 0.00138552 0 0.00138544 0 0.00138554 3.3 0.0013854599999999998 3.3 0.0013855599999999999 0 0.00138548 0 0.00138558 3.3 0.0013855 3.3 0.0013856 0 0.00138552 0 0.00138562 3.3 0.00138554 3.3 0.00138564 0 0.0013855599999999999 0 0.00138566 3.3 0.00138558 3.3 0.00138568 0 0.0013855999999999999 0 0.0013857 3.3 0.00138562 3.3 0.00138572 0 0.0013856399999999998 0 0.0013857399999999999 3.3 0.00138566 3.3 0.00138576 0 0.0013856799999999998 0 0.0013857799999999999 3.3 0.0013857 3.3 0.0013858 0 0.00138572 0 0.00138582 3.3 0.0013857399999999999 3.3 0.00138584 0 0.00138576 0 0.00138586 3.3 0.0013857799999999999 3.3 0.00138588 0 0.0013858 0 0.0013859 3.3 0.0013858199999999998 3.3 0.00138592 0 0.00138584 0 0.00138594 3.3 0.0013858599999999998 3.3 0.0013859599999999999 0 0.00138588 0 0.00138598 3.3 0.0013859 3.3 0.001386 0 0.00138592 0 0.00138602 3.3 0.00138594 3.3 0.00138604 0 0.0013859599999999999 0 0.00138606 3.3 0.00138598 3.3 0.00138608 0 0.0013859999999999999 0 0.0013861 3.3 0.00138602 3.3 0.00138612 0 0.0013860399999999998 0 0.00138614 3.3 0.00138606 3.3 0.00138616 0 0.0013860799999999998 0 0.0013861799999999999 3.3 0.0013861 3.3 0.0013862 0 0.00138612 0 0.00138622 3.3 0.00138614 3.3 0.00138624 0 0.00138616 0 0.00138626 3.3 0.0013861799999999999 3.3 0.00138628 0 0.0013862 0 0.0013863 3.3 0.0013862199999999999 3.3 0.00138632 0 0.00138624 0 0.00138634 3.3 0.0013862599999999998 3.3 0.00138636 0 0.00138628 0 0.00138638 3.3 0.0013862999999999998 3.3 0.0013863999999999999 0 0.00138632 0 0.00138642 3.3 0.00138634 3.3 0.00138644 0 0.00138636 0 0.00138646 3.3 0.00138638 3.3 0.00138648 0 0.0013863999999999999 0 0.0013865 3.3 0.00138642 3.3 0.00138652 0 0.0013864399999999999 0 0.00138654 3.3 0.00138646 3.3 0.00138656 0 0.0013864799999999998 0 0.0013865799999999999 3.3 0.0013865 3.3 0.0013866 0 0.0013865199999999998 0 0.0013866199999999999 3.3 0.00138654 3.3 0.00138664 0 0.00138656 0 0.00138666 3.3 0.0013865799999999999 3.3 0.00138668 0 0.0013866 0 0.0013867 3.3 0.0013866199999999999 3.3 0.00138672 0 0.00138664 0 0.00138674 3.3 0.0013866599999999998 3.3 0.00138676 0 0.00138668 0 0.00138678 3.3 0.0013866999999999998 3.3 0.0013867999999999999 0 0.00138672 0 0.00138682 3.3 0.00138674 3.3 0.00138684 0 0.00138676 0 0.00138686 3.3 0.00138678 3.3 0.00138688 0 0.0013867999999999999 0 0.0013869 3.3 0.00138682 3.3 0.00138692 0 0.0013868399999999999 0 0.00138694 3.3 0.00138686 3.3 0.00138696 0 0.0013868799999999998 0 0.00138698 3.3 0.0013869 3.3 0.001387 0 0.0013869199999999998 0 0.0013870199999999999 3.3 0.00138694 3.3 0.00138704 0 0.00138696 0 0.00138706 3.3 0.00138698 3.3 0.00138708 0 0.001387 0 0.0013871 3.3 0.0013870199999999999 3.3 0.00138712 0 0.00138704 0 0.00138714 3.3 0.0013870599999999999 3.3 0.00138716 0 0.00138708 0 0.00138718 3.3 0.0013870999999999998 3.3 0.0013871999999999999 0 0.00138712 0 0.00138722 3.3 0.0013871399999999998 3.3 0.0013872399999999999 0 0.00138716 0 0.00138726 3.3 0.00138718 3.3 0.00138728 0 0.0013871999999999999 0 0.0013873 3.3 0.00138722 3.3 0.00138732 0 0.0013872399999999999 0 0.00138734 3.3 0.00138726 3.3 0.00138736 0 0.0013872799999999999 0 0.00138738 3.3 0.0013873 3.3 0.0013874 0 0.0013873199999999998 0 0.0013874199999999999 3.3 0.00138734 3.3 0.00138744 0 0.0013873599999999998 0 0.0013874599999999999 3.3 0.00138738 3.3 0.00138748 0 0.0013874 0 0.0013875 3.3 0.0013874199999999999 3.3 0.00138752 0 0.00138744 0 0.00138754 3.3 0.0013874599999999999 3.3 0.00138756 0 0.00138748 0 0.00138758 3.3 0.0013874999999999998 3.3 0.0013876 0 0.00138752 0 0.00138762 3.3 0.0013875399999999998 3.3 0.0013876399999999999 0 0.00138756 0 0.00138766 3.3 0.00138758 3.3 0.00138768 0 0.0013876 0 0.0013877 3.3 0.00138762 3.3 0.00138772 0 0.0013876399999999999 0 0.00138774 3.3 0.00138766 3.3 0.00138776 0 0.0013876799999999999 0 0.00138778 3.3 0.0013877 3.3 0.0013878 0 0.0013877199999999998 0 0.00138782 3.3 0.00138774 3.3 0.00138784 0 0.0013877599999999998 0 0.0013878599999999999 3.3 0.00138778 3.3 0.00138788 0 0.0013878 0 0.0013879 3.3 0.00138782 3.3 0.00138792 0 0.00138784 0 0.00138794 3.3 0.0013878599999999999 3.3 0.00138796 0 0.00138788 0 0.00138798 3.3 0.0013878999999999999 3.3 0.001388 0 0.00138792 0 0.00138802 3.3 0.0013879399999999998 3.3 0.0013880399999999999 0 0.00138796 0 0.00138806 3.3 0.0013879799999999998 3.3 0.0013880799999999999 0 0.001388 0 0.0013881 3.3 0.00138802 3.3 0.00138812 0 0.0013880399999999999 0 0.00138814 3.3 0.00138806 3.3 0.00138816 0 0.0013880799999999999 0 0.00138818 3.3 0.0013881 3.3 0.0013882 0 0.0013881199999999998 0 0.00138822 3.3 0.00138814 3.3 0.00138824 0 0.0013881599999999998 0 0.0013882599999999999 3.3 0.00138818 3.3 0.00138828 0 0.0013881999999999998 0 0.0013882999999999999 3.3 0.00138822 3.3 0.00138832 0 0.00138824 0 0.00138834 3.3 0.0013882599999999999 3.3 0.00138836 0 0.00138828 0 0.00138838 3.3 0.0013882999999999999 3.3 0.0013884 0 0.00138832 0 0.00138842 3.3 0.0013883399999999998 3.3 0.00138844 0 0.00138836 0 0.00138846 3.3 0.0013883799999999998 3.3 0.0013884799999999999 0 0.0013884 0 0.0013885 3.3 0.00138842 3.3 0.00138852 0 0.00138844 0 0.00138854 3.3 0.00138846 3.3 0.00138856 0 0.0013884799999999999 0 0.00138858 3.3 0.0013885 3.3 0.0013886 0 0.0013885199999999999 0 0.00138862 3.3 0.00138854 3.3 0.00138864 0 0.0013885599999999998 0 0.00138866 3.3 0.00138858 3.3 0.00138868 0 0.0013885999999999998 0 0.0013886999999999999 3.3 0.00138862 3.3 0.00138872 0 0.00138864 0 0.00138874 3.3 0.00138866 3.3 0.00138876 0 0.00138868 0 0.00138878 3.3 0.0013886999999999999 3.3 0.0013888 0 0.00138872 0 0.00138882 3.3 0.0013887399999999999 3.3 0.00138884 0 0.00138876 0 0.00138886 3.3 0.0013887799999999998 3.3 0.0013888799999999999 0 0.0013888 0 0.0013889 3.3 0.0013888199999999998 3.3 0.0013889199999999999 0 0.00138884 0 0.00138894 3.3 0.00138886 3.3 0.00138896 0 0.0013888799999999999 0 0.00138898 3.3 0.0013889 3.3 0.001389 0 0.0013889199999999999 0 0.00138902 3.3 0.00138894 3.3 0.00138904 0 0.0013889599999999998 0 0.00138906 3.3 0.00138898 3.3 0.00138908 0 0.0013889999999999998 0 0.0013890999999999999 3.3 0.00138902 3.3 0.00138912 0 0.00138904 0 0.00138914 3.3 0.00138906 3.3 0.00138916 0 0.00138908 0 0.00138918 3.3 0.0013890999999999999 3.3 0.0013892 0 0.00138912 0 0.00138922 3.3 0.0013891399999999999 3.3 0.00138924 0 0.00138916 0 0.00138926 3.3 0.0013891799999999998 3.3 0.00138928 0 0.0013892 0 0.0013893 3.3 0.0013892199999999998 3.3 0.0013893199999999999 0 0.00138924 0 0.00138934 3.3 0.00138926 3.3 0.00138936 0 0.00138928 0 0.00138938 3.3 0.0013893 3.3 0.0013894 0 0.0013893199999999999 0 0.00138942 3.3 0.00138934 3.3 0.00138944 0 0.0013893599999999999 0 0.00138946 3.3 0.00138938 3.3 0.00138948 0 0.0013893999999999998 0 0.0013895 3.3 0.00138942 3.3 0.00138952 0 0.0013894399999999998 0 0.0013895399999999999 3.3 0.00138946 3.3 0.00138956 0 0.00138948 0 0.00138958 3.3 0.0013895 3.3 0.0013896 0 0.00138952 0 0.00138962 3.3 0.0013895399999999999 3.3 0.00138964 0 0.00138956 0 0.00138966 3.3 0.0013895799999999999 3.3 0.00138968 0 0.0013896 0 0.0013897 3.3 0.0013896199999999998 3.3 0.0013897199999999999 0 0.00138964 0 0.00138974 3.3 0.0013896599999999998 3.3 0.0013897599999999999 0 0.00138968 0 0.00138978 3.3 0.0013897 3.3 0.0013898 0 0.0013897199999999999 0 0.00138982 3.3 0.00138974 3.3 0.00138984 0 0.0013897599999999999 0 0.00138986 3.3 0.00138978 3.3 0.00138988 0 0.0013897999999999998 0 0.0013899 3.3 0.00138982 3.3 0.00138992 0 0.0013898399999999998 0 0.0013899399999999999 3.3 0.00138986 3.3 0.00138996 0 0.00138988 0 0.00138998 3.3 0.0013899 3.3 0.00139 0 0.00138992 0 0.00139002 3.3 0.0013899399999999999 3.3 0.00139004 0 0.00138996 0 0.00139006 3.3 0.0013899799999999999 3.3 0.00139008 0 0.00139 0 0.0013901 3.3 0.0013900199999999998 3.3 0.00139012 0 0.00139004 0 0.00139014 3.3 0.0013900599999999998 3.3 0.0013901599999999999 0 0.00139008 0 0.00139018 3.3 0.0013901 3.3 0.0013902 0 0.00139012 0 0.00139022 3.3 0.00139014 3.3 0.00139024 0 0.0013901599999999999 0 0.00139026 3.3 0.00139018 3.3 0.00139028 0 0.0013901999999999999 0 0.0013903 3.3 0.00139022 3.3 0.00139032 0 0.0013902399999999998 0 0.00139034 3.3 0.00139026 3.3 0.00139036 0 0.0013902799999999998 0 0.0013903799999999999 3.3 0.0013903 3.3 0.0013904 0 0.00139032 0 0.00139042 3.3 0.00139034 3.3 0.00139044 0 0.00139036 0 0.00139046 3.3 0.0013903799999999999 3.3 0.00139048 0 0.0013904 0 0.0013905 3.3 0.0013904199999999999 3.3 0.00139052 0 0.00139044 0 0.00139054 3.3 0.0013904599999999998 3.3 0.0013905599999999999 0 0.00139048 0 0.00139058 3.3 0.0013904999999999998 3.3 0.0013905999999999999 0 0.00139052 0 0.00139062 3.3 0.00139054 3.3 0.00139064 0 0.0013905599999999999 0 0.00139066 3.3 0.00139058 3.3 0.00139068 0 0.0013905999999999999 0 0.0013907 3.3 0.00139062 3.3 0.00139072 0 0.0013906399999999998 0 0.00139074 3.3 0.00139066 3.3 0.00139076 0 0.0013906799999999998 0 0.0013907799999999999 3.3 0.0013907 3.3 0.0013908 0 0.00139072 0 0.00139082 3.3 0.00139074 3.3 0.00139084 0 0.00139076 0 0.00139086 3.3 0.0013907799999999999 3.3 0.00139088 0 0.0013908 0 0.0013909 3.3 0.0013908199999999999 3.3 0.00139092 0 0.00139084 0 0.00139094 3.3 0.0013908599999999998 3.3 0.00139096 0 0.00139088 0 0.00139098 3.3 0.0013908999999999998 3.3 0.0013909999999999999 0 0.00139092 0 0.00139102 3.3 0.00139094 3.3 0.00139104 0 0.00139096 0 0.00139106 3.3 0.00139098 3.3 0.00139108 0 0.0013909999999999999 0 0.0013911 3.3 0.00139102 3.3 0.00139112 0 0.0013910399999999999 0 0.00139114 3.3 0.00139106 3.3 0.00139116 0 0.0013910799999999998 0 0.0013911799999999999 3.3 0.0013911 3.3 0.0013912 0 0.0013911199999999998 0 0.0013912199999999999 3.3 0.00139114 3.3 0.00139124 0 0.00139116 0 0.00139126 3.3 0.0013911799999999999 3.3 0.00139128 0 0.0013912 0 0.0013913 3.3 0.0013912199999999999 3.3 0.00139132 0 0.00139124 0 0.00139134 3.3 0.0013912599999999998 3.3 0.00139136 0 0.00139128 0 0.00139138 3.3 0.0013912999999999998 3.3 0.0013913999999999999 0 0.00139132 0 0.00139142 3.3 0.0013913399999999998 3.3 0.0013914399999999999 0 0.00139136 0 0.00139146 3.3 0.00139138 3.3 0.00139148 0 0.0013913999999999999 0 0.0013915 3.3 0.00139142 3.3 0.00139152 0 0.0013914399999999999 0 0.00139154 3.3 0.00139146 3.3 0.00139156 0 0.0013914799999999998 0 0.00139158 3.3 0.0013915 3.3 0.0013916 0 0.0013915199999999998 0 0.0013916199999999999 3.3 0.00139154 3.3 0.00139164 0 0.00139156 0 0.00139166 3.3 0.00139158 3.3 0.00139168 0 0.0013916 0 0.0013917 3.3 0.0013916199999999999 3.3 0.00139172 0 0.00139164 0 0.00139174 3.3 0.0013916599999999999 3.3 0.00139176 0 0.00139168 0 0.00139178 3.3 0.0013916999999999998 3.3 0.0013918 0 0.00139172 0 0.00139182 3.3 0.0013917399999999998 3.3 0.0013918399999999999 0 0.00139176 0 0.00139186 3.3 0.00139178 3.3 0.00139188 0 0.0013918 0 0.0013919 3.3 0.00139182 3.3 0.00139192 0 0.0013918399999999999 0 0.00139194 3.3 0.00139186 3.3 0.00139196 0 0.0013918799999999999 0 0.00139198 3.3 0.0013919 3.3 0.001392 0 0.0013919199999999998 0 0.0013920199999999999 3.3 0.00139194 3.3 0.00139204 0 0.0013919599999999998 0 0.0013920599999999999 3.3 0.00139198 3.3 0.00139208 0 0.001392 0 0.0013921 3.3 0.0013920199999999999 3.3 0.00139212 0 0.00139204 0 0.00139214 3.3 0.0013920599999999999 3.3 0.00139216 0 0.00139208 0 0.00139218 3.3 0.0013920999999999998 3.3 0.0013922 0 0.00139212 0 0.00139222 3.3 0.0013921399999999998 3.3 0.0013922399999999999 0 0.00139216 0 0.00139226 3.3 0.00139218 3.3 0.00139228 0 0.0013922 0 0.0013923 3.3 0.00139222 3.3 0.00139232 0 0.0013922399999999999 0 0.00139234 3.3 0.00139226 3.3 0.00139236 0 0.0013922799999999999 0 0.00139238 3.3 0.0013923 3.3 0.0013924 0 0.0013923199999999998 0 0.00139242 3.3 0.00139234 3.3 0.00139244 0 0.0013923599999999998 0 0.0013924599999999999 3.3 0.00139238 3.3 0.00139248 0 0.0013924 0 0.0013925 3.3 0.00139242 3.3 0.00139252 0 0.00139244 0 0.00139254 3.3 0.0013924599999999999 3.3 0.00139256 0 0.00139248 0 0.00139258 3.3 0.0013924999999999999 3.3 0.0013926 0 0.00139252 0 0.00139262 3.3 0.0013925399999999998 3.3 0.00139264 0 0.00139256 0 0.00139266 3.3 0.0013925799999999998 3.3 0.0013926799999999999 0 0.0013926 0 0.0013927 3.3 0.00139262 3.3 0.00139272 0 0.00139264 0 0.00139274 3.3 0.00139266 3.3 0.00139276 0 0.0013926799999999999 0 0.00139278 3.3 0.0013927 3.3 0.0013928 0 0.0013927199999999999 0 0.00139282 3.3 0.00139274 3.3 0.00139284 0 0.0013927599999999998 0 0.0013928599999999999 3.3 0.00139278 3.3 0.00139288 0 0.0013927999999999998 0 0.0013928999999999999 3.3 0.00139282 3.3 0.00139292 0 0.00139284 0 0.00139294 3.3 0.0013928599999999999 3.3 0.00139296 0 0.00139288 0 0.00139298 3.3 0.0013928999999999999 3.3 0.001393 0 0.00139292 0 0.00139302 3.3 0.0013929399999999998 3.3 0.00139304 0 0.00139296 0 0.00139306 3.3 0.0013929799999999998 3.3 0.0013930799999999999 0 0.001393 0 0.0013931 3.3 0.00139302 3.3 0.00139312 0 0.00139304 0 0.00139314 3.3 0.00139306 3.3 0.00139316 0 0.0013930799999999999 0 0.00139318 3.3 0.0013931 3.3 0.0013932 0 0.0013931199999999999 0 0.00139322 3.3 0.00139314 3.3 0.00139324 0 0.0013931599999999998 0 0.00139326 3.3 0.00139318 3.3 0.00139328 0 0.0013931999999999998 0 0.0013932999999999999 3.3 0.00139322 3.3 0.00139332 0 0.00139324 0 0.00139334 3.3 0.00139326 3.3 0.00139336 0 0.00139328 0 0.00139338 3.3 0.0013932999999999999 3.3 0.0013934 0 0.00139332 0 0.00139342 3.3 0.0013933399999999999 3.3 0.00139344 0 0.00139336 0 0.00139346 3.3 0.0013933799999999998 3.3 0.00139348 0 0.0013934 0 0.0013935 3.3 0.0013934199999999998 3.3 0.0013935199999999999 0 0.00139344 0 0.00139354 3.3 0.00139346 3.3 0.00139356 0 0.00139348 0 0.00139358 3.3 0.0013935 3.3 0.0013936 0 0.0013935199999999999 0 0.00139362 3.3 0.00139354 3.3 0.00139364 0 0.0013935599999999999 0 0.00139366 3.3 0.00139358 3.3 0.00139368 0 0.0013935999999999998 0 0.0013936999999999999 3.3 0.00139362 3.3 0.00139372 0 0.0013936399999999998 0 0.0013937399999999999 3.3 0.00139366 3.3 0.00139376 0 0.00139368 0 0.00139378 3.3 0.0013936999999999999 3.3 0.0013938 0 0.00139372 0 0.00139382 3.3 0.0013937399999999999 3.3 0.00139384 0 0.00139376 0 0.00139386 3.3 0.0013937799999999998 3.3 0.00139388 0 0.0013938 0 0.0013939 3.3 0.0013938199999999998 3.3 0.0013939199999999999 0 0.00139384 0 0.00139394 3.3 0.00139386 3.3 0.00139396 0 0.00139388 0 0.00139398 3.3 0.0013939 3.3 0.001394 0 0.0013939199999999999 0 0.00139402 3.3 0.00139394 3.3 0.00139404 0 0.0013939599999999999 0 0.00139406 3.3 0.00139398 3.3 0.00139408 0 0.0013939999999999998 0 0.0013941 3.3 0.00139402 3.3 0.00139412 0 0.0013940399999999998 0 0.0013941399999999999 3.3 0.00139406 3.3 0.00139416 0 0.00139408 0 0.00139418 3.3 0.0013941 3.3 0.0013942 0 0.00139412 0 0.00139422 3.3 0.0013941399999999999 3.3 0.00139424 0 0.00139416 0 0.00139426 3.3 0.0013941799999999999 3.3 0.00139428 0 0.0013942 0 0.0013943 3.3 0.0013942199999999998 3.3 0.0013943199999999999 0 0.00139424 0 0.00139434 3.3 0.0013942599999999998 3.3 0.0013943599999999999 0 0.00139428 0 0.00139438 3.3 0.0013943 3.3 0.0013944 0 0.0013943199999999999 0 0.00139442 3.3 0.00139434 3.3 0.00139444 0 0.0013943599999999999 0 0.00139446 3.3 0.00139438 3.3 0.00139448 0 0.0013943999999999998 0 0.0013945 3.3 0.00139442 3.3 0.00139452 0 0.0013944399999999998 0 0.0013945399999999999 3.3 0.00139446 3.3 0.00139456 0 0.0013944799999999998 0 0.0013945799999999999 3.3 0.0013945 3.3 0.0013946 0 0.00139452 0 0.00139462 3.3 0.0013945399999999999 3.3 0.00139464 0 0.00139456 0 0.00139466 3.3 0.0013945799999999999 3.3 0.00139468 0 0.0013946 0 0.0013947 3.3 0.0013946199999999998 3.3 0.00139472 0 0.00139464 0 0.00139474 3.3 0.0013946599999999998 3.3 0.0013947599999999999 0 0.00139468 0 0.00139478 3.3 0.0013947 3.3 0.0013948 0 0.00139472 0 0.00139482 3.3 0.00139474 3.3 0.00139484 0 0.0013947599999999999 0 0.00139486 3.3 0.00139478 3.3 0.00139488 0 0.0013947999999999999 0 0.0013949 3.3 0.00139482 3.3 0.00139492 0 0.0013948399999999998 0 0.00139494 3.3 0.00139486 3.3 0.00139496 0 0.0013948799999999998 0 0.0013949799999999999 3.3 0.0013949 3.3 0.001395 0 0.00139492 0 0.00139502 3.3 0.00139494 3.3 0.00139504 0 0.00139496 0 0.00139506 3.3 0.0013949799999999999 3.3 0.00139508 0 0.001395 0 0.0013951 3.3 0.0013950199999999999 3.3 0.00139512 0 0.00139504 0 0.00139514 3.3 0.0013950599999999998 3.3 0.0013951599999999999 0 0.00139508 0 0.00139518 3.3 0.0013950999999999998 3.3 0.0013951999999999999 0 0.00139512 0 0.00139522 3.3 0.00139514 3.3 0.00139524 0 0.0013951599999999999 0 0.00139526 3.3 0.00139518 3.3 0.00139528 0 0.0013951999999999999 0 0.0013953 3.3 0.00139522 3.3 0.00139532 0 0.0013952399999999998 0 0.00139534 3.3 0.00139526 3.3 0.00139536 0 0.0013952799999999998 0 0.0013953799999999999 3.3 0.0013953 3.3 0.0013954 0 0.0013953199999999998 0 0.0013954199999999999 3.3 0.00139534 3.3 0.00139544 0 0.00139536 0 0.00139546 3.3 0.0013953799999999999 3.3 0.00139548 0 0.0013954 0 0.0013955 3.3 0.0013954199999999999 3.3 0.00139552 0 0.00139544 0 0.00139554 3.3 0.0013954599999999998 3.3 0.00139556 0 0.00139548 0 0.00139558 3.3 0.0013954999999999998 3.3 0.0013955999999999999 0 0.00139552 0 0.00139562 3.3 0.00139554 3.3 0.00139564 0 0.00139556 0 0.00139566 3.3 0.00139558 3.3 0.00139568 0 0.0013955999999999999 0 0.0013957 3.3 0.00139562 3.3 0.00139572 0 0.0013956399999999999 0 0.00139574 3.3 0.00139566 3.3 0.00139576 0 0.0013956799999999998 0 0.00139578 3.3 0.0013957 3.3 0.0013958 0 0.0013957199999999998 0 0.0013958199999999999 3.3 0.00139574 3.3 0.00139584 0 0.00139576 0 0.00139586 3.3 0.00139578 3.3 0.00139588 0 0.0013958 0 0.0013959 3.3 0.0013958199999999999 3.3 0.00139592 0 0.00139584 0 0.00139594 3.3 0.0013958599999999999 3.3 0.00139596 0 0.00139588 0 0.00139598 3.3 0.0013958999999999998 3.3 0.0013959999999999999 0 0.00139592 0 0.00139602 3.3 0.0013959399999999998 3.3 0.0013960399999999999 0 0.00139596 0 0.00139606 3.3 0.00139598 3.3 0.00139608 0 0.0013959999999999999 0 0.0013961 3.3 0.00139602 3.3 0.00139612 0 0.0013960399999999999 0 0.00139614 3.3 0.00139606 3.3 0.00139616 0 0.0013960799999999998 0 0.00139618 3.3 0.0013961 3.3 0.0013962 0 0.0013961199999999998 0 0.0013962199999999999 3.3 0.00139614 3.3 0.00139624 0 0.00139616 0 0.00139626 3.3 0.00139618 3.3 0.00139628 0 0.0013962 0 0.0013963 3.3 0.0013962199999999999 3.3 0.00139632 0 0.00139624 0 0.00139634 3.3 0.0013962599999999999 3.3 0.00139636 0 0.00139628 0 0.00139638 3.3 0.0013962999999999998 3.3 0.0013964 0 0.00139632 0 0.00139642 3.3 0.0013963399999999998 3.3 0.0013964399999999999 0 0.00139636 0 0.00139646 3.3 0.00139638 3.3 0.00139648 0 0.0013964 0 0.0013965 3.3 0.00139642 3.3 0.00139652 0 0.0013964399999999999 0 0.00139654 3.3 0.00139646 3.3 0.00139656 0 0.0013964799999999999 0 0.00139658 3.3 0.0013965 3.3 0.0013966 0 0.0013965199999999998 0 0.00139662 3.3 0.00139654 3.3 0.00139664 0 0.0013965599999999998 0 0.0013966599999999999 3.3 0.00139658 3.3 0.00139668 0 0.0013966 0 0.0013967 3.3 0.00139662 3.3 0.00139672 0 0.00139664 0 0.00139674 3.3 0.0013966599999999999 3.3 0.00139676 0 0.00139668 0 0.00139678 3.3 0.0013966999999999999 3.3 0.0013968 0 0.00139672 0 0.00139682 3.3 0.0013967399999999998 3.3 0.0013968399999999999 0 0.00139676 0 0.00139686 3.3 0.0013967799999999998 3.3 0.0013968799999999999 0 0.0013968 0 0.0013969 3.3 0.00139682 3.3 0.00139692 0 0.0013968399999999999 0 0.00139694 3.3 0.00139686 3.3 0.00139696 0 0.0013968799999999999 0 0.00139698 3.3 0.0013969 3.3 0.001397 0 0.0013969199999999998 0 0.00139702 3.3 0.00139694 3.3 0.00139704 0 0.0013969599999999998 0 0.0013970599999999999 3.3 0.00139698 3.3 0.00139708 0 0.001397 0 0.0013971 3.3 0.00139702 3.3 0.00139712 0 0.00139704 0 0.00139714 3.3 0.0013970599999999999 3.3 0.00139716 0 0.00139708 0 0.00139718 3.3 0.0013970999999999999 3.3 0.0013972 0 0.00139712 0 0.00139722 3.3 0.0013971399999999998 3.3 0.00139724 0 0.00139716 0 0.00139726 3.3 0.0013971799999999998 3.3 0.0013972799999999999 0 0.0013972 0 0.0013973 3.3 0.00139722 3.3 0.00139732 0 0.00139724 0 0.00139734 3.3 0.00139726 3.3 0.00139736 0 0.0013972799999999999 0 0.00139738 3.3 0.0013973 3.3 0.0013974 0 0.0013973199999999999 0 0.00139742 3.3 0.00139734 3.3 0.00139744 0 0.0013973599999999998 0 0.0013974599999999999 3.3 0.00139738 3.3 0.00139748 0 0.0013973999999999998 0 0.0013974999999999999 3.3 0.00139742 3.3 0.00139752 0 0.00139744 0 0.00139754 3.3 0.0013974599999999999 3.3 0.00139756 0 0.00139748 0 0.00139758 3.3 0.0013974999999999999 3.3 0.0013976 0 0.00139752 0 0.00139762 3.3 0.0013975399999999999 3.3 0.00139764 0 0.00139756 0 0.00139766 3.3 0.0013975799999999998 3.3 0.0013976799999999999 0 0.0013976 0 0.0013977 3.3 0.0013976199999999998 3.3 0.0013977199999999999 0 0.00139764 0 0.00139774 3.3 0.00139766 3.3 0.00139776 0 0.0013976799999999999 0 0.00139778 3.3 0.0013977 3.3 0.0013978 0 0.0013977199999999999 0 0.00139782 3.3 0.00139774 3.3 0.00139784 0 0.0013977599999999998 0 0.00139786 3.3 0.00139778 3.3 0.00139788 0 0.0013977999999999998 0 0.0013978999999999999 3.3 0.00139782 3.3 0.00139792 0 0.00139784 0 0.00139794 3.3 0.00139786 3.3 0.00139796 0 0.00139788 0 0.00139798 3.3 0.0013978999999999999 3.3 0.001398 0 0.00139792 0 0.00139802 3.3 0.0013979399999999999 3.3 0.00139804 0 0.00139796 0 0.00139806 3.3 0.0013979799999999998 3.3 0.00139808 0 0.001398 0 0.0013981 3.3 0.0013980199999999998 3.3 0.0013981199999999999 0 0.00139804 0 0.00139814 3.3 0.00139806 3.3 0.00139816 0 0.00139808 0 0.00139818 3.3 0.0013981 3.3 0.0013982 0 0.0013981199999999999 0 0.00139822 3.3 0.00139814 3.3 0.00139824 0 0.0013981599999999999 0 0.00139826 3.3 0.00139818 3.3 0.00139828 0 0.0013981999999999998 0 0.0013982999999999999 3.3 0.00139822 3.3 0.00139832 0 0.0013982399999999998 0 0.0013983399999999999 3.3 0.00139826 3.3 0.00139836 0 0.00139828 0 0.00139838 3.3 0.0013982999999999999 3.3 0.0013984 0 0.00139832 0 0.00139842 3.3 0.0013983399999999999 3.3 0.00139844 0 0.00139836 0 0.00139846 3.3 0.0013983799999999998 3.3 0.00139848 0 0.0013984 0 0.0013985 3.3 0.0013984199999999998 3.3 0.0013985199999999999 0 0.00139844 0 0.00139854 3.3 0.0013984599999999998 3.3 0.0013985599999999999 0 0.00139848 0 0.00139858 3.3 0.0013985 3.3 0.0013986 0 0.0013985199999999999 0 0.00139862 3.3 0.00139854 3.3 0.00139864 0 0.0013985599999999999 0 0.00139866 3.3 0.00139858 3.3 0.00139868 0 0.0013985999999999998 0 0.0013987 3.3 0.00139862 3.3 0.00139872 0 0.0013986399999999998 0 0.0013987399999999999 3.3 0.00139866 3.3 0.00139876 0 0.00139868 0 0.00139878 3.3 0.0013987 3.3 0.0013988 0 0.00139872 0 0.00139882 3.3 0.0013987399999999999 3.3 0.00139884 0 0.00139876 0 0.00139886 3.3 0.0013987799999999999 3.3 0.00139888 0 0.0013988 0 0.0013989 3.3 0.0013988199999999998 3.3 0.00139892 0 0.00139884 0 0.00139894 3.3 0.0013988599999999998 3.3 0.0013989599999999999 0 0.00139888 0 0.00139898 3.3 0.0013989 3.3 0.001399 0 0.00139892 0 0.00139902 3.3 0.00139894 3.3 0.00139904 0 0.0013989599999999999 0 0.00139906 3.3 0.00139898 3.3 0.00139908 0 0.0013989999999999999 0 0.0013991 3.3 0.00139902 3.3 0.00139912 0 0.0013990399999999998 0 0.0013991399999999999 3.3 0.00139906 3.3 0.00139916 0 0.0013990799999999998 0 0.0013991799999999999 3.3 0.0013991 3.3 0.0013992 0 0.00139912 0 0.00139922 3.3 0.0013991399999999999 3.3 0.00139924 0 0.00139916 0 0.00139926 3.3 0.0013991799999999999 3.3 0.00139928 0 0.0013992 0 0.0013993 3.3 0.0013992199999999998 3.3 0.00139932 0 0.00139924 0 0.00139934 3.3 0.0013992599999999998 3.3 0.0013993599999999999 0 0.00139928 0 0.00139938 3.3 0.0013993 3.3 0.0013994 0 0.00139932 0 0.00139942 3.3 0.00139934 3.3 0.00139944 0 0.0013993599999999999 0 0.00139946 3.3 0.00139938 3.3 0.00139948 0 0.0013993999999999999 0 0.0013995 3.3 0.00139942 3.3 0.00139952 0 0.0013994399999999998 0 0.00139954 3.3 0.00139946 3.3 0.00139956 0 0.0013994799999999998 0 0.0013995799999999999 3.3 0.0013995 3.3 0.0013996 0 0.00139952 0 0.00139962 3.3 0.00139954 3.3 0.00139964 0 0.00139956 0 0.00139966 3.3 0.0013995799999999999 3.3 0.00139968 0 0.0013996 0 0.0013997 3.3 0.0013996199999999999 3.3 0.00139972 0 0.00139964 0 0.00139974 3.3 0.0013996599999999998 3.3 0.00139976 0 0.00139968 0 0.00139978 3.3 0.0013996999999999998 3.3 0.0013997999999999999 0 0.00139972 0 0.00139982 3.3 0.00139974 3.3 0.00139984 0 0.00139976 0 0.00139986 3.3 0.00139978 3.3 0.00139988 0 0.0013997999999999999 0 0.0013999 3.3 0.00139982 3.3 0.00139992 0 0.0013998399999999999 0 0.00139994 3.3 0.00139986 3.3 0.00139996 0 0.0013998799999999998 0 0.0013999799999999999 3.3 0.0013999 3.3 0.0014 0 0.0013999199999999998 0 0.0014000199999999999 3.3 0.00139994 3.3 0.00140004 0 0.00139996 0 0.00140006 3.3 0.0013999799999999999 3.3 0.00140008 0 0.0014 0 0.0014001 3.3 0.0014000199999999999 3.3 0.00140012 0 0.00140004 0 0.00140014 3.3 0.0014000599999999998 3.3 0.00140016 0 0.00140008 0 0.00140018 3.3 0.0014000999999999998 3.3 0.0014001999999999999 0 0.00140012 0 0.00140022 3.3 0.00140014 3.3 0.00140024 0 0.00140016 0 0.00140026 3.3 0.00140018 3.3 0.00140028 0 0.0014001999999999999 0 0.0014003 3.3 0.00140022 3.3 0.00140032 0 0.0014002399999999999 0 0.00140034 3.3 0.00140026 3.3 0.00140036 0 0.0014002799999999998 0 0.00140038 3.3 0.0014003 3.3 0.0014004 0 0.0014003199999999998 0 0.0014004199999999999 3.3 0.00140034 3.3 0.00140044 0 0.00140036 0 0.00140046 3.3 0.00140038 3.3 0.00140048 0 0.0014004 0 0.0014005 3.3 0.0014004199999999999 3.3 0.00140052 0 0.00140044 0 0.00140054 3.3 0.0014004599999999999 3.3 0.00140056 0 0.00140048 0 0.00140058 3.3 0.0014004999999999998 3.3 0.0014006 0 0.00140052 0 0.00140062 3.3 0.0014005399999999998 3.3 0.0014006399999999999 0 0.00140056 0 0.00140066 3.3 0.00140058 3.3 0.00140068 0 0.0014006 0 0.0014007 3.3 0.00140062 3.3 0.00140072 0 0.0014006399999999999 0 0.00140074 3.3 0.00140066 3.3 0.00140076 0 0.0014006799999999999 0 0.00140078 3.3 0.0014007 3.3 0.0014008 0 0.0014007199999999998 0 0.0014008199999999999 3.3 0.00140074 3.3 0.00140084 0 0.0014007599999999998 0 0.0014008599999999999 3.3 0.00140078 3.3 0.00140088 0 0.0014008 0 0.0014009 3.3 0.0014008199999999999 3.3 0.00140092 0 0.00140084 0 0.00140094 3.3 0.0014008599999999999 3.3 0.00140096 0 0.00140088 0 0.00140098 3.3 0.0014008999999999998 3.3 0.001401 0 0.00140092 0 0.00140102 3.3 0.0014009399999999998 3.3 0.0014010399999999999 0 0.00140096 0 0.00140106 3.3 0.00140098 3.3 0.00140108 0 0.001401 0 0.0014011 3.3 0.00140102 3.3 0.00140112 0 0.0014010399999999999 0 0.00140114 3.3 0.00140106 3.3 0.00140116 0 0.0014010799999999999 0 0.00140118 3.3 0.0014011 3.3 0.0014012 0 0.0014011199999999998 0 0.00140122 3.3 0.00140114 3.3 0.00140124 0 0.0014011599999999998 0 0.0014012599999999999 3.3 0.00140118 3.3 0.00140128 0 0.0014012 0 0.0014013 3.3 0.00140122 3.3 0.00140132 0 0.00140124 0 0.00140134 3.3 0.0014012599999999999 3.3 0.00140136 0 0.00140128 0 0.00140138 3.3 0.0014012999999999999 3.3 0.0014014 0 0.00140132 0 0.00140142 3.3 0.0014013399999999998 3.3 0.0014014399999999999 0 0.00140136 0 0.00140146 3.3 0.0014013799999999998 3.3 0.0014014799999999999 0 0.0014014 0 0.0014015 3.3 0.00140142 3.3 0.00140152 0 0.0014014399999999999 0 0.00140154 3.3 0.00140146 3.3 0.00140156 0 0.0014014799999999999 0 0.00140158 3.3 0.0014015 3.3 0.0014016 0 0.0014015199999999998 0 0.00140162 3.3 0.00140154 3.3 0.00140164 0 0.0014015599999999998 0 0.0014016599999999999 3.3 0.00140158 3.3 0.00140168 0 0.0014015999999999998 0 0.0014016999999999999 3.3 0.00140162 3.3 0.00140172 0 0.00140164 0 0.00140174 3.3 0.0014016599999999999 3.3 0.00140176 0 0.00140168 0 0.00140178 3.3 0.0014016999999999999 3.3 0.0014018 0 0.00140172 0 0.00140182 3.3 0.0014017399999999998 3.3 0.00140184 0 0.00140176 0 0.00140186 3.3 0.0014017799999999998 3.3 0.0014018799999999999 0 0.0014018 0 0.0014019 3.3 0.00140182 3.3 0.00140192 0 0.00140184 0 0.00140194 3.3 0.00140186 3.3 0.00140196 0 0.0014018799999999999 0 0.00140198 3.3 0.0014019 3.3 0.001402 0 0.0014019199999999999 0 0.00140202 3.3 0.00140194 3.3 0.00140204 0 0.0014019599999999998 0 0.00140206 3.3 0.00140198 3.3 0.00140208 0 0.0014019999999999998 0 0.0014020999999999999 3.3 0.00140202 3.3 0.00140212 0 0.00140204 0 0.00140214 3.3 0.00140206 3.3 0.00140216 0 0.00140208 0 0.00140218 3.3 0.0014020999999999999 3.3 0.0014022 0 0.00140212 0 0.00140222 3.3 0.0014021399999999999 3.3 0.00140224 0 0.00140216 0 0.00140226 3.3 0.0014021799999999998 3.3 0.0014022799999999999 0 0.0014022 0 0.0014023 3.3 0.0014022199999999998 3.3 0.0014023199999999999 0 0.00140224 0 0.00140234 3.3 0.00140226 3.3 0.00140236 0 0.0014022799999999999 0 0.00140238 3.3 0.0014023 3.3 0.0014024 0 0.0014023199999999999 0 0.00140242 3.3 0.00140234 3.3 0.00140244 0 0.0014023599999999998 0 0.00140246 3.3 0.00140238 3.3 0.00140248 0 0.0014023999999999998 0 0.0014024999999999999 3.3 0.00140242 3.3 0.00140252 0 0.00140244 0 0.00140254 3.3 0.00140246 3.3 0.00140256 0 0.00140248 0 0.00140258 3.3 0.0014024999999999999 3.3 0.0014026 0 0.00140252 0 0.00140262 3.3 0.0014025399999999999 3.3 0.00140264 0 0.00140256 0 0.00140266 3.3 0.0014025799999999998 3.3 0.00140268 0 0.0014026 0 0.0014027 3.3 0.0014026199999999998 3.3 0.0014027199999999999 0 0.00140264 0 0.00140274 3.3 0.00140266 3.3 0.00140276 0 0.00140268 0 0.00140278 3.3 0.0014027 3.3 0.0014028 0 0.0014027199999999999 0 0.00140282 3.3 0.00140274 3.3 0.00140284 0 0.0014027599999999999 0 0.00140286 3.3 0.00140278 3.3 0.00140288 0 0.0014027999999999998 0 0.0014029 3.3 0.00140282 3.3 0.00140292 0 0.0014028399999999998 0 0.0014029399999999999 3.3 0.00140286 3.3 0.00140296 0 0.00140288 0 0.00140298 3.3 0.0014029 3.3 0.001403 0 0.00140292 0 0.00140302 3.3 0.0014029399999999999 3.3 0.00140304 0 0.00140296 0 0.00140306 3.3 0.0014029799999999999 3.3 0.00140308 0 0.001403 0 0.0014031 3.3 0.0014030199999999998 3.3 0.0014031199999999999 0 0.00140304 0 0.00140314 3.3 0.0014030599999999998 3.3 0.0014031599999999999 0 0.00140308 0 0.00140318 3.3 0.0014031 3.3 0.0014032 0 0.0014031199999999999 0 0.00140322 3.3 0.00140314 3.3 0.00140324 0 0.0014031599999999999 0 0.00140326 3.3 0.00140318 3.3 0.00140328 0 0.0014031999999999998 0 0.0014033 3.3 0.00140322 3.3 0.00140332 0 0.0014032399999999998 0 0.0014033399999999999 3.3 0.00140326 3.3 0.00140336 0 0.00140328 0 0.00140338 3.3 0.0014033 3.3 0.0014034 0 0.00140332 0 0.00140342 3.3 0.0014033399999999999 3.3 0.00140344 0 0.00140336 0 0.00140346 3.3 0.0014033799999999999 3.3 0.00140348 0 0.0014034 0 0.0014035 3.3 0.0014034199999999998 3.3 0.00140352 0 0.00140344 0 0.00140354 3.3 0.0014034599999999998 3.3 0.0014035599999999999 0 0.00140348 0 0.00140358 3.3 0.0014035 3.3 0.0014036 0 0.00140352 0 0.00140362 3.3 0.00140354 3.3 0.00140364 0 0.0014035599999999999 0 0.00140366 3.3 0.00140358 3.3 0.00140368 0 0.0014035999999999999 0 0.0014037 3.3 0.00140362 3.3 0.00140372 0 0.0014036399999999998 0 0.00140374 3.3 0.00140366 3.3 0.00140376 0 0.0014036799999999998 0 0.0014037799999999999 3.3 0.0014037 3.3 0.0014038 0 0.00140372 0 0.00140382 3.3 0.00140374 3.3 0.00140384 0 0.00140376 0 0.00140386 3.3 0.0014037799999999999 3.3 0.00140388 0 0.0014038 0 0.0014039 3.3 0.0014038199999999999 3.3 0.00140392 0 0.00140384 0 0.00140394 3.3 0.0014038599999999998 3.3 0.0014039599999999999 0 0.00140388 0 0.00140398 3.3 0.0014038999999999998 3.3 0.0014039999999999999 0 0.00140392 0 0.00140402 3.3 0.00140394 3.3 0.00140404 0 0.0014039599999999999 0 0.00140406 3.3 0.00140398 3.3 0.00140408 0 0.0014039999999999999 0 0.0014041 3.3 0.00140402 3.3 0.00140412 0 0.0014040399999999998 0 0.00140414 3.3 0.00140406 3.3 0.00140416 0 0.0014040799999999998 0 0.0014041799999999999 3.3 0.0014041 3.3 0.0014042 0 0.00140412 0 0.00140422 3.3 0.00140414 3.3 0.00140424 0 0.00140416 0 0.00140426 3.3 0.0014041799999999999 3.3 0.00140428 0 0.0014042 0 0.0014043 3.3 0.0014042199999999999 3.3 0.00140432 0 0.00140424 0 0.00140434 3.3 0.0014042599999999998 3.3 0.00140436 0 0.00140428 0 0.00140438 3.3 0.0014042999999999998 3.3 0.0014043999999999999 0 0.00140432 0 0.00140442 3.3 0.00140434 3.3 0.00140444 0 0.00140436 0 0.00140446 3.3 0.00140438 3.3 0.00140448 0 0.0014043999999999999 0 0.0014045 3.3 0.00140442 3.3 0.00140452 0 0.0014044399999999999 0 0.00140454 3.3 0.00140446 3.3 0.00140456 0 0.0014044799999999998 0 0.0014045799999999999 3.3 0.0014045 3.3 0.0014046 0 0.0014045199999999998 0 0.0014046199999999999 3.3 0.00140454 3.3 0.00140464 0 0.00140456 0 0.00140466 3.3 0.0014045799999999999 3.3 0.00140468 0 0.0014046 0 0.0014047 3.3 0.0014046199999999999 3.3 0.00140472 0 0.00140464 0 0.00140474 3.3 0.0014046599999999998 3.3 0.00140476 0 0.00140468 0 0.00140478 3.3 0.0014046999999999998 3.3 0.0014047999999999999 0 0.00140472 0 0.00140482 3.3 0.0014047399999999998 3.3 0.0014048399999999999 0 0.00140476 0 0.00140486 3.3 0.00140478 3.3 0.00140488 0 0.0014047999999999999 0 0.0014049 3.3 0.00140482 3.3 0.00140492 0 0.0014048399999999999 0 0.00140494 3.3 0.00140486 3.3 0.00140496 0 0.0014048799999999998 0 0.00140498 3.3 0.0014049 3.3 0.001405 0 0.0014049199999999998 0 0.0014050199999999999 3.3 0.00140494 3.3 0.00140504 0 0.00140496 0 0.00140506 3.3 0.00140498 3.3 0.00140508 0 0.001405 0 0.0014051 3.3 0.0014050199999999999 3.3 0.00140512 0 0.00140504 0 0.00140514 3.3 0.0014050599999999999 3.3 0.00140516 0 0.00140508 0 0.00140518 3.3 0.0014050999999999998 3.3 0.0014052 0 0.00140512 0 0.00140522 3.3 0.0014051399999999998 3.3 0.0014052399999999999 0 0.00140516 0 0.00140526 3.3 0.00140518 3.3 0.00140528 0 0.0014052 0 0.0014053 3.3 0.00140522 3.3 0.00140532 0 0.0014052399999999999 0 0.00140534 3.3 0.00140526 3.3 0.00140536 0 0.0014052799999999999 0 0.00140538 3.3 0.0014053 3.3 0.0014054 0 0.0014053199999999998 0 0.0014054199999999999 3.3 0.00140534 3.3 0.00140544 0 0.0014053599999999998 0 0.0014054599999999999 3.3 0.00140538 3.3 0.00140548 0 0.0014054 0 0.0014055 3.3 0.0014054199999999999 3.3 0.00140552 0 0.00140544 0 0.00140554 3.3 0.0014054599999999999 3.3 0.00140556 0 0.00140548 0 0.00140558 3.3 0.0014054999999999998 3.3 0.0014056 0 0.00140552 0 0.00140562 3.3 0.0014055399999999998 3.3 0.0014056399999999999 0 0.00140556 0 0.00140566 3.3 0.0014055799999999998 3.3 0.0014056799999999999 0 0.0014056 0 0.0014057 3.3 0.00140562 3.3 0.00140572 0 0.0014056399999999999 0 0.00140574 3.3 0.00140566 3.3 0.00140576 0 0.0014056799999999999 0 0.00140578 3.3 0.0014057 3.3 0.0014058 0 0.0014057199999999998 0 0.00140582 3.3 0.00140574 3.3 0.00140584 0 0.0014057599999999998 0 0.0014058599999999999 3.3 0.00140578 3.3 0.00140588 0 0.0014058 0 0.0014059 3.3 0.00140582 3.3 0.00140592 0 0.00140584 0 0.00140594 3.3 0.0014058599999999999 3.3 0.00140596 0 0.00140588 0 0.00140598 3.3 0.0014058999999999999 3.3 0.001406 0 0.00140592 0 0.00140602 3.3 0.0014059399999999998 3.3 0.00140604 0 0.00140596 0 0.00140606 3.3 0.0014059799999999998 3.3 0.0014060799999999999 0 0.001406 0 0.0014061 3.3 0.00140602 3.3 0.00140612 0 0.00140604 0 0.00140614 3.3 0.00140606 3.3 0.00140616 0 0.0014060799999999999 0 0.00140618 3.3 0.0014061 3.3 0.0014062 0 0.0014061199999999999 0 0.00140622 3.3 0.00140614 3.3 0.00140624 0 0.0014061599999999998 0 0.0014062599999999999 3.3 0.00140618 3.3 0.00140628 0 0.0014061999999999998 0 0.0014062999999999999 3.3 0.00140622 3.3 0.00140632 0 0.00140624 0 0.00140634 3.3 0.0014062599999999999 3.3 0.00140636 0 0.00140628 0 0.00140638 3.3 0.0014062999999999999 3.3 0.0014064 0 0.00140632 0 0.00140642 3.3 0.0014063399999999998 3.3 0.00140644 0 0.00140636 0 0.00140646 3.3 0.0014063799999999998 3.3 0.0014064799999999999 0 0.0014064 0 0.0014065 3.3 0.00140642 3.3 0.00140652 0 0.00140644 0 0.00140654 3.3 0.00140646 3.3 0.00140656 0 0.0014064799999999999 0 0.00140658 3.3 0.0014065 3.3 0.0014066 0 0.0014065199999999999 0 0.00140662 3.3 0.00140654 3.3 0.00140664 0 0.0014065599999999998 0 0.00140666 3.3 0.00140658 3.3 0.00140668 0 0.0014065999999999998 0 0.0014066999999999999 3.3 0.00140662 3.3 0.00140672 0 0.00140664 0 0.00140674 3.3 0.00140666 3.3 0.00140676 0 0.00140668 0 0.00140678 3.3 0.0014066999999999999 3.3 0.0014068 0 0.00140672 0 0.00140682 3.3 0.0014067399999999999 3.3 0.00140684 0 0.00140676 0 0.00140686 3.3 0.0014067799999999998 3.3 0.00140688 0 0.0014068 0 0.0014069 3.3 0.0014068199999999998 3.3 0.0014069199999999999 0 0.00140684 0 0.00140694 3.3 0.00140686 3.3 0.00140696 0 0.00140688 0 0.00140698 3.3 0.0014069 3.3 0.001407 0 0.0014069199999999999 0 0.00140702 3.3 0.00140694 3.3 0.00140704 0 0.0014069599999999999 0 0.00140706 3.3 0.00140698 3.3 0.00140708 0 0.0014069999999999998 0 0.0014070999999999999 3.3 0.00140702 3.3 0.00140712 0 0.0014070399999999998 0 0.0014071399999999999 3.3 0.00140706 3.3 0.00140716 0 0.00140708 0 0.00140718 3.3 0.0014070999999999999 3.3 0.0014072 0 0.00140712 0 0.00140722 3.3 0.0014071399999999999 3.3 0.00140724 0 0.00140716 0 0.00140726 3.3 0.0014071799999999998 3.3 0.00140728 0 0.0014072 0 0.0014073 3.3 0.0014072199999999998 3.3 0.0014073199999999999 0 0.00140724 0 0.00140734 3.3 0.00140726 3.3 0.00140736 0 0.00140728 0 0.00140738 3.3 0.0014073 3.3 0.0014074 0 0.0014073199999999999 0 0.00140742 3.3 0.00140734 3.3 0.00140744 0 0.0014073599999999999 0 0.00140746 3.3 0.00140738 3.3 0.00140748 0 0.0014073999999999998 0 0.0014075 3.3 0.00140742 3.3 0.00140752 0 0.0014074399999999998 0 0.0014075399999999999 3.3 0.00140746 3.3 0.00140756 0 0.00140748 0 0.00140758 3.3 0.0014075 3.3 0.0014076 0 0.00140752 0 0.00140762 3.3 0.0014075399999999999 3.3 0.00140764 0 0.00140756 0 0.00140766 3.3 0.0014075799999999999 3.3 0.00140768 0 0.0014076 0 0.0014077 3.3 0.0014076199999999998 3.3 0.0014077199999999999 0 0.00140764 0 0.00140774 3.3 0.0014076599999999998 3.3 0.0014077599999999999 0 0.00140768 0 0.00140778 3.3 0.0014077 3.3 0.0014078 0 0.0014077199999999999 0 0.00140782 3.3 0.00140774 3.3 0.00140784 0 0.0014077599999999999 0 0.00140786 3.3 0.00140778 3.3 0.00140788 0 0.0014077999999999999 0 0.0014079 3.3 0.00140782 3.3 0.00140792 0 0.0014078399999999998 0 0.0014079399999999999 3.3 0.00140786 3.3 0.00140796 0 0.0014078799999999998 0 0.0014079799999999999 3.3 0.0014079 3.3 0.001408 0 0.00140792 0 0.00140802 3.3 0.0014079399999999999 3.3 0.00140804 0 0.00140796 0 0.00140806 3.3 0.0014079799999999999 3.3 0.00140808 0 0.001408 0 0.0014081 3.3 0.0014080199999999998 3.3 0.00140812 0 0.00140804 0 0.00140814 3.3 0.0014080599999999998 3.3 0.0014081599999999999 0 0.00140808 0 0.00140818 3.3 0.0014081 3.3 0.0014082 0 0.00140812 0 0.00140822 3.3 0.00140814 3.3 0.00140824 0 0.0014081599999999999 0 0.00140826 3.3 0.00140818 3.3 0.00140828 0 0.0014081999999999999 0 0.0014083 3.3 0.00140822 3.3 0.00140832 0 0.0014082399999999998 0 0.00140834 3.3 0.00140826 3.3 0.00140836 0 0.0014082799999999998 0 0.0014083799999999999 3.3 0.0014083 3.3 0.0014084 0 0.00140832 0 0.00140842 3.3 0.00140834 3.3 0.00140844 0 0.00140836 0 0.00140846 3.3 0.0014083799999999999 3.3 0.00140848 0 0.0014084 0 0.0014085 3.3 0.0014084199999999999 3.3 0.00140852 0 0.00140844 0 0.00140854 3.3 0.0014084599999999998 3.3 0.0014085599999999999 0 0.00140848 0 0.00140858 3.3 0.0014084999999999998 3.3 0.0014085999999999999 0 0.00140852 0 0.00140862 3.3 0.00140854 3.3 0.00140864 0 0.0014085599999999999 0 0.00140866 3.3 0.00140858 3.3 0.00140868 0 0.0014085999999999999 0 0.0014087 3.3 0.00140862 3.3 0.00140872 0 0.0014086399999999998 0 0.00140874 3.3 0.00140866 3.3 0.00140876 0 0.0014086799999999998 0 0.0014087799999999999 3.3 0.0014087 3.3 0.0014088 0 0.0014087199999999998 0 0.0014088199999999999 3.3 0.00140874 3.3 0.00140884 0 0.00140876 0 0.00140886 3.3 0.0014087799999999999 3.3 0.00140888 0 0.0014088 0 0.0014089 3.3 0.0014088199999999999 3.3 0.00140892 0 0.00140884 0 0.00140894 3.3 0.0014088599999999998 3.3 0.00140896 0 0.00140888 0 0.00140898 3.3 0.0014088999999999998 3.3 0.0014089999999999999 0 0.00140892 0 0.00140902 3.3 0.00140894 3.3 0.00140904 0 0.00140896 0 0.00140906 3.3 0.00140898 3.3 0.00140908 0 0.0014089999999999999 0 0.0014091 3.3 0.00140902 3.3 0.00140912 0 0.0014090399999999999 0 0.00140914 3.3 0.00140906 3.3 0.00140916 0 0.0014090799999999998 0 0.00140918 3.3 0.0014091 3.3 0.0014092 0 0.0014091199999999998 0 0.0014092199999999999 3.3 0.00140914 3.3 0.00140924 0 0.00140916 0 0.00140926 3.3 0.00140918 3.3 0.00140928 0 0.0014092 0 0.0014093 3.3 0.0014092199999999999 3.3 0.00140932 0 0.00140924 0 0.00140934 3.3 0.0014092599999999999 3.3 0.00140936 0 0.00140928 0 0.00140938 3.3 0.0014092999999999998 3.3 0.0014093999999999999 0 0.00140932 0 0.00140942 3.3 0.0014093399999999998 3.3 0.0014094399999999999 0 0.00140936 0 0.00140946 3.3 0.00140938 3.3 0.00140948 0 0.0014093999999999999 0 0.0014095 3.3 0.00140942 3.3 0.00140952 0 0.0014094399999999999 0 0.00140954 3.3 0.00140946 3.3 0.00140956 0 0.0014094799999999998 0 0.00140958 3.3 0.0014095 3.3 0.0014096 0 0.0014095199999999998 0 0.0014096199999999999 3.3 0.00140954 3.3 0.00140964 0 0.00140956 0 0.00140966 3.3 0.00140958 3.3 0.00140968 0 0.0014096 0 0.0014097 3.3 0.0014096199999999999 3.3 0.00140972 0 0.00140964 0 0.00140974 3.3 0.0014096599999999999 3.3 0.00140976 0 0.00140968 0 0.00140978 3.3 0.0014096999999999998 3.3 0.0014098 0 0.00140972 0 0.00140982 3.3 0.0014097399999999998 3.3 0.0014098399999999999 0 0.00140976 0 0.00140986 3.3 0.00140978 3.3 0.00140988 0 0.0014098 0 0.0014099 3.3 0.00140982 3.3 0.00140992 0 0.0014098399999999999 0 0.00140994 3.3 0.00140986 3.3 0.00140996 0 0.0014098799999999999 0 0.00140998 3.3 0.0014099 3.3 0.00141 0 0.0014099199999999998 0 0.00141002 3.3 0.00140994 3.3 0.00141004 0 0.0014099599999999998 0 0.0014100599999999999 3.3 0.00140998 3.3 0.00141008 0 0.00141 0 0.0014101 3.3 0.00141002 3.3 0.00141012 0 0.00141004 0 0.00141014 3.3 0.0014100599999999999 3.3 0.00141016 0 0.00141008 0 0.00141018 3.3 0.0014100999999999999 3.3 0.0014102 0 0.00141012 0 0.00141022 3.3 0.0014101399999999998 3.3 0.0014102399999999999 0 0.00141016 0 0.00141026 3.3 0.0014101799999999998 3.3 0.0014102799999999999 0 0.0014102 0 0.0014103 3.3 0.00141022 3.3 0.00141032 0 0.0014102399999999999 0 0.00141034 3.3 0.00141026 3.3 0.00141036 0 0.0014102799999999999 0 0.00141038 3.3 0.0014103 3.3 0.0014104 0 0.0014103199999999998 0 0.00141042 3.3 0.00141034 3.3 0.00141044 0 0.0014103599999999998 0 0.0014104599999999999 3.3 0.00141038 3.3 0.00141048 0 0.0014104 0 0.0014105 3.3 0.00141042 3.3 0.00141052 0 0.00141044 0 0.00141054 3.3 0.0014104599999999999 3.3 0.00141056 0 0.00141048 0 0.00141058 3.3 0.0014104999999999999 3.3 0.0014106 0 0.00141052 0 0.00141062 3.3 0.0014105399999999998 3.3 0.00141064 0 0.00141056 0 0.00141066 3.3 0.0014105799999999998 3.3 0.0014106799999999999 0 0.0014106 0 0.0014107 3.3 0.00141062 3.3 0.00141072 0 0.00141064 0 0.00141074 3.3 0.00141066 3.3 0.00141076 0 0.0014106799999999999 0 0.00141078 3.3 0.0014107 3.3 0.0014108 0 0.0014107199999999999 0 0.00141082 3.3 0.00141074 3.3 0.00141084 0 0.0014107599999999998 0 0.00141086 3.3 0.00141078 3.3 0.00141088 0 0.0014107999999999998 0 0.0014108999999999999 3.3 0.00141082 3.3 0.00141092 0 0.00141084 0 0.00141094 3.3 0.00141086 3.3 0.00141096 0 0.00141088 0 0.00141098 3.3 0.0014108999999999999 3.3 0.001411 0 0.00141092 0 0.00141102 3.3 0.0014109399999999999 3.3 0.00141104 0 0.00141096 0 0.00141106 3.3 0.0014109799999999998 3.3 0.0014110799999999999 0 0.001411 0 0.0014111 3.3 0.0014110199999999998 3.3 0.0014111199999999999 0 0.00141104 0 0.00141114 3.3 0.00141106 3.3 0.00141116 0 0.0014110799999999999 0 0.00141118 3.3 0.0014111 3.3 0.0014112 0 0.0014111199999999999 0 0.00141122 3.3 0.00141114 3.3 0.00141124 0 0.0014111599999999998 0 0.00141126 3.3 0.00141118 3.3 0.00141128 0 0.0014111999999999998 0 0.0014112999999999999 3.3 0.00141122 3.3 0.00141132 0 0.00141124 0 0.00141134 3.3 0.00141126 3.3 0.00141136 0 0.00141128 0 0.00141138 3.3 0.0014112999999999999 3.3 0.0014114 0 0.00141132 0 0.00141142 3.3 0.0014113399999999999 3.3 0.00141144 0 0.00141136 0 0.00141146 3.3 0.0014113799999999998 3.3 0.00141148 0 0.0014114 0 0.0014115 3.3 0.0014114199999999998 3.3 0.0014115199999999999 0 0.00141144 0 0.00141154 3.3 0.00141146 3.3 0.00141156 0 0.00141148 0 0.00141158 3.3 0.0014115 3.3 0.0014116 0 0.0014115199999999999 0 0.00141162 3.3 0.00141154 3.3 0.00141164 0 0.0014115599999999999 0 0.00141166 3.3 0.00141158 3.3 0.00141168 0 0.0014115999999999998 0 0.0014116999999999999 3.3 0.00141162 3.3 0.00141172 0 0.0014116399999999998 0 0.0014117399999999999 3.3 0.00141166 3.3 0.00141176 0 0.00141168 0 0.00141178 3.3 0.0014116999999999999 3.3 0.0014118 0 0.00141172 0 0.00141182 3.3 0.0014117399999999999 3.3 0.00141184 0 0.00141176 0 0.00141186 3.3 0.0014117799999999998 3.3 0.00141188 0 0.0014118 0 0.0014119 3.3 0.0014118199999999998 3.3 0.0014119199999999999 0 0.00141184 0 0.00141194 3.3 0.0014118599999999998 3.3 0.0014119599999999999 0 0.00141188 0 0.00141198 3.3 0.0014119 3.3 0.001412 0 0.0014119199999999999 0 0.00141202 3.3 0.00141194 3.3 0.00141204 0 0.0014119599999999999 0 0.00141206 3.3 0.00141198 3.3 0.00141208 0 0.0014119999999999998 0 0.0014121 3.3 0.00141202 3.3 0.00141212 0 0.0014120399999999998 0 0.0014121399999999999 3.3 0.00141206 3.3 0.00141216 0 0.00141208 0 0.00141218 3.3 0.0014121 3.3 0.0014122 0 0.00141212 0 0.00141222 3.3 0.0014121399999999999 3.3 0.00141224 0 0.00141216 0 0.00141226 3.3 0.0014121799999999999 3.3 0.00141228 0 0.0014122 0 0.0014123 3.3 0.0014122199999999998 3.3 0.00141232 0 0.00141224 0 0.00141234 3.3 0.0014122599999999998 3.3 0.0014123599999999999 0 0.00141228 0 0.00141238 3.3 0.0014123 3.3 0.0014124 0 0.00141232 0 0.00141242 3.3 0.00141234 3.3 0.00141244 0 0.0014123599999999999 0 0.00141246 3.3 0.00141238 3.3 0.00141248 0 0.0014123999999999999 0 0.0014125 3.3 0.00141242 3.3 0.00141252 0 0.0014124399999999998 0 0.0014125399999999999 3.3 0.00141246 3.3 0.00141256 0 0.0014124799999999998 0 0.0014125799999999999 3.3 0.0014125 3.3 0.0014126 0 0.00141252 0 0.00141262 3.3 0.0014125399999999999 3.3 0.00141264 0 0.00141256 0 0.00141266 3.3 0.0014125799999999999 3.3 0.00141268 0 0.0014126 0 0.0014127 3.3 0.0014126199999999998 3.3 0.00141272 0 0.00141264 0 0.00141274 3.3 0.0014126599999999998 3.3 0.0014127599999999999 0 0.00141268 0 0.00141278 3.3 0.0014126999999999998 3.3 0.0014127999999999999 0 0.00141272 0 0.00141282 3.3 0.00141274 3.3 0.00141284 0 0.0014127599999999999 0 0.00141286 3.3 0.00141278 3.3 0.00141288 0 0.0014127999999999999 0 0.0014129 3.3 0.00141282 3.3 0.00141292 0 0.0014128399999999998 0 0.00141294 3.3 0.00141286 3.3 0.00141296 0 0.0014128799999999998 0 0.0014129799999999999 3.3 0.0014129 3.3 0.001413 0 0.00141292 0 0.00141302 3.3 0.00141294 3.3 0.00141304 0 0.00141296 0 0.00141306 3.3 0.0014129799999999999 3.3 0.00141308 0 0.001413 0 0.0014131 3.3 0.0014130199999999999 3.3 0.00141312 0 0.00141304 0 0.00141314 3.3 0.0014130599999999998 3.3 0.00141316 0 0.00141308 0 0.00141318 3.3 0.0014130999999999998 3.3 0.0014131999999999999 0 0.00141312 0 0.00141322 3.3 0.00141314 3.3 0.00141324 0 0.00141316 0 0.00141326 3.3 0.00141318 3.3 0.00141328 0 0.0014131999999999999 0 0.0014133 3.3 0.00141322 3.3 0.00141332 0 0.0014132399999999999 0 0.00141334 3.3 0.00141326 3.3 0.00141336 0 0.0014132799999999998 0 0.0014133799999999999 3.3 0.0014133 3.3 0.0014134 0 0.0014133199999999998 0 0.0014134199999999999 3.3 0.00141334 3.3 0.00141344 0 0.00141336 0 0.00141346 3.3 0.0014133799999999999 3.3 0.00141348 0 0.0014134 0 0.0014135 3.3 0.0014134199999999999 3.3 0.00141352 0 0.00141344 0 0.00141354 3.3 0.0014134599999999998 3.3 0.00141356 0 0.00141348 0 0.00141358 3.3 0.0014134999999999998 3.3 0.0014135999999999999 0 0.00141352 0 0.00141362 3.3 0.00141354 3.3 0.00141364 0 0.00141356 0 0.00141366 3.3 0.00141358 3.3 0.00141368 0 0.0014135999999999999 0 0.0014137 3.3 0.00141362 3.3 0.00141372 0 0.0014136399999999999 0 0.00141374 3.3 0.00141366 3.3 0.00141376 0 0.0014136799999999998 0 0.00141378 3.3 0.0014137 3.3 0.0014138 0 0.0014137199999999998 0 0.0014138199999999999 3.3 0.00141374 3.3 0.00141384 0 0.00141376 0 0.00141386 3.3 0.00141378 3.3 0.00141388 0 0.0014138 0 0.0014139 3.3 0.0014138199999999999 3.3 0.00141392 0 0.00141384 0 0.00141394 3.3 0.0014138599999999999 3.3 0.00141396 0 0.00141388 0 0.00141398 3.3 0.0014138999999999998 3.3 0.001414 0 0.00141392 0 0.00141402 3.3 0.0014139399999999998 3.3 0.0014140399999999999 0 0.00141396 0 0.00141406 3.3 0.00141398 3.3 0.00141408 0 0.001414 0 0.0014141 3.3 0.00141402 3.3 0.00141412 0 0.0014140399999999999 0 0.00141414 3.3 0.00141406 3.3 0.00141416 0 0.0014140799999999999 0 0.00141418 3.3 0.0014141 3.3 0.0014142 0 0.0014141199999999998 0 0.0014142199999999999 3.3 0.00141414 3.3 0.00141424 0 0.0014141599999999998 0 0.0014142599999999999 3.3 0.00141418 3.3 0.00141428 0 0.0014142 0 0.0014143 3.3 0.0014142199999999999 3.3 0.00141432 0 0.00141424 0 0.00141434 3.3 0.0014142599999999999 3.3 0.00141436 0 0.00141428 0 0.00141438 3.3 0.0014142999999999998 3.3 0.0014144 0 0.00141432 0 0.00141442 3.3 0.0014143399999999998 3.3 0.0014144399999999999 0 0.00141436 0 0.00141446 3.3 0.00141438 3.3 0.00141448 0 0.0014144 0 0.0014145 3.3 0.00141442 3.3 0.00141452 0 0.0014144399999999999 0 0.00141454 3.3 0.00141446 3.3 0.00141456 0 0.0014144799999999999 0 0.00141458 3.3 0.0014145 3.3 0.0014146 0 0.0014145199999999998 0 0.00141462 3.3 0.00141454 3.3 0.00141464 0 0.0014145599999999998 0 0.0014146599999999999 3.3 0.00141458 3.3 0.00141468 0 0.0014146 0 0.0014147 3.3 0.00141462 3.3 0.00141472 0 0.00141464 0 0.00141474 3.3 0.0014146599999999999 3.3 0.00141476 0 0.00141468 0 0.00141478 3.3 0.0014146999999999999 3.3 0.0014148 0 0.00141472 0 0.00141482 3.3 0.0014147399999999998 3.3 0.0014148399999999999 0 0.00141476 0 0.00141486 3.3 0.0014147799999999998 3.3 0.0014148799999999999 0 0.0014148 0 0.0014149 3.3 0.00141482 3.3 0.00141492 0 0.0014148399999999999 0 0.00141494 3.3 0.00141486 3.3 0.00141496 0 0.0014148799999999999 0 0.00141498 3.3 0.0014149 3.3 0.001415 0 0.0014149199999999998 0 0.00141502 3.3 0.00141494 3.3 0.00141504 0 0.0014149599999999998 0 0.0014150599999999999 3.3 0.00141498 3.3 0.00141508 0 0.0014149999999999998 0 0.0014150999999999999 3.3 0.00141502 3.3 0.00141512 0 0.00141504 0 0.00141514 3.3 0.0014150599999999999 3.3 0.00141516 0 0.00141508 0 0.00141518 3.3 0.0014150999999999999 3.3 0.0014152 0 0.00141512 0 0.00141522 3.3 0.0014151399999999998 3.3 0.00141524 0 0.00141516 0 0.00141526 3.3 0.0014151799999999998 3.3 0.0014152799999999999 0 0.0014152 0 0.0014153 3.3 0.00141522 3.3 0.00141532 0 0.00141524 0 0.00141534 3.3 0.00141526 3.3 0.00141536 0 0.0014152799999999999 0 0.00141538 3.3 0.0014153 3.3 0.0014154 0 0.0014153199999999999 0 0.00141542 3.3 0.00141534 3.3 0.00141544 0 0.0014153599999999998 0 0.00141546 3.3 0.00141538 3.3 0.00141548 0 0.0014153999999999998 0 0.0014154999999999999 3.3 0.00141542 3.3 0.00141552 0 0.00141544 0 0.00141554 3.3 0.00141546 3.3 0.00141556 0 0.00141548 0 0.00141558 3.3 0.0014154999999999999 3.3 0.0014156 0 0.00141552 0 0.00141562 3.3 0.0014155399999999999 3.3 0.00141564 0 0.00141556 0 0.00141566 3.3 0.0014155799999999998 3.3 0.0014156799999999999 0 0.0014156 0 0.0014157 3.3 0.0014156199999999998 3.3 0.0014157199999999999 0 0.00141564 0 0.00141574 3.3 0.00141566 3.3 0.00141576 0 0.0014156799999999999 0 0.00141578 3.3 0.0014157 3.3 0.0014158 0 0.0014157199999999999 0 0.00141582 3.3 0.00141574 3.3 0.00141584 0 0.0014157599999999998 0 0.00141586 3.3 0.00141578 3.3 0.00141588 0 0.0014157999999999998 0 0.0014158999999999999 3.3 0.00141582 3.3 0.00141592 0 0.0014158399999999998 0 0.0014159399999999999 3.3 0.00141586 3.3 0.00141596 0 0.00141588 0 0.00141598 3.3 0.0014158999999999999 3.3 0.001416 0 0.00141592 0 0.00141602 3.3 0.0014159399999999999 3.3 0.00141604 0 0.00141596 0 0.00141606 3.3 0.0014159799999999998 3.3 0.00141608 0 0.001416 0 0.0014161 3.3 0.0014160199999999998 3.3 0.0014161199999999999 0 0.00141604 0 0.00141614 3.3 0.00141606 3.3 0.00141616 0 0.00141608 0 0.00141618 3.3 0.0014161 3.3 0.0014162 0 0.0014161199999999999 0 0.00141622 3.3 0.00141614 3.3 0.00141624 0 0.0014161599999999999 0 0.00141626 3.3 0.00141618 3.3 0.00141628 0 0.0014161999999999998 0 0.0014163 3.3 0.00141622 3.3 0.00141632 0 0.0014162399999999998 0 0.0014163399999999999 3.3 0.00141626 3.3 0.00141636 0 0.00141628 0 0.00141638 3.3 0.0014163 3.3 0.0014164 0 0.00141632 0 0.00141642 3.3 0.0014163399999999999 3.3 0.00141644 0 0.00141636 0 0.00141646 3.3 0.0014163799999999999 3.3 0.00141648 0 0.0014164 0 0.0014165 3.3 0.0014164199999999998 3.3 0.0014165199999999999 0 0.00141644 0 0.00141654 3.3 0.0014164599999999998 3.3 0.0014165599999999999 0 0.00141648 0 0.00141658 3.3 0.0014165 3.3 0.0014166 0 0.0014165199999999999 0 0.00141662 3.3 0.00141654 3.3 0.00141664 0 0.0014165599999999999 0 0.00141666 3.3 0.00141658 3.3 0.00141668 0 0.0014165999999999998 0 0.0014167 3.3 0.00141662 3.3 0.00141672 0 0.0014166399999999998 0 0.0014167399999999999 3.3 0.00141666 3.3 0.00141676 0 0.00141668 0 0.00141678 3.3 0.0014167 3.3 0.0014168 0 0.00141672 0 0.00141682 3.3 0.0014167399999999999 3.3 0.00141684 0 0.00141676 0 0.00141686 3.3 0.0014167799999999999 3.3 0.00141688 0 0.0014168 0 0.0014169 3.3 0.0014168199999999998 3.3 0.00141692 0 0.00141684 0 0.00141694 3.3 0.0014168599999999998 3.3 0.0014169599999999999 0 0.00141688 0 0.00141698 3.3 0.0014169 3.3 0.001417 0 0.00141692 0 0.00141702 3.3 0.00141694 3.3 0.00141704 0 0.0014169599999999999 0 0.00141706 3.3 0.00141698 3.3 0.00141708 0 0.0014169999999999999 0 0.0014171 3.3 0.00141702 3.3 0.00141712 0 0.0014170399999999998 0 0.00141714 3.3 0.00141706 3.3 0.00141716 0 0.0014170799999999998 0 0.0014171799999999999 3.3 0.0014171 3.3 0.0014172 0 0.00141712 0 0.00141722 3.3 0.00141714 3.3 0.00141724 0 0.00141716 0 0.00141726 3.3 0.0014171799999999999 3.3 0.00141728 0 0.0014172 0 0.0014173 3.3 0.0014172199999999999 3.3 0.00141732 0 0.00141724 0 0.00141734 3.3 0.0014172599999999998 3.3 0.0014173599999999999 0 0.00141728 0 0.00141738 3.3 0.0014172999999999998 3.3 0.0014173999999999999 0 0.00141732 0 0.00141742 3.3 0.00141734 3.3 0.00141744 0 0.0014173599999999999 0 0.00141746 3.3 0.00141738 3.3 0.00141748 0 0.0014173999999999999 0 0.0014175 3.3 0.00141742 3.3 0.00141752 0 0.0014174399999999998 0 0.00141754 3.3 0.00141746 3.3 0.00141756 0 0.0014174799999999998 0 0.0014175799999999999 3.3 0.0014175 3.3 0.0014176 0 0.00141752 0 0.00141762 3.3 0.00141754 3.3 0.00141764 0 0.00141756 0 0.00141766 3.3 0.0014175799999999999 3.3 0.00141768 0 0.0014176 0 0.0014177 3.3 0.0014176199999999999 3.3 0.00141772 0 0.00141764 0 0.00141774 3.3 0.0014176599999999998 3.3 0.00141776 0 0.00141768 0 0.00141778 3.3 0.0014176999999999998 3.3 0.0014177999999999999 0 0.00141772 0 0.00141782 3.3 0.00141774 3.3 0.00141784 0 0.00141776 0 0.00141786 3.3 0.00141778 3.3 0.00141788 0 0.0014177999999999999 0 0.0014179 3.3 0.00141782 3.3 0.00141792 0 0.0014178399999999999 0 0.00141794 3.3 0.00141786 3.3 0.00141796 0 0.0014178799999999998 0 0.0014179799999999999 3.3 0.0014179 3.3 0.001418 0 0.0014179199999999998 0 0.0014180199999999999 3.3 0.00141794 3.3 0.00141804 0 0.00141796 0 0.00141806 3.3 0.0014179799999999999 3.3 0.00141808 0 0.001418 0 0.0014181 3.3 0.0014180199999999999 3.3 0.00141812 0 0.00141804 0 0.00141814 3.3 0.0014180599999999999 3.3 0.00141816 0 0.00141808 0 0.00141818 3.3 0.0014180999999999998 3.3 0.0014181999999999999 0 0.00141812 0 0.00141822 3.3 0.0014181399999999998 3.3 0.0014182399999999999 0 0.00141816 0 0.00141826 3.3 0.00141818 3.3 0.00141828 0 0.0014181999999999999 0 0.0014183 3.3 0.00141822 3.3 0.00141832 0 0.0014182399999999999 0 0.00141834 3.3 0.00141826 3.3 0.00141836 0 0.0014182799999999998 0 0.00141838 3.3 0.0014183 3.3 0.0014184 0 0.0014183199999999998 0 0.0014184199999999999 3.3 0.00141834 3.3 0.00141844 0 0.00141836 0 0.00141846 3.3 0.00141838 3.3 0.00141848 0 0.0014184 0 0.0014185 3.3 0.0014184199999999999 3.3 0.00141852 0 0.00141844 0 0.00141854 3.3 0.0014184599999999999 3.3 0.00141856 0 0.00141848 0 0.00141858 3.3 0.0014184999999999998 3.3 0.0014186 0 0.00141852 0 0.00141862 3.3 0.0014185399999999998 3.3 0.0014186399999999999 0 0.00141856 0 0.00141866 3.3 0.00141858 3.3 0.00141868 0 0.0014186 0 0.0014187 3.3 0.00141862 3.3 0.00141872 0 0.0014186399999999999 0 0.00141874 3.3 0.00141866 3.3 0.00141876 0 0.0014186799999999999 0 0.00141878 3.3 0.0014187 3.3 0.0014188 0 0.0014187199999999998 0 0.0014188199999999999 3.3 0.00141874 3.3 0.00141884 0 0.0014187599999999998 0 0.0014188599999999999 3.3 0.00141878 3.3 0.00141888 0 0.0014188 0 0.0014189 3.3 0.0014188199999999999 3.3 0.00141892 0 0.00141884 0 0.00141894 3.3 0.0014188599999999999 3.3 0.00141896 0 0.00141888 0 0.00141898 3.3 0.0014188999999999998 3.3 0.001419 0 0.00141892 0 0.00141902 3.3 0.0014189399999999998 3.3 0.0014190399999999999 0 0.00141896 0 0.00141906 3.3 0.0014189799999999998 3.3 0.0014190799999999999 0 0.001419 0 0.0014191 3.3 0.00141902 3.3 0.00141912 0 0.0014190399999999999 0 0.00141914 3.3 0.00141906 3.3 0.00141916 0 0.0014190799999999999 0 0.00141918 3.3 0.0014191 3.3 0.0014192 0 0.0014191199999999998 0 0.00141922 3.3 0.00141914 3.3 0.00141924 0 0.0014191599999999998 0 0.0014192599999999999 3.3 0.00141918 3.3 0.00141928 0 0.0014192 0 0.0014193 3.3 0.00141922 3.3 0.00141932 0 0.00141924 0 0.00141934 3.3 0.0014192599999999999 3.3 0.00141936 0 0.00141928 0 0.00141938 3.3 0.0014192999999999999 3.3 0.0014194 0 0.00141932 0 0.00141942 3.3 0.0014193399999999998 3.3 0.00141944 0 0.00141936 0 0.00141946 3.3 0.0014193799999999998 3.3 0.0014194799999999999 0 0.0014194 0 0.0014195 3.3 0.00141942 3.3 0.00141952 0 0.00141944 0 0.00141954 3.3 0.00141946 3.3 0.00141956 0 0.0014194799999999999 0 0.00141958 3.3 0.0014195 3.3 0.0014196 0 0.0014195199999999999 0 0.00141962 3.3 0.00141954 3.3 0.00141964 0 0.0014195599999999998 0 0.0014196599999999999 3.3 0.00141958 3.3 0.00141968 0 0.0014195999999999998 0 0.0014196999999999999 3.3 0.00141962 3.3 0.00141972 0 0.00141964 0 0.00141974 3.3 0.0014196599999999999 3.3 0.00141976 0 0.00141968 0 0.00141978 3.3 0.0014196999999999999 3.3 0.0014198 0 0.00141972 0 0.00141982 3.3 0.0014197399999999998 3.3 0.00141984 0 0.00141976 0 0.00141986 3.3 0.0014197799999999998 3.3 0.0014198799999999999 0 0.0014198 0 0.0014199 3.3 0.00141982 3.3 0.00141992 0 0.00141984 0 0.00141994 3.3 0.00141986 3.3 0.00141996 0 0.0014198799999999999 0 0.00141998 3.3 0.0014199 3.3 0.00142 0 0.0014199199999999999 0 0.00142002 3.3 0.00141994 3.3 0.00142004 0 0.0014199599999999998 0 0.00142006 3.3 0.00141998 3.3 0.00142008 0 0.0014199999999999998 0 0.0014200999999999999 3.3 0.00142002 3.3 0.00142012 0 0.00142004 0 0.00142014 3.3 0.00142006 3.3 0.00142016 0 0.00142008 0 0.00142018 3.3 0.0014200999999999999 3.3 0.0014202 0 0.00142012 0 0.00142022 3.3 0.0014201399999999999 3.3 0.00142024 0 0.00142016 0 0.00142026 3.3 0.0014201799999999998 3.3 0.00142028 0 0.0014202 0 0.0014203 3.3 0.0014202199999999998 3.3 0.0014203199999999999 0 0.00142024 0 0.00142034 3.3 0.00142026 3.3 0.00142036 0 0.00142028 0 0.00142038 3.3 0.0014203 3.3 0.0014204 0 0.0014203199999999999 0 0.00142042 3.3 0.00142034 3.3 0.00142044 0 0.0014203599999999999 0 0.00142046 3.3 0.00142038 3.3 0.00142048 0 0.0014203999999999998 0 0.0014204999999999999 3.3 0.00142042 3.3 0.00142052 0 0.0014204399999999998 0 0.0014205399999999999 3.3 0.00142046 3.3 0.00142056 0 0.00142048 0 0.00142058 3.3 0.0014204999999999999 3.3 0.0014206 0 0.00142052 0 0.00142062 3.3 0.0014205399999999999 3.3 0.00142064 0 0.00142056 0 0.00142066 3.3 0.0014205799999999998 3.3 0.00142068 0 0.0014206 0 0.0014207 3.3 0.0014206199999999998 3.3 0.0014207199999999999 0 0.00142064 0 0.00142074 3.3 0.00142066 3.3 0.00142076 0 0.00142068 0 0.00142078 3.3 0.0014207 3.3 0.0014208 0 0.0014207199999999999 0 0.00142082 3.3 0.00142074 3.3 0.00142084 0 0.0014207599999999999 0 0.00142086 3.3 0.00142078 3.3 0.00142088 0 0.0014207999999999998 0 0.0014209 3.3 0.00142082 3.3 0.00142092 0 0.0014208399999999998 0 0.0014209399999999999 3.3 0.00142086 3.3 0.00142096 0 0.00142088 0 0.00142098 3.3 0.0014209 3.3 0.001421 0 0.00142092 0 0.00142102 3.3 0.0014209399999999999 3.3 0.00142104 0 0.00142096 0 0.00142106 3.3 0.0014209799999999999 3.3 0.00142108 0 0.001421 0 0.0014211 3.3 0.0014210199999999998 3.3 0.00142112 0 0.00142104 0 0.00142114 3.3 0.0014210599999999998 3.3 0.0014211599999999999 0 0.00142108 0 0.00142118 3.3 0.0014211 3.3 0.0014212 0 0.00142112 0 0.00142122 3.3 0.00142114 3.3 0.00142124 0 0.0014211599999999999 0 0.00142126 3.3 0.00142118 3.3 0.00142128 0 0.0014211999999999999 0 0.0014213 3.3 0.00142122 3.3 0.00142132 0 0.0014212399999999998 0 0.0014213399999999999 3.3 0.00142126 3.3 0.00142136 0 0.0014212799999999998 0 0.0014213799999999999 3.3 0.0014213 3.3 0.0014214 0 0.00142132 0 0.00142142 3.3 0.0014213399999999999 3.3 0.00142144 0 0.00142136 0 0.00142146 3.3 0.0014213799999999999 3.3 0.00142148 0 0.0014214 0 0.0014215 3.3 0.0014214199999999998 3.3 0.00142152 0 0.00142144 0 0.00142154 3.3 0.0014214599999999998 3.3 0.0014215599999999999 0 0.00142148 0 0.00142158 3.3 0.0014215 3.3 0.0014216 0 0.00142152 0 0.00142162 3.3 0.00142154 3.3 0.00142164 0 0.0014215599999999999 0 0.00142166 3.3 0.00142158 3.3 0.00142168 0 0.0014215999999999999 0 0.0014217 3.3 0.00142162 3.3 0.00142172 0 0.0014216399999999998 0 0.00142174 3.3 0.00142166 3.3 0.00142176 0 0.0014216799999999998 0 0.0014217799999999999 3.3 0.0014217 3.3 0.0014218 0 0.00142172 0 0.00142182 3.3 0.00142174 3.3 0.00142184 0 0.00142176 0 0.00142186 3.3 0.0014217799999999999 3.3 0.00142188 0 0.0014218 0 0.0014219 3.3 0.0014218199999999999 3.3 0.00142192 0 0.00142184 0 0.00142194 3.3 0.0014218599999999998 3.3 0.0014219599999999999 0 0.00142188 0 0.00142198 3.3 0.0014218999999999998 3.3 0.0014219999999999999 0 0.00142192 0 0.00142202 3.3 0.00142194 3.3 0.00142204 0 0.0014219599999999999 0 0.00142206 3.3 0.00142198 3.3 0.00142208 0 0.0014219999999999999 0 0.0014221 3.3 0.00142202 3.3 0.00142212 0 0.0014220399999999998 0 0.00142214 3.3 0.00142206 3.3 0.00142216 0 0.0014220799999999998 0 0.0014221799999999999 3.3 0.0014221 3.3 0.0014222 0 0.0014221199999999998 0 0.0014222199999999999 3.3 0.00142214 3.3 0.00142224 0 0.00142216 0 0.00142226 3.3 0.0014221799999999999 3.3 0.00142228 0 0.0014222 0 0.0014223 3.3 0.0014222199999999999 3.3 0.00142232 0 0.00142224 0 0.00142234 3.3 0.0014222599999999998 3.3 0.00142236 0 0.00142228 0 0.00142238 3.3 0.0014222999999999998 3.3 0.0014223999999999999 0 0.00142232 0 0.00142242 3.3 0.00142234 3.3 0.00142244 0 0.00142236 0 0.00142246 3.3 0.00142238 3.3 0.00142248 0 0.0014223999999999999 0 0.0014225 3.3 0.00142242 3.3 0.00142252 0 0.0014224399999999999 0 0.00142254 3.3 0.00142246 3.3 0.00142256 0 0.0014224799999999998 0 0.00142258 3.3 0.0014225 3.3 0.0014226 0 0.0014225199999999998 0 0.0014226199999999999 3.3 0.00142254 3.3 0.00142264 0 0.00142256 0 0.00142266 3.3 0.00142258 3.3 0.00142268 0 0.0014226 0 0.0014227 3.3 0.0014226199999999999 3.3 0.00142272 0 0.00142264 0 0.00142274 3.3 0.0014226599999999999 3.3 0.00142276 0 0.00142268 0 0.00142278 3.3 0.0014226999999999998 3.3 0.0014227999999999999 0 0.00142272 0 0.00142282 3.3 0.0014227399999999998 3.3 0.0014228399999999999 0 0.00142276 0 0.00142286 3.3 0.00142278 3.3 0.00142288 0 0.0014227999999999999 0 0.0014229 3.3 0.00142282 3.3 0.00142292 0 0.0014228399999999999 0 0.00142294 3.3 0.00142286 3.3 0.00142296 0 0.0014228799999999998 0 0.00142298 3.3 0.0014229 3.3 0.001423 0 0.0014229199999999998 0 0.0014230199999999999 3.3 0.00142294 3.3 0.00142304 0 0.0014229599999999998 0 0.0014230599999999999 3.3 0.00142298 3.3 0.00142308 0 0.001423 0 0.0014231 3.3 0.0014230199999999999 3.3 0.00142312 0 0.00142304 0 0.00142314 3.3 0.0014230599999999999 3.3 0.00142316 0 0.00142308 0 0.00142318 3.3 0.0014230999999999998 3.3 0.0014232 0 0.00142312 0 0.00142322 3.3 0.0014231399999999998 3.3 0.0014232399999999999 0 0.00142316 0 0.00142326 3.3 0.00142318 3.3 0.00142328 0 0.0014232 0 0.0014233 3.3 0.00142322 3.3 0.00142332 0 0.0014232399999999999 0 0.00142334 3.3 0.00142326 3.3 0.00142336 0 0.0014232799999999999 0 0.00142338 3.3 0.0014233 3.3 0.0014234 0 0.0014233199999999998 0 0.00142342 3.3 0.00142334 3.3 0.00142344 0 0.0014233599999999998 0 0.0014234599999999999 3.3 0.00142338 3.3 0.00142348 0 0.0014234 0 0.0014235 3.3 0.00142342 3.3 0.00142352 0 0.00142344 0 0.00142354 3.3 0.0014234599999999999 3.3 0.00142356 0 0.00142348 0 0.00142358 3.3 0.0014234999999999999 3.3 0.0014236 0 0.00142352 0 0.00142362 3.3 0.0014235399999999998 3.3 0.0014236399999999999 0 0.00142356 0 0.00142366 3.3 0.0014235799999999998 3.3 0.0014236799999999999 0 0.0014236 0 0.0014237 3.3 0.00142362 3.3 0.00142372 0 0.0014236399999999999 0 0.00142374 3.3 0.00142366 3.3 0.00142376 0 0.0014236799999999999 0 0.00142378 3.3 0.0014237 3.3 0.0014238 0 0.0014237199999999998 0 0.00142382 3.3 0.00142374 3.3 0.00142384 0 0.0014237599999999998 0 0.0014238599999999999 3.3 0.00142378 3.3 0.00142388 0 0.0014238 0 0.0014239 3.3 0.00142382 3.3 0.00142392 0 0.00142384 0 0.00142394 3.3 0.0014238599999999999 3.3 0.00142396 0 0.00142388 0 0.00142398 3.3 0.0014238999999999999 3.3 0.001424 0 0.00142392 0 0.00142402 3.3 0.0014239399999999998 3.3 0.00142404 0 0.00142396 0 0.00142406 3.3 0.0014239799999999998 3.3 0.0014240799999999999 0 0.001424 0 0.0014241 3.3 0.00142402 3.3 0.00142412 0 0.00142404 0 0.00142414 3.3 0.00142406 3.3 0.00142416 0 0.0014240799999999999 0 0.00142418 3.3 0.0014241 3.3 0.0014242 0 0.0014241199999999999 0 0.00142422 3.3 0.00142414 3.3 0.00142424 0 0.0014241599999999998 0 0.00142426 3.3 0.00142418 3.3 0.00142428 0 0.0014241999999999998 0 0.0014242999999999999 3.3 0.00142422 3.3 0.00142432 0 0.00142424 0 0.00142434 3.3 0.00142426 3.3 0.00142436 0 0.00142428 0 0.00142438 3.3 0.0014242999999999999 3.3 0.0014244 0 0.00142432 0 0.00142442 3.3 0.0014243399999999999 3.3 0.00142444 0 0.00142436 0 0.00142446 3.3 0.0014243799999999998 3.3 0.0014244799999999999 0 0.0014244 0 0.0014245 3.3 0.0014244199999999998 3.3 0.0014245199999999999 0 0.00142444 0 0.00142454 3.3 0.00142446 3.3 0.00142456 0 0.0014244799999999999 0 0.00142458 3.3 0.0014245 3.3 0.0014246 0 0.0014245199999999999 0 0.00142462 3.3 0.00142454 3.3 0.00142464 0 0.0014245599999999998 0 0.00142466 3.3 0.00142458 3.3 0.00142468 0 0.0014245999999999998 0 0.0014246999999999999 3.3 0.00142462 3.3 0.00142472 0 0.00142464 0 0.00142474 3.3 0.00142466 3.3 0.00142476 0 0.00142468 0 0.00142478 3.3 0.0014246999999999999 3.3 0.0014248 0 0.00142472 0 0.00142482 3.3 0.0014247399999999999 3.3 0.00142484 0 0.00142476 0 0.00142486 3.3 0.0014247799999999998 3.3 0.00142488 0 0.0014248 0 0.0014249 3.3 0.0014248199999999998 3.3 0.0014249199999999999 0 0.00142484 0 0.00142494 3.3 0.00142486 3.3 0.00142496 0 0.00142488 0 0.00142498 3.3 0.0014249 3.3 0.001425 0 0.0014249199999999999 0 0.00142502 3.3 0.00142494 3.3 0.00142504 0 0.0014249599999999999 0 0.00142506 3.3 0.00142498 3.3 0.00142508 0 0.0014249999999999998 0 0.0014250999999999999 3.3 0.00142502 3.3 0.00142512 0 0.0014250399999999998 0 0.0014251399999999999 3.3 0.00142506 3.3 0.00142516 0 0.00142508 0 0.00142518 3.3 0.0014250999999999999 3.3 0.0014252 0 0.00142512 0 0.00142522 3.3 0.0014251399999999999 3.3 0.00142524 0 0.00142516 0 0.00142526 3.3 0.0014251799999999998 3.3 0.00142528 0 0.0014252 0 0.0014253 3.3 0.0014252199999999998 3.3 0.0014253199999999999 0 0.00142524 0 0.00142534 3.3 0.0014252599999999998 3.3 0.0014253599999999999 0 0.00142528 0 0.00142538 3.3 0.0014253 3.3 0.0014254 0 0.0014253199999999999 0 0.00142542 3.3 0.00142534 3.3 0.00142544 0 0.0014253599999999999 0 0.00142546 3.3 0.00142538 3.3 0.00142548 0 0.0014253999999999998 0 0.0014255 3.3 0.00142542 3.3 0.00142552 0 0.0014254399999999998 0 0.0014255399999999999 3.3 0.00142546 3.3 0.00142556 0 0.00142548 0 0.00142558 3.3 0.0014255 3.3 0.0014256 0 0.00142552 0 0.00142562 3.3 0.0014255399999999999 3.3 0.00142564 0 0.00142556 0 0.00142566 3.3 0.0014255799999999999 3.3 0.00142568 0 0.0014256 0 0.0014257 3.3 0.0014256199999999998 3.3 0.00142572 0 0.00142564 0 0.00142574 3.3 0.0014256599999999998 3.3 0.0014257599999999999 0 0.00142568 0 0.00142578 3.3 0.0014257 3.3 0.0014258 0 0.00142572 0 0.00142582 3.3 0.00142574 3.3 0.00142584 0 0.0014257599999999999 0 0.00142586 3.3 0.00142578 3.3 0.00142588 0 0.0014257999999999999 0 0.0014259 3.3 0.00142582 3.3 0.00142592 0 0.0014258399999999998 0 0.0014259399999999999 3.3 0.00142586 3.3 0.00142596 0 0.0014258799999999998 0 0.0014259799999999999 3.3 0.0014259 3.3 0.001426 0 0.00142592 0 0.00142602 3.3 0.0014259399999999999 3.3 0.00142604 0 0.00142596 0 0.00142606 3.3 0.0014259799999999999 3.3 0.00142608 0 0.001426 0 0.0014261 3.3 0.0014260199999999998 3.3 0.00142612 0 0.00142604 0 0.00142614 3.3 0.0014260599999999998 3.3 0.0014261599999999999 0 0.00142608 0 0.00142618 3.3 0.0014260999999999998 3.3 0.0014261999999999999 0 0.00142612 0 0.00142622 3.3 0.00142614 3.3 0.00142624 0 0.0014261599999999999 0 0.00142626 3.3 0.00142618 3.3 0.00142628 0 0.0014261999999999999 0 0.0014263 3.3 0.00142622 3.3 0.00142632 0 0.0014262399999999998 0 0.00142634 3.3 0.00142626 3.3 0.00142636 0 0.0014262799999999998 0 0.0014263799999999999 3.3 0.0014263 3.3 0.0014264 0 0.00142632 0 0.00142642 3.3 0.00142634 3.3 0.00142644 0 0.00142636 0 0.00142646 3.3 0.0014263799999999999 3.3 0.00142648 0 0.0014264 0 0.0014265 3.3 0.0014264199999999999 3.3 0.00142652 0 0.00142644 0 0.00142654 3.3 0.0014264599999999998 3.3 0.00142656 0 0.00142648 0 0.00142658 3.3 0.0014264999999999998 3.3 0.0014265999999999999 0 0.00142652 0 0.00142662 3.3 0.00142654 3.3 0.00142664 0 0.00142656 0 0.00142666 3.3 0.00142658 3.3 0.00142668 0 0.0014265999999999999 0 0.0014267 3.3 0.00142662 3.3 0.00142672 0 0.0014266399999999999 0 0.00142674 3.3 0.00142666 3.3 0.00142676 0 0.0014266799999999998 0 0.0014267799999999999 3.3 0.0014267 3.3 0.0014268 0 0.0014267199999999998 0 0.0014268199999999999 3.3 0.00142674 3.3 0.00142684 0 0.00142676 0 0.00142686 3.3 0.0014267799999999999 3.3 0.00142688 0 0.0014268 0 0.0014269 3.3 0.0014268199999999999 3.3 0.00142692 0 0.00142684 0 0.00142694 3.3 0.0014268599999999998 3.3 0.00142696 0 0.00142688 0 0.00142698 3.3 0.0014268999999999998 3.3 0.0014269999999999999 0 0.00142692 0 0.00142702 3.3 0.00142694 3.3 0.00142704 0 0.00142696 0 0.00142706 3.3 0.00142698 3.3 0.00142708 0 0.0014269999999999999 0 0.0014271 3.3 0.00142702 3.3 0.00142712 0 0.0014270399999999999 0 0.00142714 3.3 0.00142706 3.3 0.00142716 0 0.0014270799999999998 0 0.00142718 3.3 0.0014271 3.3 0.0014272 0 0.0014271199999999998 0 0.0014272199999999999 3.3 0.00142714 3.3 0.00142724 0 0.00142716 0 0.00142726 3.3 0.00142718 3.3 0.00142728 0 0.0014272 0 0.0014273 3.3 0.0014272199999999999 3.3 0.00142732 0 0.00142724 0 0.00142734 3.3 0.0014272599999999999 3.3 0.00142736 0 0.00142728 0 0.00142738 3.3 0.0014272999999999998 3.3 0.0014274 0 0.00142732 0 0.00142742 3.3 0.0014273399999999998 3.3 0.0014274399999999999 0 0.00142736 0 0.00142746 3.3 0.00142738 3.3 0.00142748 0 0.0014274 0 0.0014275 3.3 0.00142742 3.3 0.00142752 0 0.0014274399999999999 0 0.00142754 3.3 0.00142746 3.3 0.00142756 0 0.0014274799999999999 0 0.00142758 3.3 0.0014275 3.3 0.0014276 0 0.0014275199999999998 0 0.0014276199999999999 3.3 0.00142754 3.3 0.00142764 0 0.0014275599999999998 0 0.0014276599999999999 3.3 0.00142758 3.3 0.00142768 0 0.0014276 0 0.0014277 3.3 0.0014276199999999999 3.3 0.00142772 0 0.00142764 0 0.00142774 3.3 0.0014276599999999999 3.3 0.00142776 0 0.00142768 0 0.00142778 3.3 0.0014276999999999998 3.3 0.0014278 0 0.00142772 0 0.00142782 3.3 0.0014277399999999998 3.3 0.0014278399999999999 0 0.00142776 0 0.00142786 3.3 0.00142778 3.3 0.00142788 0 0.0014278 0 0.0014279 3.3 0.00142782 3.3 0.00142792 0 0.0014278399999999999 0 0.00142794 3.3 0.00142786 3.3 0.00142796 0 0.0014278799999999999 0 0.00142798 3.3 0.0014279 3.3 0.001428 0 0.0014279199999999998 0 0.00142802 3.3 0.00142794 3.3 0.00142804 0 0.0014279599999999998 0 0.0014280599999999999 3.3 0.00142798 3.3 0.00142808 0 0.001428 0 0.0014281 3.3 0.00142802 3.3 0.00142812 0 0.00142804 0 0.00142814 3.3 0.0014280599999999999 3.3 0.00142816 0 0.00142808 0 0.00142818 3.3 0.0014280999999999999 3.3 0.0014282 0 0.00142812 0 0.00142822 3.3 0.0014281399999999998 3.3 0.0014282399999999999 0 0.00142816 0 0.00142826 3.3 0.0014281799999999998 3.3 0.0014282799999999999 0 0.0014282 0 0.0014283 3.3 0.00142822 3.3 0.00142832 0 0.0014282399999999999 0 0.00142834 3.3 0.00142826 3.3 0.00142836 0 0.0014282799999999999 0 0.00142838 3.3 0.0014283 3.3 0.0014284 0 0.0014283199999999999 0 0.00142842 3.3 0.00142834 3.3 0.00142844 0 0.0014283599999999998 0 0.0014284599999999999 3.3 0.00142838 3.3 0.00142848 0 0.0014283999999999998 0 0.0014284999999999999 3.3 0.00142842 3.3 0.00142852 0 0.00142844 0 0.00142854 3.3 0.0014284599999999999 3.3 0.00142856 0 0.00142848 0 0.00142858 3.3 0.0014284999999999999 3.3 0.0014286 0 0.00142852 0 0.00142862 3.3 0.0014285399999999998 3.3 0.00142864 0 0.00142856 0 0.00142866 3.3 0.0014285799999999998 3.3 0.0014286799999999999 0 0.0014286 0 0.0014287 3.3 0.00142862 3.3 0.00142872 0 0.00142864 0 0.00142874 3.3 0.00142866 3.3 0.00142876 0 0.0014286799999999999 0 0.00142878 3.3 0.0014287 3.3 0.0014288 0 0.0014287199999999999 0 0.00142882 3.3 0.00142874 3.3 0.00142884 0 0.0014287599999999998 0 0.00142886 3.3 0.00142878 3.3 0.00142888 0 0.0014287999999999998 0 0.0014288999999999999 3.3 0.00142882 3.3 0.00142892 0 0.00142884 0 0.00142894 3.3 0.00142886 3.3 0.00142896 0 0.00142888 0 0.00142898 3.3 0.0014288999999999999 3.3 0.001429 0 0.00142892 0 0.00142902 3.3 0.0014289399999999999 3.3 0.00142904 0 0.00142896 0 0.00142906 3.3 0.0014289799999999998 3.3 0.0014290799999999999 0 0.001429 0 0.0014291 3.3 0.0014290199999999998 3.3 0.0014291199999999999 0 0.00142904 0 0.00142914 3.3 0.00142906 3.3 0.00142916 0 0.0014290799999999999 0 0.00142918 3.3 0.0014291 3.3 0.0014292 0 0.0014291199999999999 0 0.00142922 3.3 0.00142914 3.3 0.00142924 0 0.0014291599999999998 0 0.00142926 3.3 0.00142918 3.3 0.00142928 0 0.0014291999999999998 0 0.0014292999999999999 3.3 0.00142922 3.3 0.00142932 0 0.0014292399999999998 0 0.0014293399999999999 3.3 0.00142926 3.3 0.00142936 0 0.00142928 0 0.00142938 3.3 0.0014292999999999999 3.3 0.0014294 0 0.00142932 0 0.00142942 3.3 0.0014293399999999999 3.3 0.00142944 0 0.00142936 0 0.00142946 3.3 0.0014293799999999998 3.3 0.00142948 0 0.0014294 0 0.0014295 3.3 0.0014294199999999998 3.3 0.0014295199999999999 0 0.00142944 0 0.00142954 3.3 0.00142946 3.3 0.00142956 0 0.00142948 0 0.00142958 3.3 0.0014295 3.3 0.0014296 0 0.0014295199999999999 0 0.00142962 3.3 0.00142954 3.3 0.00142964 0 0.0014295599999999999 0 0.00142966 3.3 0.00142958 3.3 0.00142968 0 0.0014295999999999998 0 0.0014297 3.3 0.00142962 3.3 0.00142972 0 0.0014296399999999998 0 0.0014297399999999999 3.3 0.00142966 3.3 0.00142976 0 0.00142968 0 0.00142978 3.3 0.0014297 3.3 0.0014298 0 0.00142972 0 0.00142982 3.3 0.0014297399999999999 3.3 0.00142984 0 0.00142976 0 0.00142986 3.3 0.0014297799999999999 3.3 0.00142988 0 0.0014298 0 0.0014299 3.3 0.0014298199999999998 3.3 0.0014299199999999999 0 0.00142984 0 0.00142994 3.3 0.0014298599999999998 3.3 0.0014299599999999999 0 0.00142988 0 0.00142998 3.3 0.0014299 3.3 0.00143 0 0.0014299199999999999 0 0.00143002 3.3 0.00142994 3.3 0.00143004 0 0.0014299599999999999 0 0.00143006 3.3 0.00142998 3.3 0.00143008 0 0.0014299999999999998 0 0.0014301 3.3 0.00143002 3.3 0.00143012 0 0.0014300399999999998 0 0.0014301399999999999 3.3 0.00143006 3.3 0.00143016 0 0.0014300799999999998 0 0.0014301799999999999 3.3 0.0014301 3.3 0.0014302 0 0.00143012 0 0.00143022 3.3 0.0014301399999999999 3.3 0.00143024 0 0.00143016 0 0.00143026 3.3 0.0014301799999999999 3.3 0.00143028 0 0.0014302 0 0.0014303 3.3 0.0014302199999999998 3.3 0.00143032 0 0.00143024 0 0.00143034 3.3 0.0014302599999999998 3.3 0.0014303599999999999 0 0.00143028 0 0.00143038 3.3 0.0014303 3.3 0.0014304 0 0.00143032 0 0.00143042 3.3 0.00143034 3.3 0.00143044 0 0.0014303599999999999 0 0.00143046 3.3 0.00143038 3.3 0.00143048 0 0.0014303999999999999 0 0.0014305 3.3 0.00143042 3.3 0.00143052 0 0.0014304399999999998 0 0.00143054 3.3 0.00143046 3.3 0.00143056 0 0.0014304799999999998 0 0.0014305799999999999 3.3 0.0014305 3.3 0.0014306 0 0.00143052 0 0.00143062 3.3 0.00143054 3.3 0.00143064 0 0.00143056 0 0.00143066 3.3 0.0014305799999999999 3.3 0.00143068 0 0.0014306 0 0.0014307 3.3 0.0014306199999999999 3.3 0.00143072 0 0.00143064 0 0.00143074 3.3 0.0014306599999999998 3.3 0.0014307599999999999 0 0.00143068 0 0.00143078 3.3 0.0014306999999999998 3.3 0.0014307999999999999 0 0.00143072 0 0.00143082 3.3 0.00143074 3.3 0.00143084 0 0.0014307599999999999 0 0.00143086 3.3 0.00143078 3.3 0.00143088 0 0.0014307999999999999 0 0.0014309 3.3 0.00143082 3.3 0.00143092 0 0.0014308399999999998 0 0.00143094 3.3 0.00143086 3.3 0.00143096 0 0.0014308799999999998 0 0.0014309799999999999 3.3 0.0014309 3.3 0.001431 0 0.00143092 0 0.00143102 3.3 0.00143094 3.3 0.00143104 0 0.00143096 0 0.00143106 3.3 0.0014309799999999999 3.3 0.00143108 0 0.001431 0 0.0014311 3.3 0.0014310199999999999 3.3 0.00143112 0 0.00143104 0 0.00143114 3.3 0.0014310599999999998 3.3 0.00143116 0 0.00143108 0 0.00143118 3.3 0.0014310999999999998 3.3 0.0014311999999999999 0 0.00143112 0 0.00143122 3.3 0.00143114 3.3 0.00143124 0 0.00143116 0 0.00143126 3.3 0.00143118 3.3 0.00143128 0 0.0014311999999999999 0 0.0014313 3.3 0.00143122 3.3 0.00143132 0 0.0014312399999999999 0 0.00143134 3.3 0.00143126 3.3 0.00143136 0 0.0014312799999999998 0 0.00143138 3.3 0.0014313 3.3 0.0014314 0 0.0014313199999999998 0 0.0014314199999999999 3.3 0.00143134 3.3 0.00143144 0 0.00143136 0 0.00143146 3.3 0.00143138 3.3 0.00143148 0 0.0014314 0 0.0014315 3.3 0.0014314199999999999 3.3 0.00143152 0 0.00143144 0 0.00143154 3.3 0.0014314599999999999 3.3 0.00143156 0 0.00143148 0 0.00143158 3.3 0.0014314999999999998 3.3 0.0014315999999999999 0 0.00143152 0 0.00143162 3.3 0.0014315399999999998 3.3 0.0014316399999999999 0 0.00143156 0 0.00143166 3.3 0.00143158 3.3 0.00143168 0 0.0014315999999999999 0 0.0014317 3.3 0.00143162 3.3 0.00143172 0 0.0014316399999999999 0 0.00143174 3.3 0.00143166 3.3 0.00143176 0 0.0014316799999999998 0 0.00143178 3.3 0.0014317 3.3 0.0014318 0 0.0014317199999999998 0 0.0014318199999999999 3.3 0.00143174 3.3 0.00143184 0 0.00143176 0 0.00143186 3.3 0.00143178 3.3 0.00143188 0 0.0014318 0 0.0014319 3.3 0.0014318199999999999 3.3 0.00143192 0 0.00143184 0 0.00143194 3.3 0.0014318599999999999 3.3 0.00143196 0 0.00143188 0 0.00143198 3.3 0.0014318999999999998 3.3 0.001432 0 0.00143192 0 0.00143202 3.3 0.0014319399999999998 3.3 0.0014320399999999999 0 0.00143196 0 0.00143206 3.3 0.00143198 3.3 0.00143208 0 0.001432 0 0.0014321 3.3 0.00143202 3.3 0.00143212 0 0.0014320399999999999 0 0.00143214 3.3 0.00143206 3.3 0.00143216 0 0.0014320799999999999 0 0.00143218 3.3 0.0014321 3.3 0.0014322 0 0.0014321199999999998 0 0.0014322199999999999 3.3 0.00143214 3.3 0.00143224 0 0.0014321599999999998 0 0.0014322599999999999 3.3 0.00143218 3.3 0.00143228 0 0.0014322 0 0.0014323 3.3 0.0014322199999999999 3.3 0.00143232 0 0.00143224 0 0.00143234 3.3 0.0014322599999999999 3.3 0.00143236 0 0.00143228 0 0.00143238 3.3 0.0014322999999999998 3.3 0.0014324 0 0.00143232 0 0.00143242 3.3 0.0014323399999999998 3.3 0.0014324399999999999 0 0.00143236 0 0.00143246 3.3 0.0014323799999999998 3.3 0.0014324799999999999 0 0.0014324 0 0.0014325 3.3 0.00143242 3.3 0.00143252 0 0.0014324399999999999 0 0.00143254 3.3 0.00143246 3.3 0.00143256 0 0.0014324799999999999 0 0.00143258 3.3 0.0014325 3.3 0.0014326 0 0.0014325199999999998 0 0.00143262 3.3 0.00143254 3.3 0.00143264 0 0.0014325599999999998 0 0.0014326599999999999 3.3 0.00143258 3.3 0.00143268 0 0.0014326 0 0.0014327 3.3 0.00143262 3.3 0.00143272 0 0.00143264 0 0.00143274 3.3 0.0014326599999999999 3.3 0.00143276 0 0.00143268 0 0.00143278 3.3 0.0014326999999999999 3.3 0.0014328 0 0.00143272 0 0.00143282 3.3 0.0014327399999999998 3.3 0.00143284 0 0.00143276 0 0.00143286 3.3 0.0014327799999999998 3.3 0.0014328799999999999 0 0.0014328 0 0.0014329 3.3 0.00143282 3.3 0.00143292 0 0.00143284 0 0.00143294 3.3 0.00143286 3.3 0.00143296 0 0.0014328799999999999 0 0.00143298 3.3 0.0014329 3.3 0.001433 0 0.0014329199999999999 0 0.00143302 3.3 0.00143294 3.3 0.00143304 0 0.0014329599999999998 0 0.0014330599999999999 3.3 0.00143298 3.3 0.00143308 0 0.0014329999999999998 0 0.0014330999999999999 3.3 0.00143302 3.3 0.00143312 0 0.00143304 0 0.00143314 3.3 0.0014330599999999999 3.3 0.00143316 0 0.00143308 0 0.00143318 3.3 0.0014330999999999999 3.3 0.0014332 0 0.00143312 0 0.00143322 3.3 0.0014331399999999998 3.3 0.00143324 0 0.00143316 0 0.00143326 3.3 0.0014331799999999998 3.3 0.0014332799999999999 0 0.0014332 0 0.0014333 3.3 0.0014332199999999998 3.3 0.0014333199999999999 0 0.00143324 0 0.00143334 3.3 0.00143326 3.3 0.00143336 0 0.0014332799999999999 0 0.00143338 3.3 0.0014333 3.3 0.0014334 0 0.0014333199999999999 0 0.00143342 3.3 0.00143334 3.3 0.00143344 0 0.0014333599999999998 0 0.00143346 3.3 0.00143338 3.3 0.00143348 0 0.0014333999999999998 0 0.0014334999999999999 3.3 0.00143342 3.3 0.00143352 0 0.00143344 0 0.00143354 3.3 0.00143346 3.3 0.00143356 0 0.00143348 0 0.00143358 3.3 0.0014334999999999999 3.3 0.0014336 0 0.00143352 0 0.00143362 3.3 0.0014335399999999999 3.3 0.00143364 0 0.00143356 0 0.00143366 3.3 0.0014335799999999998 3.3 0.00143368 0 0.0014336 0 0.0014337 3.3 0.0014336199999999998 3.3 0.0014337199999999999 0 0.00143364 0 0.00143374 3.3 0.00143366 3.3 0.00143376 0 0.00143368 0 0.00143378 3.3 0.0014337 3.3 0.0014338 0 0.0014337199999999999 0 0.00143382 3.3 0.00143374 3.3 0.00143384 0 0.0014337599999999999 0 0.00143386 3.3 0.00143378 3.3 0.00143388 0 0.0014337999999999998 0 0.0014338999999999999 3.3 0.00143382 3.3 0.00143392 0 0.0014338399999999998 0 0.0014339399999999999 3.3 0.00143386 3.3 0.00143396 0 0.00143388 0 0.00143398 3.3 0.0014338999999999999 3.3 0.001434 0 0.00143392 0 0.00143402 3.3 0.0014339399999999999 3.3 0.00143404 0 0.00143396 0 0.00143406 3.3 0.0014339799999999998 3.3 0.00143408 0 0.001434 0 0.0014341 3.3 0.0014340199999999998 3.3 0.0014341199999999999 0 0.00143404 0 0.00143414 3.3 0.00143406 3.3 0.00143416 0 0.00143408 0 0.00143418 3.3 0.0014341 3.3 0.0014342 0 0.0014341199999999999 0 0.00143422 3.3 0.00143414 3.3 0.00143424 0 0.0014341599999999999 0 0.00143426 3.3 0.00143418 3.3 0.00143428 0 0.0014341999999999998 0 0.0014343 3.3 0.00143422 3.3 0.00143432 0 0.0014342399999999998 0 0.0014343399999999999 3.3 0.00143426 3.3 0.00143436 0 0.00143428 0 0.00143438 3.3 0.0014343 3.3 0.0014344 0 0.00143432 0 0.00143442 3.3 0.0014343399999999999 3.3 0.00143444 0 0.00143436 0 0.00143446 3.3 0.0014343799999999999 3.3 0.00143448 0 0.0014344 0 0.0014345 3.3 0.0014344199999999998 3.3 0.00143452 0 0.00143444 0 0.00143454 3.3 0.0014344599999999998 3.3 0.0014345599999999999 0 0.00143448 0 0.00143458 3.3 0.0014345 3.3 0.0014346 0 0.00143452 0 0.00143462 3.3 0.00143454 3.3 0.00143464 0 0.0014345599999999999 0 0.00143466 3.3 0.00143458 3.3 0.00143468 0 0.0014345999999999999 0 0.0014347 3.3 0.00143462 3.3 0.00143472 0 0.0014346399999999998 0 0.0014347399999999999 3.3 0.00143466 3.3 0.00143476 0 0.0014346799999999998 0 0.0014347799999999999 3.3 0.0014347 3.3 0.0014348 0 0.00143472 0 0.00143482 3.3 0.0014347399999999999 3.3 0.00143484 0 0.00143476 0 0.00143486 3.3 0.0014347799999999999 3.3 0.00143488 0 0.0014348 0 0.0014349 3.3 0.0014348199999999998 3.3 0.00143492 0 0.00143484 0 0.00143494 3.3 0.0014348599999999998 3.3 0.0014349599999999999 0 0.00143488 0 0.00143498 3.3 0.0014349 3.3 0.001435 0 0.00143492 0 0.00143502 3.3 0.00143494 3.3 0.00143504 0 0.0014349599999999999 0 0.00143506 3.3 0.00143498 3.3 0.00143508 0 0.0014349999999999999 0 0.0014351 3.3 0.00143502 3.3 0.00143512 0 0.0014350399999999998 0 0.00143514 3.3 0.00143506 3.3 0.00143516 0 0.0014350799999999998 0 0.0014351799999999999 3.3 0.0014351 3.3 0.0014352 0 0.00143512 0 0.00143522 3.3 0.00143514 3.3 0.00143524 0 0.00143516 0 0.00143526 3.3 0.0014351799999999999 3.3 0.00143528 0 0.0014352 0 0.0014353 3.3 0.0014352199999999999 3.3 0.00143532 0 0.00143524 0 0.00143534 3.3 0.0014352599999999998 3.3 0.0014353599999999999 0 0.00143528 0 0.00143538 3.3 0.0014352999999999998 3.3 0.0014353999999999999 0 0.00143532 0 0.00143542 3.3 0.00143534 3.3 0.00143544 0 0.0014353599999999999 0 0.00143546 3.3 0.00143538 3.3 0.00143548 0 0.0014353999999999999 0 0.0014355 3.3 0.00143542 3.3 0.00143552 0 0.0014354399999999998 0 0.00143554 3.3 0.00143546 3.3 0.00143556 0 0.0014354799999999998 0 0.0014355799999999999 3.3 0.0014355 3.3 0.0014356 0 0.0014355199999999998 0 0.0014356199999999999 3.3 0.00143554 3.3 0.00143564 0 0.00143556 0 0.00143566 3.3 0.0014355799999999999 3.3 0.00143568 0 0.0014356 0 0.0014357 3.3 0.0014356199999999999 3.3 0.00143572 0 0.00143564 0 0.00143574 3.3 0.0014356599999999998 3.3 0.00143576 0 0.00143568 0 0.00143578 3.3 0.0014356999999999998 3.3 0.0014357999999999999 0 0.00143572 0 0.00143582 3.3 0.00143574 3.3 0.00143584 0 0.00143576 0 0.00143586 3.3 0.00143578 3.3 0.00143588 0 0.0014357999999999999 0 0.0014359 3.3 0.00143582 3.3 0.00143592 0 0.0014358399999999999 0 0.00143594 3.3 0.00143586 3.3 0.00143596 0 0.0014358799999999998 0 0.00143598 3.3 0.0014359 3.3 0.001436 0 0.0014359199999999998 0 0.0014360199999999999 3.3 0.00143594 3.3 0.00143604 0 0.00143596 0 0.00143606 3.3 0.00143598 3.3 0.00143608 0 0.001436 0 0.0014361 3.3 0.0014360199999999999 3.3 0.00143612 0 0.00143604 0 0.00143614 3.3 0.0014360599999999999 3.3 0.00143616 0 0.00143608 0 0.00143618 3.3 0.0014360999999999998 3.3 0.0014361999999999999 0 0.00143612 0 0.00143622 3.3 0.0014361399999999998 3.3 0.0014362399999999999 0 0.00143616 0 0.00143626 3.3 0.00143618 3.3 0.00143628 0 0.0014361999999999999 0 0.0014363 3.3 0.00143622 3.3 0.00143632 0 0.0014362399999999999 0 0.00143634 3.3 0.00143626 3.3 0.00143636 0 0.0014362799999999998 0 0.00143638 3.3 0.0014363 3.3 0.0014364 0 0.0014363199999999998 0 0.0014364199999999999 3.3 0.00143634 3.3 0.00143644 0 0.0014363599999999998 0 0.0014364599999999999 3.3 0.00143638 3.3 0.00143648 0 0.0014364 0 0.0014365 3.3 0.0014364199999999999 3.3 0.00143652 0 0.00143644 0 0.00143654 3.3 0.0014364599999999999 3.3 0.00143656 0 0.00143648 0 0.00143658 3.3 0.0014364999999999998 3.3 0.0014366 0 0.00143652 0 0.00143662 3.3 0.0014365399999999998 3.3 0.0014366399999999999 0 0.00143656 0 0.00143666 3.3 0.00143658 3.3 0.00143668 0 0.0014366 0 0.0014367 3.3 0.00143662 3.3 0.00143672 0 0.0014366399999999999 0 0.00143674 3.3 0.00143666 3.3 0.00143676 0 0.0014366799999999999 0 0.00143678 3.3 0.0014367 3.3 0.0014368 0 0.0014367199999999998 0 0.00143682 3.3 0.00143674 3.3 0.00143684 0 0.0014367599999999998 0 0.0014368599999999999 3.3 0.00143678 3.3 0.00143688 0 0.0014368 0 0.0014369 3.3 0.00143682 3.3 0.00143692 0 0.00143684 0 0.00143694 3.3 0.0014368599999999999 3.3 0.00143696 0 0.00143688 0 0.00143698 3.3 0.0014368999999999999 3.3 0.001437 0 0.00143692 0 0.00143702 3.3 0.0014369399999999998 3.3 0.0014370399999999999 0 0.00143696 0 0.00143706 3.3 0.0014369799999999998 3.3 0.0014370799999999999 0 0.001437 0 0.0014371 3.3 0.00143702 3.3 0.00143712 0 0.0014370399999999999 0 0.00143714 3.3 0.00143706 3.3 0.00143716 0 0.0014370799999999999 0 0.00143718 3.3 0.0014371 3.3 0.0014372 0 0.0014371199999999998 0 0.00143722 3.3 0.00143714 3.3 0.00143724 0 0.0014371599999999998 0 0.0014372599999999999 3.3 0.00143718 3.3 0.00143728 0 0.0014372 0 0.0014373 3.3 0.00143722 3.3 0.00143732 0 0.00143724 0 0.00143734 3.3 0.0014372599999999999 3.3 0.00143736 0 0.00143728 0 0.00143738 3.3 0.0014372999999999999 3.3 0.0014374 0 0.00143732 0 0.00143742 3.3 0.0014373399999999998 3.3 0.00143744 0 0.00143736 0 0.00143746 3.3 0.0014373799999999998 3.3 0.0014374799999999999 0 0.0014374 0 0.0014375 3.3 0.00143742 3.3 0.00143752 0 0.00143744 0 0.00143754 3.3 0.00143746 3.3 0.00143756 0 0.0014374799999999999 0 0.00143758 3.3 0.0014375 3.3 0.0014376 0 0.0014375199999999999 0 0.00143762 3.3 0.00143754 3.3 0.00143764 0 0.0014375599999999998 0 0.00143766 3.3 0.00143758 3.3 0.00143768 0 0.0014375999999999998 0 0.0014376999999999999 3.3 0.00143762 3.3 0.00143772 0 0.00143764 0 0.00143774 3.3 0.00143766 3.3 0.00143776 0 0.00143768 0 0.00143778 3.3 0.0014376999999999999 3.3 0.0014378 0 0.00143772 0 0.00143782 3.3 0.0014377399999999999 3.3 0.00143784 0 0.00143776 0 0.00143786 3.3 0.0014377799999999998 3.3 0.0014378799999999999 0 0.0014378 0 0.0014379 3.3 0.0014378199999999998 3.3 0.0014379199999999999 0 0.00143784 0 0.00143794 3.3 0.00143786 3.3 0.00143796 0 0.0014378799999999999 0 0.00143798 3.3 0.0014379 3.3 0.001438 0 0.0014379199999999999 0 0.00143802 3.3 0.00143794 3.3 0.00143804 0 0.0014379599999999998 0 0.00143806 3.3 0.00143798 3.3 0.00143808 0 0.0014379999999999998 0 0.0014380999999999999 3.3 0.00143802 3.3 0.00143812 0 0.00143804 0 0.00143814 3.3 0.00143806 3.3 0.00143816 0 0.00143808 0 0.00143818 3.3 0.0014380999999999999 3.3 0.0014382 0 0.00143812 0 0.00143822 3.3 0.0014381399999999999 3.3 0.00143824 0 0.00143816 0 0.00143826 3.3 0.0014381799999999998 3.3 0.00143828 0 0.0014382 0 0.0014383 3.3 0.0014382199999999998 3.3 0.0014383199999999999 0 0.00143824 0 0.00143834 3.3 0.00143826 3.3 0.00143836 0 0.00143828 0 0.00143838 3.3 0.0014383 3.3 0.0014384 0 0.0014383199999999999 0 0.00143842 3.3 0.00143834 3.3 0.00143844 0 0.0014383599999999999 0 0.00143846 3.3 0.00143838 3.3 0.00143848 0 0.0014383999999999998 0 0.0014385 3.3 0.00143842 3.3 0.00143852 0 0.0014384399999999998 0 0.0014385399999999999 3.3 0.00143846 3.3 0.00143856 0 0.00143848 0 0.00143858 3.3 0.0014385 3.3 0.0014386 0 0.00143852 0 0.00143862 3.3 0.0014385399999999999 3.3 0.00143864 0 0.00143856 0 0.00143866 3.3 0.0014385799999999999 3.3 0.00143868 0 0.0014386 0 0.0014387 3.3 0.0014386199999999998 3.3 0.0014387199999999999 0 0.00143864 0 0.00143874 3.3 0.0014386599999999998 3.3 0.0014387599999999999 0 0.00143868 0 0.00143878 3.3 0.0014387 3.3 0.0014388 0 0.0014387199999999999 0 0.00143882 3.3 0.00143874 3.3 0.00143884 0 0.0014387599999999999 0 0.00143886 3.3 0.00143878 3.3 0.00143888 0 0.0014387999999999998 0 0.0014389 3.3 0.00143882 3.3 0.00143892 0 0.0014388399999999998 0 0.0014389399999999999 3.3 0.00143886 3.3 0.00143896 0 0.00143888 0 0.00143898 3.3 0.0014389 3.3 0.001439 0 0.00143892 0 0.00143902 3.3 0.0014389399999999999 3.3 0.00143904 0 0.00143896 0 0.00143906 3.3 0.0014389799999999999 3.3 0.00143908 0 0.001439 0 0.0014391 3.3 0.0014390199999999998 3.3 0.00143912 0 0.00143904 0 0.00143914 3.3 0.0014390599999999998 3.3 0.0014391599999999999 0 0.00143908 0 0.00143918 3.3 0.0014391 3.3 0.0014392 0 0.00143912 0 0.00143922 3.3 0.00143914 3.3 0.00143924 0 0.0014391599999999999 0 0.00143926 3.3 0.00143918 3.3 0.00143928 0 0.0014391999999999999 0 0.0014393 3.3 0.00143922 3.3 0.00143932 0 0.0014392399999999998 0 0.0014393399999999999 3.3 0.00143926 3.3 0.00143936 0 0.0014392799999999998 0 0.0014393799999999999 3.3 0.0014393 3.3 0.0014394 0 0.00143932 0 0.00143942 3.3 0.0014393399999999999 3.3 0.00143944 0 0.00143936 0 0.00143946 3.3 0.0014393799999999999 3.3 0.00143948 0 0.0014394 0 0.0014395 3.3 0.0014394199999999998 3.3 0.00143952 0 0.00143944 0 0.00143954 3.3 0.0014394599999999998 3.3 0.0014395599999999999 0 0.00143948 0 0.00143958 3.3 0.0014394999999999998 3.3 0.0014395999999999999 0 0.00143952 0 0.00143962 3.3 0.00143954 3.3 0.00143964 0 0.0014395599999999999 0 0.00143966 3.3 0.00143958 3.3 0.00143968 0 0.0014395999999999999 0 0.0014397 3.3 0.00143962 3.3 0.00143972 0 0.0014396399999999998 0 0.00143974 3.3 0.00143966 3.3 0.00143976 0 0.0014396799999999998 0 0.0014397799999999999 3.3 0.0014397 3.3 0.0014398 0 0.00143972 0 0.00143982 3.3 0.00143974 3.3 0.00143984 0 0.00143976 0 0.00143986 3.3 0.0014397799999999999 3.3 0.00143988 0 0.0014398 0 0.0014399 3.3 0.0014398199999999999 3.3 0.00143992 0 0.00143984 0 0.00143994 3.3 0.0014398599999999998 3.3 0.00143996 0 0.00143988 0 0.00143998 3.3 0.0014398999999999998 3.3 0.0014399999999999999 0 0.00143992 0 0.00144002 3.3 0.00143994 3.3 0.00144004 0 0.00143996 0 0.00144006 3.3 0.00143998 3.3 0.00144008 0 0.0014399999999999999 0 0.0014401 3.3 0.00144002 3.3 0.00144012 0 0.0014400399999999999 0 0.00144014 3.3 0.00144006 3.3 0.00144016 0 0.0014400799999999998 0 0.0014401799999999999 3.3 0.0014401 3.3 0.0014402 0 0.0014401199999999998 0 0.0014402199999999999 3.3 0.00144014 3.3 0.00144024 0 0.00144016 0 0.00144026 3.3 0.0014401799999999999 3.3 0.00144028 0 0.0014402 0 0.0014403 3.3 0.0014402199999999999 3.3 0.00144032 0 0.00144024 0 0.00144034 3.3 0.0014402599999999998 3.3 0.00144036 0 0.00144028 0 0.00144038 3.3 0.0014402999999999998 3.3 0.0014403999999999999 0 0.00144032 0 0.00144042 3.3 0.0014403399999999998 3.3 0.0014404399999999999 0 0.00144036 0 0.00144046 3.3 0.00144038 3.3 0.00144048 0 0.0014403999999999999 0 0.0014405 3.3 0.00144042 3.3 0.00144052 0 0.0014404399999999999 0 0.00144054 3.3 0.00144046 3.3 0.00144056 0 0.0014404799999999998 0 0.00144058 3.3 0.0014405 3.3 0.0014406 0 0.0014405199999999998 0 0.0014406199999999999 3.3 0.00144054 3.3 0.00144064 0 0.00144056 0 0.00144066 3.3 0.00144058 3.3 0.00144068 0 0.0014406 0 0.0014407 3.3 0.0014406199999999999 3.3 0.00144072 0 0.00144064 0 0.00144074 3.3 0.0014406599999999999 3.3 0.00144076 0 0.00144068 0 0.00144078 3.3 0.0014406999999999998 3.3 0.0014408 0 0.00144072 0 0.00144082 3.3 0.0014407399999999998 3.3 0.0014408399999999999 0 0.00144076 0 0.00144086 3.3 0.00144078 3.3 0.00144088 0 0.0014408 0 0.0014409 3.3 0.00144082 3.3 0.00144092 0 0.0014408399999999999 0 0.00144094 3.3 0.00144086 3.3 0.00144096 0 0.0014408799999999999 0 0.00144098 3.3 0.0014409 3.3 0.001441 0 0.0014409199999999998 0 0.0014410199999999999 3.3 0.00144094 3.3 0.00144104 0 0.0014409599999999998 0 0.0014410599999999999 3.3 0.00144098 3.3 0.00144108 0 0.001441 0 0.0014411 3.3 0.0014410199999999999 3.3 0.00144112 0 0.00144104 0 0.00144114 3.3 0.0014410599999999999 3.3 0.00144116 0 0.00144108 0 0.00144118 3.3 0.0014410999999999998 3.3 0.0014412 0 0.00144112 0 0.00144122 3.3 0.0014411399999999998 3.3 0.0014412399999999999 0 0.00144116 0 0.00144126 3.3 0.00144118 3.3 0.00144128 0 0.0014412 0 0.0014413 3.3 0.00144122 3.3 0.00144132 0 0.0014412399999999999 0 0.00144134 3.3 0.00144126 3.3 0.00144136 0 0.0014412799999999999 0 0.00144138 3.3 0.0014413 3.3 0.0014414 0 0.0014413199999999998 0 0.00144142 3.3 0.00144134 3.3 0.00144144 0 0.0014413599999999998 0 0.0014414599999999999 3.3 0.00144138 3.3 0.00144148 0 0.0014414 0 0.0014415 3.3 0.00144142 3.3 0.00144152 0 0.00144144 0 0.00144154 3.3 0.0014414599999999999 3.3 0.00144156 0 0.00144148 0 0.00144158 3.3 0.0014414999999999999 3.3 0.0014416 0 0.00144152 0 0.00144162 3.3 0.0014415399999999998 3.3 0.00144164 0 0.00144156 0 0.00144166 3.3 0.0014415799999999998 3.3 0.0014416799999999999 0 0.0014416 0 0.0014417 3.3 0.00144162 3.3 0.00144172 0 0.00144164 0 0.00144174 3.3 0.00144166 3.3 0.00144176 0 0.0014416799999999999 0 0.00144178 3.3 0.0014417 3.3 0.0014418 0 0.0014417199999999999 0 0.00144182 3.3 0.00144174 3.3 0.00144184 0 0.0014417599999999998 0 0.0014418599999999999 3.3 0.00144178 3.3 0.00144188 0 0.0014417999999999998 0 0.0014418999999999999 3.3 0.00144182 3.3 0.00144192 0 0.00144184 0 0.00144194 3.3 0.0014418599999999999 3.3 0.00144196 0 0.00144188 0 0.00144198 3.3 0.0014418999999999999 3.3 0.001442 0 0.00144192 0 0.00144202 3.3 0.0014419399999999998 3.3 0.00144204 0 0.00144196 0 0.00144206 3.3 0.0014419799999999998 3.3 0.0014420799999999999 0 0.001442 0 0.0014421 3.3 0.00144202 3.3 0.00144212 0 0.00144204 0 0.00144214 3.3 0.00144206 3.3 0.00144216 0 0.0014420799999999999 0 0.00144218 3.3 0.0014421 3.3 0.0014422 0 0.0014421199999999999 0 0.00144222 3.3 0.00144214 3.3 0.00144224 0 0.0014421599999999998 0 0.00144226 3.3 0.00144218 3.3 0.00144228 0 0.0014421999999999998 0 0.0014422999999999999 3.3 0.00144222 3.3 0.00144232 0 0.00144224 0 0.00144234 3.3 0.00144226 3.3 0.00144236 0 0.00144228 0 0.00144238 3.3 0.0014422999999999999 3.3 0.0014424 0 0.00144232 0 0.00144242 3.3 0.0014423399999999999 3.3 0.00144244 0 0.00144236 0 0.00144246 3.3 0.0014423799999999998 3.3 0.0014424799999999999 0 0.0014424 0 0.0014425 3.3 0.0014424199999999998 3.3 0.0014425199999999999 0 0.00144244 0 0.00144254 3.3 0.00144246 3.3 0.00144256 0 0.0014424799999999999 0 0.00144258 3.3 0.0014425 3.3 0.0014426 0 0.0014425199999999999 0 0.00144262 3.3 0.00144254 3.3 0.00144264 0 0.0014425599999999998 0 0.00144266 3.3 0.00144258 3.3 0.00144268 0 0.0014425999999999998 0 0.0014426999999999999 3.3 0.00144262 3.3 0.00144272 0 0.0014426399999999998 0 0.0014427399999999999 3.3 0.00144266 3.3 0.00144276 0 0.00144268 0 0.00144278 3.3 0.0014426999999999999 3.3 0.0014428 0 0.00144272 0 0.00144282 3.3 0.0014427399999999999 3.3 0.00144284 0 0.00144276 0 0.00144286 3.3 0.0014427799999999998 3.3 0.00144288 0 0.0014428 0 0.0014429 3.3 0.0014428199999999998 3.3 0.0014429199999999999 0 0.00144284 0 0.00144294 3.3 0.00144286 3.3 0.00144296 0 0.00144288 0 0.00144298 3.3 0.0014429 3.3 0.001443 0 0.0014429199999999999 0 0.00144302 3.3 0.00144294 3.3 0.00144304 0 0.0014429599999999999 0 0.00144306 3.3 0.00144298 3.3 0.00144308 0 0.0014429999999999998 0 0.0014431 3.3 0.00144302 3.3 0.00144312 0 0.0014430399999999998 0 0.0014431399999999999 3.3 0.00144306 3.3 0.00144316 0 0.00144308 0 0.00144318 3.3 0.0014431 3.3 0.0014432 0 0.00144312 0 0.00144322 3.3 0.0014431399999999999 3.3 0.00144324 0 0.00144316 0 0.00144326 3.3 0.0014431799999999999 3.3 0.00144328 0 0.0014432 0 0.0014433 3.3 0.0014432199999999998 3.3 0.0014433199999999999 0 0.00144324 0 0.00144334 3.3 0.0014432599999999998 3.3 0.0014433599999999999 0 0.00144328 0 0.00144338 3.3 0.0014433 3.3 0.0014434 0 0.0014433199999999999 0 0.00144342 3.3 0.00144334 3.3 0.00144344 0 0.0014433599999999999 0 0.00144346 3.3 0.00144338 3.3 0.00144348 0 0.0014433999999999998 0 0.0014435 3.3 0.00144342 3.3 0.00144352 0 0.0014434399999999998 0 0.0014435399999999999 3.3 0.00144346 3.3 0.00144356 0 0.0014434799999999998 0 0.0014435799999999999 3.3 0.0014435 3.3 0.0014436 0 0.00144352 0 0.00144362 3.3 0.0014435399999999999 3.3 0.00144364 0 0.00144356 0 0.00144366 3.3 0.0014435799999999999 3.3 0.00144368 0 0.0014436 0 0.0014437 3.3 0.0014436199999999998 3.3 0.00144372 0 0.00144364 0 0.00144374 3.3 0.0014436599999999998 3.3 0.0014437599999999999 0 0.00144368 0 0.00144378 3.3 0.0014437 3.3 0.0014438 0 0.00144372 0 0.00144382 3.3 0.00144374 3.3 0.00144384 0 0.0014437599999999999 0 0.00144386 3.3 0.00144378 3.3 0.00144388 0 0.0014437999999999999 0 0.0014439 3.3 0.00144382 3.3 0.00144392 0 0.0014438399999999998 0 0.00144394 3.3 0.00144386 3.3 0.00144396 0 0.0014438799999999998 0 0.0014439799999999999 3.3 0.0014439 3.3 0.001444 0 0.00144392 0 0.00144402 3.3 0.00144394 3.3 0.00144404 0 0.00144396 0 0.00144406 3.3 0.0014439799999999999 3.3 0.00144408 0 0.001444 0 0.0014441 3.3 0.0014440199999999999 3.3 0.00144412 0 0.00144404 0 0.00144414 3.3 0.0014440599999999998 3.3 0.0014441599999999999 0 0.00144408 0 0.00144418 3.3 0.0014440999999999998 3.3 0.0014441999999999999 0 0.00144412 0 0.00144422 3.3 0.00144414 3.3 0.00144424 0 0.0014441599999999999 0 0.00144426 3.3 0.00144418 3.3 0.00144428 0 0.0014441999999999999 0 0.0014443 3.3 0.00144422 3.3 0.00144432 0 0.0014442399999999998 0 0.00144434 3.3 0.00144426 3.3 0.00144436 0 0.0014442799999999998 0 0.0014443799999999999 3.3 0.0014443 3.3 0.0014444 0 0.00144432 0 0.00144442 3.3 0.00144434 3.3 0.00144444 0 0.00144436 0 0.00144446 3.3 0.0014443799999999999 3.3 0.00144448 0 0.0014444 0 0.0014445 3.3 0.0014444199999999999 3.3 0.00144452 0 0.00144444 0 0.00144454 3.3 0.0014444599999999998 3.3 0.00144456 0 0.00144448 0 0.00144458 3.3 0.0014444999999999998 3.3 0.0014445999999999999 0 0.00144452 0 0.00144462 3.3 0.00144454 3.3 0.00144464 0 0.00144456 0 0.00144466 3.3 0.00144458 3.3 0.00144468 0 0.0014445999999999999 0 0.0014447 3.3 0.00144462 3.3 0.00144472 0 0.0014446399999999999 0 0.00144474 3.3 0.00144466 3.3 0.00144476 0 0.0014446799999999998 0 0.00144478 3.3 0.0014447 3.3 0.0014448 0 0.0014447199999999998 0 0.0014448199999999999 3.3 0.00144474 3.3 0.00144484 0 0.00144476 0 0.00144486 3.3 0.00144478 3.3 0.00144488 0 0.0014448 0 0.0014449 3.3 0.0014448199999999999 3.3 0.00144492 0 0.00144484 0 0.00144494 3.3 0.0014448599999999999 3.3 0.00144496 0 0.00144488 0 0.00144498 3.3 0.0014448999999999998 3.3 0.0014449999999999999 0 0.00144492 0 0.00144502 3.3 0.0014449399999999998 3.3 0.0014450399999999999 0 0.00144496 0 0.00144506 3.3 0.00144498 3.3 0.00144508 0 0.0014449999999999999 0 0.0014451 3.3 0.00144502 3.3 0.00144512 0 0.0014450399999999999 0 0.00144514 3.3 0.00144506 3.3 0.00144516 0 0.0014450799999999998 0 0.00144518 3.3 0.0014451 3.3 0.0014452 0 0.0014451199999999998 0 0.0014452199999999999 3.3 0.00144514 3.3 0.00144524 0 0.00144516 0 0.00144526 3.3 0.00144518 3.3 0.00144528 0 0.0014452 0 0.0014453 3.3 0.0014452199999999999 3.3 0.00144532 0 0.00144524 0 0.00144534 3.3 0.0014452599999999999 3.3 0.00144536 0 0.00144528 0 0.00144538 3.3 0.0014452999999999998 3.3 0.0014454 0 0.00144532 0 0.00144542 3.3 0.0014453399999999998 3.3 0.0014454399999999999 0 0.00144536 0 0.00144546 3.3 0.00144538 3.3 0.00144548 0 0.0014454 0 0.0014455 3.3 0.00144542 3.3 0.00144552 0 0.0014454399999999999 0 0.00144554 3.3 0.00144546 3.3 0.00144556 0 0.0014454799999999999 0 0.00144558 3.3 0.0014455 3.3 0.0014456 0 0.0014455199999999998 0 0.0014456199999999999 3.3 0.00144554 3.3 0.00144564 0 0.0014455599999999998 0 0.0014456599999999999 3.3 0.00144558 3.3 0.00144568 0 0.0014456 0 0.0014457 3.3 0.0014456199999999999 3.3 0.00144572 0 0.00144564 0 0.00144574 3.3 0.0014456599999999999 3.3 0.00144576 0 0.00144568 0 0.00144578 3.3 0.0014456999999999998 3.3 0.0014458 0 0.00144572 0 0.00144582 3.3 0.0014457399999999998 3.3 0.0014458399999999999 0 0.00144576 0 0.00144586 3.3 0.0014457799999999998 3.3 0.0014458799999999999 0 0.0014458 0 0.0014459 3.3 0.00144582 3.3 0.00144592 0 0.0014458399999999999 0 0.00144594 3.3 0.00144586 3.3 0.00144596 0 0.0014458799999999999 0 0.00144598 3.3 0.0014459 3.3 0.001446 0 0.0014459199999999998 0 0.00144602 3.3 0.00144594 3.3 0.00144604 0 0.0014459599999999998 0 0.0014460599999999999 3.3 0.00144598 3.3 0.00144608 0 0.001446 0 0.0014461 3.3 0.00144602 3.3 0.00144612 0 0.00144604 0 0.00144614 3.3 0.0014460599999999999 3.3 0.00144616 0 0.00144608 0 0.00144618 3.3 0.0014460999999999999 3.3 0.0014462 0 0.00144612 0 0.00144622 3.3 0.0014461399999999998 3.3 0.00144624 0 0.00144616 0 0.00144626 3.3 0.0014461799999999998 3.3 0.0014462799999999999 0 0.0014462 0 0.0014463 3.3 0.00144622 3.3 0.00144632 0 0.00144624 0 0.00144634 3.3 0.00144626 3.3 0.00144636 0 0.0014462799999999999 0 0.00144638 3.3 0.0014463 3.3 0.0014464 0 0.0014463199999999999 0 0.00144642 3.3 0.00144634 3.3 0.00144644 0 0.0014463599999999998 0 0.0014464599999999999 3.3 0.00144638 3.3 0.00144648 0 0.0014463999999999998 0 0.0014464999999999999 3.3 0.00144642 3.3 0.00144652 0 0.00144644 0 0.00144654 3.3 0.0014464599999999999 3.3 0.00144656 0 0.00144648 0 0.00144658 3.3 0.0014464999999999999 3.3 0.0014466 0 0.00144652 0 0.00144662 3.3 0.0014465399999999998 3.3 0.00144664 0 0.00144656 0 0.00144666 3.3 0.0014465799999999998 3.3 0.0014466799999999999 0 0.0014466 0 0.0014467 3.3 0.0014466199999999998 3.3 0.0014467199999999999 0 0.00144664 0 0.00144674 3.3 0.00144666 3.3 0.00144676 0 0.0014466799999999999 0 0.00144678 3.3 0.0014467 3.3 0.0014468 0 0.0014467199999999999 0 0.00144682 3.3 0.00144674 3.3 0.00144684 0 0.0014467599999999998 0 0.00144686 3.3 0.00144678 3.3 0.00144688 0 0.0014467999999999998 0 0.0014468999999999999 3.3 0.00144682 3.3 0.00144692 0 0.00144684 0 0.00144694 3.3 0.00144686 3.3 0.00144696 0 0.00144688 0 0.00144698 3.3 0.0014468999999999999 3.3 0.001447 0 0.00144692 0 0.00144702 3.3 0.0014469399999999999 3.3 0.00144704 0 0.00144696 0 0.00144706 3.3 0.0014469799999999998 3.3 0.00144708 0 0.001447 0 0.0014471 3.3 0.0014470199999999998 3.3 0.0014471199999999999 0 0.00144704 0 0.00144714 3.3 0.00144706 3.3 0.00144716 0 0.00144708 0 0.00144718 3.3 0.0014471 3.3 0.0014472 0 0.0014471199999999999 0 0.00144722 3.3 0.00144714 3.3 0.00144724 0 0.0014471599999999999 0 0.00144726 3.3 0.00144718 3.3 0.00144728 0 0.0014471999999999998 0 0.0014472999999999999 3.3 0.00144722 3.3 0.00144732 0 0.0014472399999999998 0 0.0014473399999999999 3.3 0.00144726 3.3 0.00144736 0 0.00144728 0 0.00144738 3.3 0.0014472999999999999 3.3 0.0014474 0 0.00144732 0 0.00144742 3.3 0.0014473399999999999 3.3 0.00144744 0 0.00144736 0 0.00144746 3.3 0.0014473799999999998 3.3 0.00144748 0 0.0014474 0 0.0014475 3.3 0.0014474199999999998 3.3 0.0014475199999999999 0 0.00144744 0 0.00144754 3.3 0.00144746 3.3 0.00144756 0 0.00144748 0 0.00144758 3.3 0.0014475 3.3 0.0014476 0 0.0014475199999999999 0 0.00144762 3.3 0.00144754 3.3 0.00144764 0 0.0014475599999999999 0 0.00144766 3.3 0.00144758 3.3 0.00144768 0 0.0014475999999999998 0 0.0014477 3.3 0.00144762 3.3 0.00144772 0 0.0014476399999999998 0 0.0014477399999999999 3.3 0.00144766 3.3 0.00144776 0 0.00144768 0 0.00144778 3.3 0.0014477 3.3 0.0014478 0 0.00144772 0 0.00144782 3.3 0.0014477399999999999 3.3 0.00144784 0 0.00144776 0 0.00144786 3.3 0.0014477799999999999 3.3 0.00144788 0 0.0014478 0 0.0014479 3.3 0.0014478199999999998 3.3 0.00144792 0 0.00144784 0 0.00144794 3.3 0.0014478599999999998 3.3 0.0014479599999999999 0 0.00144788 0 0.00144798 3.3 0.0014479 3.3 0.001448 0 0.00144792 0 0.00144802 3.3 0.00144794 3.3 0.00144804 0 0.0014479599999999999 0 0.00144806 3.3 0.00144798 3.3 0.00144808 0 0.0014479999999999999 0 0.0014481 3.3 0.00144802 3.3 0.00144812 0 0.0014480399999999998 0 0.0014481399999999999 3.3 0.00144806 3.3 0.00144816 0 0.0014480799999999998 0 0.0014481799999999999 3.3 0.0014481 3.3 0.0014482 0 0.00144812 0 0.00144822 3.3 0.0014481399999999999 3.3 0.00144824 0 0.00144816 0 0.00144826 3.3 0.0014481799999999999 3.3 0.00144828 0 0.0014482 0 0.0014483 3.3 0.0014482199999999998 3.3 0.00144832 0 0.00144824 0 0.00144834 3.3 0.0014482599999999998 3.3 0.0014483599999999999 0 0.00144828 0 0.00144838 3.3 0.0014483 3.3 0.0014484 0 0.00144832 0 0.00144842 3.3 0.00144834 3.3 0.00144844 0 0.0014483599999999999 0 0.00144846 3.3 0.00144838 3.3 0.00144848 0 0.0014483999999999999 0 0.0014485 3.3 0.00144842 3.3 0.00144852 0 0.0014484399999999998 0 0.00144854 3.3 0.00144846 3.3 0.00144856 0 0.0014484799999999998 0 0.0014485799999999999 3.3 0.0014485 3.3 0.0014486 0 0.00144852 0 0.00144862 3.3 0.00144854 3.3 0.00144864 0 0.00144856 0 0.00144866 3.3 0.0014485799999999999 3.3 0.00144868 0 0.0014486 0 0.0014487 3.3 0.0014486199999999999 3.3 0.00144872 0 0.00144864 0 0.00144874 3.3 0.0014486599999999998 3.3 0.00144876 0 0.00144868 0 0.00144878 3.3 0.0014486999999999998 3.3 0.0014487999999999999 0 0.00144872 0 0.00144882 3.3 0.00144874 3.3 0.00144884 0 0.00144876 0 0.00144886 3.3 0.00144878 3.3 0.00144888 0 0.0014487999999999999 0 0.0014489 3.3 0.00144882 3.3 0.00144892 0 0.0014488399999999999 0 0.00144894 3.3 0.00144886 3.3 0.00144896 0 0.0014488799999999998 0 0.0014489799999999999 3.3 0.0014489 3.3 0.001449 0 0.0014489199999999998 0 0.0014490199999999999 3.3 0.00144894 3.3 0.00144904 0 0.00144896 0 0.00144906 3.3 0.0014489799999999999 3.3 0.00144908 0 0.001449 0 0.0014491 3.3 0.0014490199999999999 3.3 0.00144912 0 0.00144904 0 0.00144914 3.3 0.0014490599999999998 3.3 0.00144916 0 0.00144908 0 0.00144918 3.3 0.0014490999999999998 3.3 0.0014491999999999999 0 0.00144912 0 0.00144922 3.3 0.00144914 3.3 0.00144924 0 0.00144916 0 0.00144926 3.3 0.00144918 3.3 0.00144928 0 0.0014491999999999999 0 0.0014493 3.3 0.00144922 3.3 0.00144932 0 0.0014492399999999999 0 0.00144934 3.3 0.00144926 3.3 0.00144936 0 0.0014492799999999998 0 0.00144938 3.3 0.0014493 3.3 0.0014494 0 0.0014493199999999998 0 0.0014494199999999999 3.3 0.00144934 3.3 0.00144944 0 0.00144936 0 0.00144946 3.3 0.00144938 3.3 0.00144948 0 0.0014494 0 0.0014495 3.3 0.0014494199999999999 3.3 0.00144952 0 0.00144944 0 0.00144954 3.3 0.0014494599999999999 3.3 0.00144956 0 0.00144948 0 0.00144958 3.3 0.0014494999999999998 3.3 0.0014495999999999999 0 0.00144952 0 0.00144962 3.3 0.0014495399999999998 3.3 0.0014496399999999999 0 0.00144956 0 0.00144966 3.3 0.00144958 3.3 0.00144968 0 0.0014495999999999999 0 0.0014497 3.3 0.00144962 3.3 0.00144972 0 0.0014496399999999999 0 0.00144974 3.3 0.00144966 3.3 0.00144976 0 0.0014496799999999998 0 0.00144978 3.3 0.0014497 3.3 0.0014498 0 0.0014497199999999998 0 0.0014498199999999999 3.3 0.00144974 3.3 0.00144984 0 0.0014497599999999998 0 0.0014498599999999999 3.3 0.00144978 3.3 0.00144988 0 0.0014498 0 0.0014499 3.3 0.0014498199999999999 3.3 0.00144992 0 0.00144984 0 0.00144994 3.3 0.0014498599999999999 3.3 0.00144996 0 0.00144988 0 0.00144998 3.3 0.0014498999999999998 3.3 0.00145 0 0.00144992 0 0.00145002 3.3 0.0014499399999999998 3.3 0.0014500399999999999 0 0.00144996 0 0.00145006 3.3 0.00144998 3.3 0.00145008 0 0.00145 0 0.0014501 3.3 0.00145002 3.3 0.00145012 0 0.0014500399999999999 0 0.00145014 3.3 0.00145006 3.3 0.00145016 0 0.0014500799999999999 0 0.00145018 3.3 0.0014501 3.3 0.0014502 0 0.0014501199999999998 0 0.00145022 3.3 0.00145014 3.3 0.00145024 0 0.0014501599999999998 0 0.0014502599999999999 3.3 0.00145018 3.3 0.00145028 0 0.0014502 0 0.0014503 3.3 0.00145022 3.3 0.00145032 0 0.00145024 0 0.00145034 3.3 0.0014502599999999999 3.3 0.00145036 0 0.00145028 0 0.00145038 3.3 0.0014502999999999999 3.3 0.0014504 0 0.00145032 0 0.00145042 3.3 0.0014503399999999998 3.3 0.0014504399999999999 0 0.00145036 0 0.00145046 3.3 0.0014503799999999998 3.3 0.0014504799999999999 0 0.0014504 0 0.0014505 3.3 0.00145042 3.3 0.00145052 0 0.0014504399999999999 0 0.00145054 3.3 0.00145046 3.3 0.00145056 0 0.0014504799999999999 0 0.00145058 3.3 0.0014505 3.3 0.0014506 0 0.0014505199999999998 0 0.00145062 3.3 0.00145054 3.3 0.00145064 0 0.0014505599999999998 0 0.0014506599999999999 3.3 0.00145058 3.3 0.00145068 0 0.0014505999999999998 0 0.0014506999999999999 3.3 0.00145062 3.3 0.00145072 0 0.00145064 0 0.00145074 3.3 0.0014506599999999999 3.3 0.00145076 0 0.00145068 0 0.00145078 3.3 0.0014506999999999999 3.3 0.0014508 0 0.00145072 0 0.00145082 3.3 0.0014507399999999998 3.3 0.00145084 0 0.00145076 0 0.00145086 3.3 0.0014507799999999998 3.3 0.0014508799999999999 0 0.0014508 0 0.0014509 3.3 0.00145082 3.3 0.00145092 0 0.00145084 0 0.00145094 3.3 0.00145086 3.3 0.00145096 0 0.0014508799999999999 0 0.00145098 3.3 0.0014509 3.3 0.001451 0 0.0014509199999999999 0 0.00145102 3.3 0.00145094 3.3 0.00145104 0 0.0014509599999999998 0 0.00145106 3.3 0.00145098 3.3 0.00145108 0 0.0014509999999999998 0 0.0014510999999999999 3.3 0.00145102 3.3 0.00145112 0 0.00145104 0 0.00145114 3.3 0.00145106 3.3 0.00145116 0 0.00145108 0 0.00145118 3.3 0.0014510999999999999 3.3 0.0014512 0 0.00145112 0 0.00145122 3.3 0.0014511399999999999 3.3 0.00145124 0 0.00145116 0 0.00145126 3.3 0.0014511799999999998 3.3 0.0014512799999999999 0 0.0014512 0 0.0014513 3.3 0.0014512199999999998 3.3 0.0014513199999999999 0 0.00145124 0 0.00145134 3.3 0.00145126 3.3 0.00145136 0 0.0014512799999999999 0 0.00145138 3.3 0.0014513 3.3 0.0014514 0 0.0014513199999999999 0 0.00145142 3.3 0.00145134 3.3 0.00145144 0 0.0014513599999999998 0 0.00145146 3.3 0.00145138 3.3 0.00145148 0 0.0014513999999999998 0 0.0014514999999999999 3.3 0.00145142 3.3 0.00145152 0 0.00145144 0 0.00145154 3.3 0.00145146 3.3 0.00145156 0 0.00145148 0 0.00145158 3.3 0.0014514999999999999 3.3 0.0014516 0 0.00145152 0 0.00145162 3.3 0.0014515399999999999 3.3 0.00145164 0 0.00145156 0 0.00145166 3.3 0.0014515799999999998 3.3 0.00145168 0 0.0014516 0 0.0014517 3.3 0.0014516199999999998 3.3 0.0014517199999999999 0 0.00145164 0 0.00145174 3.3 0.00145166 3.3 0.00145176 0 0.00145168 0 0.00145178 3.3 0.0014517 3.3 0.0014518 0 0.0014517199999999999 0 0.00145182 3.3 0.00145174 3.3 0.00145184 0 0.0014517599999999999 0 0.00145186 3.3 0.00145178 3.3 0.00145188 0 0.0014517999999999998 0 0.0014519 3.3 0.00145182 3.3 0.00145192 0 0.0014518399999999998 0 0.0014519399999999999 3.3 0.00145186 3.3 0.00145196 0 0.00145188 0 0.00145198 3.3 0.0014519 3.3 0.001452 0 0.00145192 0 0.00145202 3.3 0.0014519399999999999 3.3 0.00145204 0 0.00145196 0 0.00145206 3.3 0.0014519799999999999 3.3 0.00145208 0 0.001452 0 0.0014521 3.3 0.0014520199999999998 3.3 0.0014521199999999999 0 0.00145204 0 0.00145214 3.3 0.0014520599999999998 3.3 0.0014521599999999999 0 0.00145208 0 0.00145218 3.3 0.0014521 3.3 0.0014522 0 0.0014521199999999999 0 0.00145222 3.3 0.00145214 3.3 0.00145224 0 0.0014521599999999999 0 0.00145226 3.3 0.00145218 3.3 0.00145228 0 0.0014521999999999998 0 0.0014523 3.3 0.00145222 3.3 0.00145232 0 0.0014522399999999998 0 0.0014523399999999999 3.3 0.00145226 3.3 0.00145236 0 0.00145228 0 0.00145238 3.3 0.0014523 3.3 0.0014524 0 0.00145232 0 0.00145242 3.3 0.0014523399999999999 3.3 0.00145244 0 0.00145236 0 0.00145246 3.3 0.0014523799999999999 3.3 0.00145248 0 0.0014524 0 0.0014525 3.3 0.0014524199999999998 3.3 0.00145252 0 0.00145244 0 0.00145254 3.3 0.0014524599999999998 3.3 0.0014525599999999999 0 0.00145248 0 0.00145258 3.3 0.0014525 3.3 0.0014526 0 0.00145252 0 0.00145262 3.3 0.00145254 3.3 0.00145264 0 0.0014525599999999999 0 0.00145266 3.3 0.00145258 3.3 0.00145268 0 0.0014525999999999999 0 0.0014527 3.3 0.00145262 3.3 0.00145272 0 0.0014526399999999998 0 0.0014527399999999999 3.3 0.00145266 3.3 0.00145276 0 0.0014526799999999998 0 0.0014527799999999999 3.3 0.0014527 3.3 0.0014528 0 0.00145272 0 0.00145282 3.3 0.0014527399999999999 3.3 0.00145284 0 0.00145276 0 0.00145286 3.3 0.0014527799999999999 3.3 0.00145288 0 0.0014528 0 0.0014529 3.3 0.0014528199999999998 3.3 0.00145292 0 0.00145284 0 0.00145294 3.3 0.0014528599999999998 3.3 0.0014529599999999999 0 0.00145288 0 0.00145298 3.3 0.0014528999999999998 3.3 0.0014529999999999999 0 0.00145292 0 0.00145302 3.3 0.00145294 3.3 0.00145304 0 0.0014529599999999999 0 0.00145306 3.3 0.00145298 3.3 0.00145308 0 0.0014529999999999999 0 0.0014531 3.3 0.00145302 3.3 0.00145312 0 0.0014530399999999998 0 0.00145314 3.3 0.00145306 3.3 0.00145316 0 0.0014530799999999998 0 0.0014531799999999999 3.3 0.0014531 3.3 0.0014532 0 0.00145312 0 0.00145322 3.3 0.00145314 3.3 0.00145324 0 0.00145316 0 0.00145326 3.3 0.0014531799999999999 3.3 0.00145328 0 0.0014532 0 0.0014533 3.3 0.0014532199999999999 3.3 0.00145332 0 0.00145324 0 0.00145334 3.3 0.0014532599999999998 3.3 0.00145336 0 0.00145328 0 0.00145338 3.3 0.0014532999999999998 3.3 0.0014533999999999999 0 0.00145332 0 0.00145342 3.3 0.00145334 3.3 0.00145344 0 0.00145336 0 0.00145346 3.3 0.00145338 3.3 0.00145348 0 0.0014533999999999999 0 0.0014535 3.3 0.00145342 3.3 0.00145352 0 0.0014534399999999999 0 0.00145354 3.3 0.00145346 3.3 0.00145356 0 0.0014534799999999998 0 0.0014535799999999999 3.3 0.0014535 3.3 0.0014536 0 0.0014535199999999998 0 0.0014536199999999999 3.3 0.00145354 3.3 0.00145364 0 0.00145356 0 0.00145366 3.3 0.0014535799999999999 3.3 0.00145368 0 0.0014536 0 0.0014537 3.3 0.0014536199999999999 3.3 0.00145372 0 0.00145364 0 0.00145374 3.3 0.0014536599999999998 3.3 0.00145376 0 0.00145368 0 0.00145378 3.3 0.0014536999999999998 3.3 0.0014537999999999999 0 0.00145372 0 0.00145382 3.3 0.0014537399999999998 3.3 0.0014538399999999999 0 0.00145376 0 0.00145386 3.3 0.00145378 3.3 0.00145388 0 0.0014537999999999999 0 0.0014539 3.3 0.00145382 3.3 0.00145392 0 0.0014538399999999999 0 0.00145394 3.3 0.00145386 3.3 0.00145396 0 0.0014538799999999998 0 0.00145398 3.3 0.0014539 3.3 0.001454 0 0.0014539199999999998 0 0.0014540199999999999 3.3 0.00145394 3.3 0.00145404 0 0.00145396 0 0.00145406 3.3 0.00145398 3.3 0.00145408 0 0.001454 0 0.0014541 3.3 0.0014540199999999999 3.3 0.00145412 0 0.00145404 0 0.00145414 3.3 0.0014540599999999999 3.3 0.00145416 0 0.00145408 0 0.00145418 3.3 0.0014540999999999998 3.3 0.0014542 0 0.00145412 0 0.00145422 3.3 0.0014541399999999998 3.3 0.0014542399999999999 0 0.00145416 0 0.00145426 3.3 0.00145418 3.3 0.00145428 0 0.0014542 0 0.0014543 3.3 0.00145422 3.3 0.00145432 0 0.0014542399999999999 0 0.00145434 3.3 0.00145426 3.3 0.00145436 0 0.0014542799999999999 0 0.00145438 3.3 0.0014543 3.3 0.0014544 0 0.0014543199999999998 0 0.0014544199999999999 3.3 0.00145434 3.3 0.00145444 0 0.0014543599999999998 0 0.0014544599999999999 3.3 0.00145438 3.3 0.00145448 0 0.0014544 0 0.0014545 3.3 0.0014544199999999999 3.3 0.00145452 0 0.00145444 0 0.00145454 3.3 0.0014544599999999999 3.3 0.00145456 0 0.00145448 0 0.00145458 3.3 0.0014544999999999998 3.3 0.0014546 0 0.00145452 0 0.00145462 3.3 0.0014545399999999998 3.3 0.0014546399999999999 0 0.00145456 0 0.00145466 3.3 0.00145458 3.3 0.00145468 0 0.0014546 0 0.0014547 3.3 0.00145462 3.3 0.00145472 0 0.0014546399999999999 0 0.00145474 3.3 0.00145466 3.3 0.00145476 0 0.0014546799999999999 0 0.00145478 3.3 0.0014547 3.3 0.0014548 0 0.0014547199999999998 0 0.00145482 3.3 0.00145474 3.3 0.00145484 0 0.0014547599999999998 0 0.0014548599999999999 3.3 0.00145478 3.3 0.00145488 0 0.0014548 0 0.0014549 3.3 0.00145482 3.3 0.00145492 0 0.00145484 0 0.00145494 3.3 0.0014548599999999999 3.3 0.00145496 0 0.00145488 0 0.00145498 3.3 0.0014548999999999999 3.3 0.001455 0 0.00145492 0 0.00145502 3.3 0.0014549399999999998 3.3 0.00145504 0 0.00145496 0 0.00145506 3.3 0.0014549799999999998 3.3 0.0014550799999999999 0 0.001455 0 0.0014551 3.3 0.00145502 3.3 0.00145512 0 0.00145504 0 0.00145514 3.3 0.00145506 3.3 0.00145516 0 0.0014550799999999999 0 0.00145518 3.3 0.0014551 3.3 0.0014552 0 0.0014551199999999999 0 0.00145522 3.3 0.00145514 3.3 0.00145524 0 0.0014551599999999998 0 0.0014552599999999999 3.3 0.00145518 3.3 0.00145528 0 0.0014551999999999998 0 0.0014552999999999999 3.3 0.00145522 3.3 0.00145532 0 0.00145524 0 0.00145534 3.3 0.0014552599999999999 3.3 0.00145536 0 0.00145528 0 0.00145538 3.3 0.0014552999999999999 3.3 0.0014554 0 0.00145532 0 0.00145542 3.3 0.0014553399999999998 3.3 0.00145544 0 0.00145536 0 0.00145546 3.3 0.0014553799999999998 3.3 0.0014554799999999999 0 0.0014554 0 0.0014555 3.3 0.00145542 3.3 0.00145552 0 0.00145544 0 0.00145554 3.3 0.00145546 3.3 0.00145556 0 0.0014554799999999999 0 0.00145558 3.3 0.0014555 3.3 0.0014556 0 0.0014555199999999999 0 0.00145562 3.3 0.00145554 3.3 0.00145564 0 0.0014555599999999998 0 0.00145566 3.3 0.00145558 3.3 0.00145568 0 0.0014555999999999998 0 0.0014556999999999999 3.3 0.00145562 3.3 0.00145572 0 0.00145564 0 0.00145574 3.3 0.00145566 3.3 0.00145576 0 0.00145568 0 0.00145578 3.3 0.0014556999999999999 3.3 0.0014558 0 0.00145572 0 0.00145582 3.3 0.0014557399999999999 3.3 0.00145584 0 0.00145576 0 0.00145586 3.3 0.0014557799999999998 3.3 0.0014558799999999999 0 0.0014558 0 0.0014559 3.3 0.0014558199999999998 3.3 0.0014559199999999999 0 0.00145584 0 0.00145594 3.3 0.00145586 3.3 0.00145596 0 0.0014558799999999999 0 0.00145598 3.3 0.0014559 3.3 0.001456 0 0.0014559199999999999 0 0.00145602 3.3 0.00145594 3.3 0.00145604 0 0.0014559599999999998 0 0.00145606 3.3 0.00145598 3.3 0.00145608 0 0.0014559999999999998 0 0.0014560999999999999 3.3 0.00145602 3.3 0.00145612 0 0.0014560399999999998 0 0.0014561399999999999 3.3 0.00145606 3.3 0.00145616 0 0.00145608 0 0.00145618 3.3 0.0014560999999999999 3.3 0.0014562 0 0.00145612 0 0.00145622 3.3 0.0014561399999999999 3.3 0.00145624 0 0.00145616 0 0.00145626 3.3 0.0014561799999999998 3.3 0.00145628 0 0.0014562 0 0.0014563 3.3 0.0014562199999999998 3.3 0.0014563199999999999 0 0.00145624 0 0.00145634 3.3 0.00145626 3.3 0.00145636 0 0.00145628 0 0.00145638 3.3 0.0014563 3.3 0.0014564 0 0.0014563199999999999 0 0.00145642 3.3 0.00145634 3.3 0.00145644 0 0.0014563599999999999 0 0.00145646 3.3 0.00145638 3.3 0.00145648 0 0.0014563999999999998 0 0.0014565 3.3 0.00145642 3.3 0.00145652 0 0.0014564399999999998 0 0.0014565399999999999 3.3 0.00145646 3.3 0.00145656 0 0.00145648 0 0.00145658 3.3 0.0014565 3.3 0.0014566 0 0.00145652 0 0.00145662 3.3 0.0014565399999999999 3.3 0.00145664 0 0.00145656 0 0.00145666 3.3 0.0014565799999999999 3.3 0.00145668 0 0.0014566 0 0.0014567 3.3 0.0014566199999999998 3.3 0.0014567199999999999 0 0.00145664 0 0.00145674 3.3 0.0014566599999999998 3.3 0.0014567599999999999 0 0.00145668 0 0.00145678 3.3 0.0014567 3.3 0.0014568 0 0.0014567199999999999 0 0.00145682 3.3 0.00145674 3.3 0.00145684 0 0.0014567599999999999 0 0.00145686 3.3 0.00145678 3.3 0.00145688 0 0.0014567999999999998 0 0.0014569 3.3 0.00145682 3.3 0.00145692 0 0.0014568399999999998 0 0.0014569399999999999 3.3 0.00145686 3.3 0.00145696 0 0.0014568799999999998 0 0.0014569799999999999 3.3 0.0014569 3.3 0.001457 0 0.00145692 0 0.00145702 3.3 0.0014569399999999999 3.3 0.00145704 0 0.00145696 0 0.00145706 3.3 0.0014569799999999999 3.3 0.00145708 0 0.001457 0 0.0014571 3.3 0.0014570199999999998 3.3 0.00145712 0 0.00145704 0 0.00145714 3.3 0.0014570599999999998 3.3 0.0014571599999999999 0 0.00145708 0 0.00145718 3.3 0.0014571 3.3 0.0014572 0 0.00145712 0 0.00145722 3.3 0.00145714 3.3 0.00145724 0 0.0014571599999999999 0 0.00145726 3.3 0.00145718 3.3 0.00145728 0 0.0014571999999999999 0 0.0014573 3.3 0.00145722 3.3 0.00145732 0 0.0014572399999999998 0 0.00145734 3.3 0.00145726 3.3 0.00145736 0 0.0014572799999999998 0 0.0014573799999999999 3.3 0.0014573 3.3 0.0014574 0 0.00145732 0 0.00145742 3.3 0.00145734 3.3 0.00145744 0 0.00145736 0 0.00145746 3.3 0.0014573799999999999 3.3 0.00145748 0 0.0014574 0 0.0014575 3.3 0.0014574199999999999 3.3 0.00145752 0 0.00145744 0 0.00145754 3.3 0.0014574599999999998 3.3 0.0014575599999999999 0 0.00145748 0 0.00145758 3.3 0.0014574999999999998 3.3 0.0014575999999999999 0 0.00145752 0 0.00145762 3.3 0.00145754 3.3 0.00145764 0 0.0014575599999999999 0 0.00145766 3.3 0.00145758 3.3 0.00145768 0 0.0014575999999999999 0 0.0014577 3.3 0.00145762 3.3 0.00145772 0 0.0014576399999999998 0 0.00145774 3.3 0.00145766 3.3 0.00145776 0 0.0014576799999999998 0 0.0014577799999999999 3.3 0.0014577 3.3 0.0014578 0 0.0014577199999999998 0 0.0014578199999999999 3.3 0.00145774 3.3 0.00145784 0 0.00145776 0 0.00145786 3.3 0.0014577799999999999 3.3 0.00145788 0 0.0014578 0 0.0014579 3.3 0.0014578199999999999 3.3 0.00145792 0 0.00145784 0 0.00145794 3.3 0.0014578599999999998 3.3 0.00145796 0 0.00145788 0 0.00145798 3.3 0.0014578999999999998 3.3 0.0014579999999999999 0 0.00145792 0 0.00145802 3.3 0.00145794 3.3 0.00145804 0 0.00145796 0 0.00145806 3.3 0.00145798 3.3 0.00145808 0 0.0014579999999999999 0 0.0014581 3.3 0.00145802 3.3 0.00145812 0 0.0014580399999999999 0 0.00145814 3.3 0.00145806 3.3 0.00145816 0 0.0014580799999999998 0 0.00145818 3.3 0.0014581 3.3 0.0014582 0 0.0014581199999999998 0 0.0014582199999999999 3.3 0.00145814 3.3 0.00145824 0 0.00145816 0 0.00145826 3.3 0.00145818 3.3 0.00145828 0 0.0014582 0 0.0014583 3.3 0.0014582199999999999 3.3 0.00145832 0 0.00145824 0 0.00145834 3.3 0.0014582599999999999 3.3 0.00145836 0 0.00145828 0 0.00145838 3.3 0.0014582999999999998 3.3 0.0014583999999999999 0 0.00145832 0 0.00145842 3.3 0.0014583399999999998 3.3 0.0014584399999999999 0 0.00145836 0 0.00145846 3.3 0.00145838 3.3 0.00145848 0 0.0014583999999999999 0 0.0014585 3.3 0.00145842 3.3 0.00145852 0 0.0014584399999999999 0 0.00145854 3.3 0.00145846 3.3 0.00145856 0 0.0014584799999999998 0 0.00145858 3.3 0.0014585 3.3 0.0014586 0 0.0014585199999999998 0 0.0014586199999999999 3.3 0.00145854 3.3 0.00145864 0 0.00145856 0 0.00145866 3.3 0.00145858 3.3 0.00145868 0 0.0014586 0 0.0014587 3.3 0.0014586199999999999 3.3 0.00145872 0 0.00145864 0 0.00145874 3.3 0.0014586599999999999 3.3 0.00145876 0 0.00145868 0 0.00145878 3.3 0.0014586999999999998 3.3 0.0014588 0 0.00145872 0 0.00145882 3.3 0.0014587399999999998 3.3 0.0014588399999999999 0 0.00145876 0 0.00145886 3.3 0.00145878 3.3 0.00145888 0 0.0014588 0 0.0014589 3.3 0.00145882 3.3 0.00145892 0 0.0014588399999999999 0 0.00145894 3.3 0.00145886 3.3 0.00145896 0 0.0014588799999999999 0 0.00145898 3.3 0.0014589 3.3 0.001459 0 0.0014589199999999998 0 0.00145902 3.3 0.00145894 3.3 0.00145904 0 0.0014589599999999998 0 0.0014590599999999999 3.3 0.00145898 3.3 0.00145908 0 0.001459 0 0.0014591 3.3 0.00145902 3.3 0.00145912 0 0.00145904 0 0.00145914 3.3 0.0014590599999999999 3.3 0.00145916 0 0.00145908 0 0.00145918 3.3 0.0014590999999999999 3.3 0.0014592 0 0.00145912 0 0.00145922 3.3 0.0014591399999999998 3.3 0.0014592399999999999 0 0.00145916 0 0.00145926 3.3 0.0014591799999999998 3.3 0.0014592799999999999 0 0.0014592 0 0.0014593 3.3 0.00145922 3.3 0.00145932 0 0.0014592399999999999 0 0.00145934 3.3 0.00145926 3.3 0.00145936 0 0.0014592799999999999 0 0.00145938 3.3 0.0014593 3.3 0.0014594 0 0.0014593199999999998 0 0.00145942 3.3 0.00145934 3.3 0.00145944 0 0.0014593599999999998 0 0.0014594599999999999 3.3 0.00145938 3.3 0.00145948 0 0.0014594 0 0.0014595 3.3 0.00145942 3.3 0.00145952 0 0.00145944 0 0.00145954 3.3 0.0014594599999999999 3.3 0.00145956 0 0.00145948 0 0.00145958 3.3 0.0014594999999999999 3.3 0.0014596 0 0.00145952 0 0.00145962 3.3 0.0014595399999999998 3.3 0.00145964 0 0.00145956 0 0.00145966 3.3 0.0014595799999999998 3.3 0.0014596799999999999 0 0.0014596 0 0.0014597 3.3 0.00145962 3.3 0.00145972 0 0.00145964 0 0.00145974 3.3 0.00145966 3.3 0.00145976 0 0.0014596799999999999 0 0.00145978 3.3 0.0014597 3.3 0.0014598 0 0.0014597199999999999 0 0.00145982 3.3 0.00145974 3.3 0.00145984 0 0.0014597599999999998 0 0.0014598599999999999 3.3 0.00145978 3.3 0.00145988 0 0.0014597999999999998 0 0.0014598999999999999 3.3 0.00145982 3.3 0.00145992 0 0.00145984 0 0.00145994 3.3 0.0014598599999999999 3.3 0.00145996 0 0.00145988 0 0.00145998 3.3 0.0014598999999999999 3.3 0.00146 0 0.00145992 0 0.00146002 3.3 0.0014599399999999998 3.3 0.00146004 0 0.00145996 0 0.00146006 3.3 0.0014599799999999998 3.3 0.0014600799999999999 0 0.00146 0 0.0014601 3.3 0.0014600199999999998 3.3 0.0014601199999999999 0 0.00146004 0 0.00146014 3.3 0.00146006 3.3 0.00146016 0 0.0014600799999999999 0 0.00146018 3.3 0.0014601 3.3 0.0014602 0 0.0014601199999999999 0 0.00146022 3.3 0.00146014 3.3 0.00146024 0 0.0014601599999999998 0 0.00146026 3.3 0.00146018 3.3 0.00146028 0 0.0014601999999999998 0 0.0014602999999999999 3.3 0.00146022 3.3 0.00146032 0 0.00146024 0 0.00146034 3.3 0.00146026 3.3 0.00146036 0 0.00146028 0 0.00146038 3.3 0.0014602999999999999 3.3 0.0014604 0 0.00146032 0 0.00146042 3.3 0.0014603399999999999 3.3 0.00146044 0 0.00146036 0 0.00146046 3.3 0.0014603799999999998 3.3 0.00146048 0 0.0014604 0 0.0014605 3.3 0.0014604199999999998 3.3 0.0014605199999999999 0 0.00146044 0 0.00146054 3.3 0.00146046 3.3 0.00146056 0 0.00146048 0 0.00146058 3.3 0.0014605 3.3 0.0014606 0 0.0014605199999999999 0 0.00146062 3.3 0.00146054 3.3 0.00146064 0 0.0014605599999999999 0 0.00146066 3.3 0.00146058 3.3 0.00146068 0 0.0014605999999999998 0 0.0014606999999999999 3.3 0.00146062 3.3 0.00146072 0 0.0014606399999999998 0 0.0014607399999999999 3.3 0.00146066 3.3 0.00146076 0 0.00146068 0 0.00146078 3.3 0.0014606999999999999 3.3 0.0014608 0 0.00146072 0 0.00146082 3.3 0.0014607399999999999 3.3 0.00146084 0 0.00146076 0 0.00146086 3.3 0.0014607799999999998 3.3 0.00146088 0 0.0014608 0 0.0014609 3.3 0.0014608199999999998 3.3 0.0014609199999999999 0 0.00146084 0 0.00146094 3.3 0.0014608599999999998 3.3 0.0014609599999999999 0 0.00146088 0 0.00146098 3.3 0.0014609 3.3 0.001461 0 0.0014609199999999999 0 0.00146102 3.3 0.00146094 3.3 0.00146104 0 0.0014609599999999999 0 0.00146106 3.3 0.00146098 3.3 0.00146108 0 0.0014609999999999998 0 0.0014611 3.3 0.00146102 3.3 0.00146112 0 0.0014610399999999998 0 0.0014611399999999999 3.3 0.00146106 3.3 0.00146116 0 0.00146108 0 0.00146118 3.3 0.0014611 3.3 0.0014612 0 0.00146112 0 0.00146122 3.3 0.0014611399999999999 3.3 0.00146124 0 0.00146116 0 0.00146126 3.3 0.0014611799999999999 3.3 0.00146128 0 0.0014612 0 0.0014613 3.3 0.0014612199999999998 3.3 0.00146132 0 0.00146124 0 0.00146134 3.3 0.0014612599999999998 3.3 0.0014613599999999999 0 0.00146128 0 0.00146138 3.3 0.0014613 3.3 0.0014614 0 0.00146132 0 0.00146142 3.3 0.00146134 3.3 0.00146144 0 0.0014613599999999999 0 0.00146146 3.3 0.00146138 3.3 0.00146148 0 0.0014613999999999999 0 0.0014615 3.3 0.00146142 3.3 0.00146152 0 0.0014614399999999998 0 0.0014615399999999999 3.3 0.00146146 3.3 0.00146156 0 0.0014614799999999998 0 0.0014615799999999999 3.3 0.0014615 3.3 0.0014616 0 0.00146152 0 0.00146162 3.3 0.0014615399999999999 3.3 0.00146164 0 0.00146156 0 0.00146166 3.3 0.0014615799999999999 3.3 0.00146168 0 0.0014616 0 0.0014617 3.3 0.0014616199999999998 3.3 0.00146172 0 0.00146164 0 0.00146174 3.3 0.0014616599999999998 3.3 0.0014617599999999999 0 0.00146168 0 0.00146178 3.3 0.0014617 3.3 0.0014618 0 0.00146172 0 0.00146182 3.3 0.00146174 3.3 0.00146184 0 0.0014617599999999999 0 0.00146186 3.3 0.00146178 3.3 0.00146188 0 0.0014617999999999999 0 0.0014619 3.3 0.00146182 3.3 0.00146192 0 0.0014618399999999998 0 0.00146194 3.3 0.00146186 3.3 0.00146196 0 0.0014618799999999998 0 0.0014619799999999999 3.3 0.0014619 3.3 0.001462 0 0.00146192 0 0.00146202 3.3 0.00146194 3.3 0.00146204 0 0.00146196 0 0.00146206 3.3 0.0014619799999999999 3.3 0.00146208 0 0.001462 0 0.0014621 3.3 0.0014620199999999999 3.3 0.00146212 0 0.00146204 0 0.00146214 3.3 0.0014620599999999998 3.3 0.00146216 0 0.00146208 0 0.00146218 3.3 0.0014620999999999998 3.3 0.0014621999999999999 0 0.00146212 0 0.00146222 3.3 0.00146214 3.3 0.00146224 0 0.00146216 0 0.00146226 3.3 0.00146218 3.3 0.00146228 0 0.0014621999999999999 0 0.0014623 3.3 0.00146222 3.3 0.00146232 0 0.0014622399999999999 0 0.00146234 3.3 0.00146226 3.3 0.00146236 0 0.0014622799999999998 0 0.0014623799999999999 3.3 0.0014623 3.3 0.0014624 0 0.0014623199999999998 0 0.0014624199999999999 3.3 0.00146234 3.3 0.00146244 0 0.00146236 0 0.00146246 3.3 0.0014623799999999999 3.3 0.00146248 0 0.0014624 0 0.0014625 3.3 0.0014624199999999999 3.3 0.00146252 0 0.00146244 0 0.00146254 3.3 0.0014624599999999998 3.3 0.00146256 0 0.00146248 0 0.00146258 3.3 0.0014624999999999998 3.3 0.0014625999999999999 0 0.00146252 0 0.00146262 3.3 0.00146254 3.3 0.00146264 0 0.00146256 0 0.00146266 3.3 0.00146258 3.3 0.00146268 0 0.0014625999999999999 0 0.0014627 3.3 0.00146262 3.3 0.00146272 0 0.0014626399999999999 0 0.00146274 3.3 0.00146266 3.3 0.00146276 0 0.0014626799999999998 0 0.00146278 3.3 0.0014627 3.3 0.0014628 0 0.0014627199999999998 0 0.0014628199999999999 3.3 0.00146274 3.3 0.00146284 0 0.00146276 0 0.00146286 3.3 0.00146278 3.3 0.00146288 0 0.0014628 0 0.0014629 3.3 0.0014628199999999999 3.3 0.00146292 0 0.00146284 0 0.00146294 3.3 0.0014628599999999999 3.3 0.00146296 0 0.00146288 0 0.00146298 3.3 0.0014628999999999998 3.3 0.0014629999999999999 0 0.00146292 0 0.00146302 3.3 0.0014629399999999998 3.3 0.0014630399999999999 0 0.00146296 0 0.00146306 3.3 0.00146298 3.3 0.00146308 0 0.0014629999999999999 0 0.0014631 3.3 0.00146302 3.3 0.00146312 0 0.0014630399999999999 0 0.00146314 3.3 0.00146306 3.3 0.00146316 0 0.0014630799999999998 0 0.00146318 3.3 0.0014631 3.3 0.0014632 0 0.0014631199999999998 0 0.0014632199999999999 3.3 0.00146314 3.3 0.00146324 0 0.0014631599999999998 0 0.0014632599999999999 3.3 0.00146318 3.3 0.00146328 0 0.0014632 0 0.0014633 3.3 0.0014632199999999999 3.3 0.00146332 0 0.00146324 0 0.00146334 3.3 0.0014632599999999999 3.3 0.00146336 0 0.00146328 0 0.00146338 3.3 0.0014632999999999998 3.3 0.0014634 0 0.00146332 0 0.00146342 3.3 0.0014633399999999998 3.3 0.0014634399999999999 0 0.00146336 0 0.00146346 3.3 0.00146338 3.3 0.00146348 0 0.0014634 0 0.0014635 3.3 0.00146342 3.3 0.00146352 0 0.0014634399999999999 0 0.00146354 3.3 0.00146346 3.3 0.00146356 0 0.0014634799999999999 0 0.00146358 3.3 0.0014635 3.3 0.0014636 0 0.0014635199999999998 0 0.00146362 3.3 0.00146354 3.3 0.00146364 0 0.0014635599999999998 0 0.0014636599999999999 3.3 0.00146358 3.3 0.00146368 0 0.0014636 0 0.0014637 3.3 0.00146362 3.3 0.00146372 0 0.00146364 0 0.00146374 3.3 0.0014636599999999999 3.3 0.00146376 0 0.00146368 0 0.00146378 3.3 0.0014636999999999999 3.3 0.0014638 0 0.00146372 0 0.00146382 3.3 0.0014637399999999998 3.3 0.0014638399999999999 0 0.00146376 0 0.00146386 3.3 0.0014637799999999998 3.3 0.0014638799999999999 0 0.0014638 0 0.0014639 3.3 0.00146382 3.3 0.00146392 0 0.0014638399999999999 0 0.00146394 3.3 0.00146386 3.3 0.00146396 0 0.0014638799999999999 0 0.00146398 3.3 0.0014639 3.3 0.001464 0 0.0014639199999999998 0 0.00146402 3.3 0.00146394 3.3 0.00146404 0 0.0014639599999999998 0 0.0014640599999999999 3.3 0.00146398 3.3 0.00146408 0 0.0014639999999999998 0 0.0014640999999999999 3.3 0.00146402 3.3 0.00146412 0 0.00146404 0 0.00146414 3.3 0.0014640599999999999 3.3 0.00146416 0 0.00146408 0 0.00146418 3.3 0.0014640999999999999 3.3 0.0014642 0 0.00146412 0 0.00146422 3.3 0.0014641399999999998 3.3 0.00146424 0 0.00146416 0 0.00146426 3.3 0.0014641799999999998 3.3 0.0014642799999999999 0 0.0014642 0 0.0014643 3.3 0.00146422 3.3 0.00146432 0 0.00146424 0 0.00146434 3.3 0.00146426 3.3 0.00146436 0 0.0014642799999999999 0 0.00146438 3.3 0.0014643 3.3 0.0014644 0 0.0014643199999999999 0 0.00146442 3.3 0.00146434 3.3 0.00146444 0 0.0014643599999999998 0 0.00146446 3.3 0.00146438 3.3 0.00146448 0 0.0014643999999999998 0 0.0014644999999999999 3.3 0.00146442 3.3 0.00146452 0 0.00146444 0 0.00146454 3.3 0.00146446 3.3 0.00146456 0 0.00146448 0 0.00146458 3.3 0.0014644999999999999 3.3 0.0014646 0 0.00146452 0 0.00146462 3.3 0.0014645399999999999 3.3 0.00146464 0 0.00146456 0 0.00146466 3.3 0.0014645799999999998 3.3 0.0014646799999999999 0 0.0014646 0 0.0014647 3.3 0.0014646199999999998 3.3 0.0014647199999999999 0 0.00146464 0 0.00146474 3.3 0.00146466 3.3 0.00146476 0 0.0014646799999999999 0 0.00146478 3.3 0.0014647 3.3 0.0014648 0 0.0014647199999999999 0 0.00146482 3.3 0.00146474 3.3 0.00146484 0 0.0014647599999999998 0 0.00146486 3.3 0.00146478 3.3 0.00146488 0 0.0014647999999999998 0 0.0014648999999999999 3.3 0.00146482 3.3 0.00146492 0 0.00146484 0 0.00146494 3.3 0.00146486 3.3 0.00146496 0 0.00146488 0 0.00146498 3.3 0.0014648999999999999 3.3 0.001465 0 0.00146492 0 0.00146502 3.3 0.0014649399999999999 3.3 0.00146504 0 0.00146496 0 0.00146506 3.3 0.0014649799999999998 3.3 0.00146508 0 0.001465 0 0.0014651 3.3 0.0014650199999999998 3.3 0.0014651199999999999 0 0.00146504 0 0.00146514 3.3 0.00146506 3.3 0.00146516 0 0.00146508 0 0.00146518 3.3 0.0014651 3.3 0.0014652 0 0.0014651199999999999 0 0.00146522 3.3 0.00146514 3.3 0.00146524 0 0.0014651599999999999 0 0.00146526 3.3 0.00146518 3.3 0.00146528 0 0.0014651999999999998 0 0.0014653 3.3 0.00146522 3.3 0.00146532 0 0.0014652399999999998 0 0.0014653399999999999 3.3 0.00146526 3.3 0.00146536 0 0.00146528 0 0.00146538 3.3 0.0014653 3.3 0.0014654 0 0.00146532 0 0.00146542 3.3 0.0014653399999999999 3.3 0.00146544 0 0.00146536 0 0.00146546 3.3 0.0014653799999999999 3.3 0.00146548 0 0.0014654 0 0.0014655 3.3 0.0014654199999999998 3.3 0.0014655199999999999 0 0.00146544 0 0.00146554 3.3 0.0014654599999999998 3.3 0.0014655599999999999 0 0.00146548 0 0.00146558 3.3 0.0014655 3.3 0.0014656 0 0.0014655199999999999 0 0.00146562 3.3 0.00146554 3.3 0.00146564 0 0.0014655599999999999 0 0.00146566 3.3 0.00146558 3.3 0.00146568 0 0.0014655999999999998 0 0.0014657 3.3 0.00146562 3.3 0.00146572 0 0.0014656399999999998 0 0.0014657399999999999 3.3 0.00146566 3.3 0.00146576 0 0.00146568 0 0.00146578 3.3 0.0014657 3.3 0.0014658 0 0.00146572 0 0.00146582 3.3 0.0014657399999999999 3.3 0.00146584 0 0.00146576 0 0.00146586 3.3 0.0014657799999999999 3.3 0.00146588 0 0.0014658 0 0.0014659 3.3 0.0014658199999999998 3.3 0.00146592 0 0.00146584 0 0.00146594 3.3 0.0014658599999999998 3.3 0.0014659599999999999 0 0.00146588 0 0.00146598 3.3 0.0014659 3.3 0.001466 0 0.00146592 0 0.00146602 3.3 0.00146594 3.3 0.00146604 0 0.0014659599999999999 0 0.00146606 3.3 0.00146598 3.3 0.00146608 0 0.0014659999999999999 0 0.0014661 3.3 0.00146602 3.3 0.00146612 0 0.0014660399999999998 0 0.0014661399999999999 3.3 0.00146606 3.3 0.00146616 0 0.0014660799999999998 0 0.0014661799999999999 3.3 0.0014661 3.3 0.0014662 0 0.00146612 0 0.00146622 3.3 0.0014661399999999999 3.3 0.00146624 0 0.00146616 0 0.00146626 3.3 0.0014661799999999999 3.3 0.00146628 0 0.0014662 0 0.0014663 3.3 0.0014662199999999998 3.3 0.00146632 0 0.00146624 0 0.00146634 3.3 0.0014662599999999998 3.3 0.0014663599999999999 0 0.00146628 0 0.00146638 3.3 0.0014662999999999998 3.3 0.0014663999999999999 0 0.00146632 0 0.00146642 3.3 0.00146634 3.3 0.00146644 0 0.0014663599999999999 0 0.00146646 3.3 0.00146638 3.3 0.00146648 0 0.0014663999999999999 0 0.0014665 3.3 0.00146642 3.3 0.00146652 0 0.0014664399999999998 0 0.00146654 3.3 0.00146646 3.3 0.00146656 0 0.0014664799999999998 0 0.0014665799999999999 3.3 0.0014665 3.3 0.0014666 0 0.00146652 0 0.00146662 3.3 0.00146654 3.3 0.00146664 0 0.00146656 0 0.00146666 3.3 0.0014665799999999999 3.3 0.00146668 0 0.0014666 0 0.0014667 3.3 0.0014666199999999999 3.3 0.00146672 0 0.00146664 0 0.00146674 3.3 0.0014666599999999998 3.3 0.00146676 0 0.00146668 0 0.00146678 3.3 0.0014666999999999998 3.3 0.0014667999999999999 0 0.00146672 0 0.00146682 3.3 0.00146674 3.3 0.00146684 0 0.00146676 0 0.00146686 3.3 0.00146678 3.3 0.00146688 0 0.0014667999999999999 0 0.0014669 3.3 0.00146682 3.3 0.00146692 0 0.0014668399999999999 0 0.00146694 3.3 0.00146686 3.3 0.00146696 0 0.0014668799999999998 0 0.0014669799999999999 3.3 0.0014669 3.3 0.001467 0 0.0014669199999999998 0 0.0014670199999999999 3.3 0.00146694 3.3 0.00146704 0 0.00146696 0 0.00146706 3.3 0.0014669799999999999 3.3 0.00146708 0 0.001467 0 0.0014671 3.3 0.0014670199999999999 3.3 0.00146712 0 0.00146704 0 0.00146714 3.3 0.0014670599999999998 3.3 0.00146716 0 0.00146708 0 0.00146718 3.3 0.0014670999999999998 3.3 0.0014671999999999999 0 0.00146712 0 0.00146722 3.3 0.0014671399999999998 3.3 0.0014672399999999999 0 0.00146716 0 0.00146726 3.3 0.00146718 3.3 0.00146728 0 0.0014671999999999999 0 0.0014673 3.3 0.00146722 3.3 0.00146732 0 0.0014672399999999999 0 0.00146734 3.3 0.00146726 3.3 0.00146736 0 0.0014672799999999998 0 0.00146738 3.3 0.0014673 3.3 0.0014674 0 0.0014673199999999998 0 0.0014674199999999999 3.3 0.00146734 3.3 0.00146744 0 0.00146736 0 0.00146746 3.3 0.00146738 3.3 0.00146748 0 0.0014674 0 0.0014675 3.3 0.0014674199999999999 3.3 0.00146752 0 0.00146744 0 0.00146754 3.3 0.0014674599999999999 3.3 0.00146756 0 0.00146748 0 0.00146758 3.3 0.0014674999999999998 3.3 0.0014676 0 0.00146752 0 0.00146762 3.3 0.0014675399999999998 3.3 0.0014676399999999999 0 0.00146756 0 0.00146766 3.3 0.00146758 3.3 0.00146768 0 0.0014676 0 0.0014677 3.3 0.00146762 3.3 0.00146772 0 0.0014676399999999999 0 0.00146774 3.3 0.00146766 3.3 0.00146776 0 0.0014676799999999999 0 0.00146778 3.3 0.0014677 3.3 0.0014678 0 0.0014677199999999998 0 0.0014678199999999999 3.3 0.00146774 3.3 0.00146784 0 0.0014677599999999998 0 0.0014678599999999999 3.3 0.00146778 3.3 0.00146788 0 0.0014678 0 0.0014679 3.3 0.0014678199999999999 3.3 0.00146792 0 0.00146784 0 0.00146794 3.3 0.0014678599999999999 3.3 0.00146796 0 0.00146788 0 0.00146798 3.3 0.0014678999999999998 3.3 0.001468 0 0.00146792 0 0.00146802 3.3 0.0014679399999999998 3.3 0.0014680399999999999 0 0.00146796 0 0.00146806 3.3 0.0014679799999999998 3.3 0.0014680799999999999 0 0.001468 0 0.0014681 3.3 0.00146802 3.3 0.00146812 0 0.0014680399999999999 0 0.00146814 3.3 0.00146806 3.3 0.00146816 0 0.0014680799999999999 0 0.00146818 3.3 0.0014681 3.3 0.0014682 0 0.0014681199999999998 0 0.00146822 3.3 0.00146814 3.3 0.00146824 0 0.0014681599999999998 0 0.0014682599999999999 3.3 0.00146818 3.3 0.00146828 0 0.0014682 0 0.0014683 3.3 0.00146822 3.3 0.00146832 0 0.00146824 0 0.00146834 3.3 0.0014682599999999999 3.3 0.00146836 0 0.00146828 0 0.00146838 3.3 0.0014682999999999999 3.3 0.0014684 0 0.00146832 0 0.00146842 3.3 0.0014683399999999998 3.3 0.00146844 0 0.00146836 0 0.00146846 3.3 0.0014683799999999998 3.3 0.0014684799999999999 0 0.0014684 0 0.0014685 3.3 0.00146842 3.3 0.00146852 0 0.00146844 0 0.00146854 3.3 0.00146846 3.3 0.00146856 0 0.0014684799999999999 0 0.00146858 3.3 0.0014685 3.3 0.0014686 0 0.0014685199999999999 0 0.00146862 3.3 0.00146854 3.3 0.00146864 0 0.0014685599999999998 0 0.0014686599999999999 3.3 0.00146858 3.3 0.00146868 0 0.0014685999999999998 0 0.0014686999999999999 3.3 0.00146862 3.3 0.00146872 0 0.00146864 0 0.00146874 3.3 0.0014686599999999999 3.3 0.00146876 0 0.00146868 0 0.00146878 3.3 0.0014686999999999999 3.3 0.0014688 0 0.00146872 0 0.00146882 3.3 0.0014687399999999998 3.3 0.00146884 0 0.00146876 0 0.00146886 3.3 0.0014687799999999998 3.3 0.0014688799999999999 0 0.0014688 0 0.0014689 3.3 0.00146882 3.3 0.00146892 0 0.00146884 0 0.00146894 3.3 0.00146886 3.3 0.00146896 0 0.0014688799999999999 0 0.00146898 3.3 0.0014689 3.3 0.001469 0 0.0014689199999999999 0 0.00146902 3.3 0.00146894 3.3 0.00146904 0 0.0014689599999999998 0 0.00146906 3.3 0.00146898 3.3 0.00146908 0 0.0014689999999999998 0 0.0014690999999999999 3.3 0.00146902 3.3 0.00146912 0 0.00146904 0 0.00146914 3.3 0.00146906 3.3 0.00146916 0 0.00146908 0 0.00146918 3.3 0.0014690999999999999 3.3 0.0014692 0 0.00146912 0 0.00146922 3.3 0.0014691399999999999 3.3 0.00146924 0 0.00146916 0 0.00146926 3.3 0.0014691799999999998 3.3 0.00146928 0 0.0014692 0 0.0014693 3.3 0.0014692199999999998 3.3 0.0014693199999999999 0 0.00146924 0 0.00146934 3.3 0.00146926 3.3 0.00146936 0 0.00146928 0 0.00146938 3.3 0.0014693 3.3 0.0014694 0 0.0014693199999999999 0 0.00146942 3.3 0.00146934 3.3 0.00146944 0 0.0014693599999999999 0 0.00146946 3.3 0.00146938 3.3 0.00146948 0 0.0014693999999999998 0 0.0014694999999999999 3.3 0.00146942 3.3 0.00146952 0 0.0014694399999999998 0 0.0014695399999999999 3.3 0.00146946 3.3 0.00146956 0 0.00146948 0 0.00146958 3.3 0.0014694999999999999 3.3 0.0014696 0 0.00146952 0 0.00146962 3.3 0.0014695399999999999 3.3 0.00146964 0 0.00146956 0 0.00146966 3.3 0.0014695799999999998 3.3 0.00146968 0 0.0014696 0 0.0014697 3.3 0.0014696199999999998 3.3 0.0014697199999999999 0 0.00146964 0 0.00146974 3.3 0.00146966 3.3 0.00146976 0 0.00146968 0 0.00146978 3.3 0.0014697 3.3 0.0014698 0 0.0014697199999999999 0 0.00146982 3.3 0.00146974 3.3 0.00146984 0 0.0014697599999999999 0 0.00146986 3.3 0.00146978 3.3 0.00146988 0 0.0014697999999999998 0 0.0014699 3.3 0.00146982 3.3 0.00146992 0 0.0014698399999999998 0 0.0014699399999999999 3.3 0.00146986 3.3 0.00146996 0 0.00146988 0 0.00146998 3.3 0.0014699 3.3 0.00147 0 0.00146992 0 0.00147002 3.3 0.0014699399999999999 3.3 0.00147004 0 0.00146996 0 0.00147006 3.3 0.0014699799999999999 3.3 0.00147008 0 0.00147 0 0.0014701 3.3 0.0014700199999999998 3.3 0.0014701199999999999 0 0.00147004 0 0.00147014 3.3 0.0014700599999999998 3.3 0.0014701599999999999 0 0.00147008 0 0.00147018 3.3 0.0014701 3.3 0.0014702 0 0.0014701199999999999 0 0.00147022 3.3 0.00147014 3.3 0.00147024 0 0.0014701599999999999 0 0.00147026 3.3 0.00147018 3.3 0.00147028 0 0.0014701999999999998 0 0.0014703 3.3 0.00147022 3.3 0.00147032 0 0.0014702399999999998 0 0.0014703399999999999 3.3 0.00147026 3.3 0.00147036 0 0.0014702799999999998 0 0.0014703799999999999 3.3 0.0014703 3.3 0.0014704 0 0.00147032 0 0.00147042 3.3 0.0014703399999999999 3.3 0.00147044 0 0.00147036 0 0.00147046 3.3 0.0014703799999999999 3.3 0.00147048 0 0.0014704 0 0.0014705 3.3 0.0014704199999999998 3.3 0.00147052 0 0.00147044 0 0.00147054 3.3 0.0014704599999999998 3.3 0.0014705599999999999 0 0.00147048 0 0.00147058 3.3 0.0014705 3.3 0.0014706 0 0.00147052 0 0.00147062 3.3 0.00147054 3.3 0.00147064 0 0.0014705599999999999 0 0.00147066 3.3 0.00147058 3.3 0.00147068 0 0.0014705999999999999 0 0.0014707 3.3 0.00147062 3.3 0.00147072 0 0.0014706399999999998 0 0.00147074 3.3 0.00147066 3.3 0.00147076 0 0.0014706799999999998 0 0.0014707799999999999 3.3 0.0014707 3.3 0.0014708 0 0.00147072 0 0.00147082 3.3 0.00147074 3.3 0.00147084 0 0.00147076 0 0.00147086 3.3 0.0014707799999999999 3.3 0.00147088 0 0.0014708 0 0.0014709 3.3 0.0014708199999999999 3.3 0.00147092 0 0.00147084 0 0.00147094 3.3 0.0014708599999999998 3.3 0.0014709599999999999 0 0.00147088 0 0.00147098 3.3 0.0014708999999999998 3.3 0.0014709999999999999 0 0.00147092 0 0.00147102 3.3 0.00147094 3.3 0.00147104 0 0.0014709599999999999 0 0.00147106 3.3 0.00147098 3.3 0.00147108 0 0.0014709999999999999 0 0.0014711 3.3 0.00147102 3.3 0.00147112 0 0.0014710399999999998 0 0.00147114 3.3 0.00147106 3.3 0.00147116 0 0.0014710799999999998 0 0.0014711799999999999 3.3 0.0014711 3.3 0.0014712 0 0.0014711199999999998 0 0.0014712199999999999 3.3 0.00147114 3.3 0.00147124 0 0.00147116 0 0.00147126 3.3 0.0014711799999999999 3.3 0.00147128 0 0.0014712 0 0.0014713 3.3 0.0014712199999999999 3.3 0.00147132 0 0.00147124 0 0.00147134 3.3 0.0014712599999999998 3.3 0.00147136 0 0.00147128 0 0.00147138 3.3 0.0014712999999999998 3.3 0.0014713999999999999 0 0.00147132 0 0.00147142 3.3 0.00147134 3.3 0.00147144 0 0.00147136 0 0.00147146 3.3 0.00147138 3.3 0.00147148 0 0.0014713999999999999 0 0.0014715 3.3 0.00147142 3.3 0.00147152 0 0.0014714399999999999 0 0.00147154 3.3 0.00147146 3.3 0.00147156 0 0.0014714799999999998 0 0.00147158 3.3 0.0014715 3.3 0.0014716 0 0.0014715199999999998 0 0.0014716199999999999 3.3 0.00147154 3.3 0.00147164 0 0.00147156 0 0.00147166 3.3 0.00147158 3.3 0.00147168 0 0.0014716 0 0.0014717 3.3 0.0014716199999999999 3.3 0.00147172 0 0.00147164 0 0.00147174 3.3 0.0014716599999999999 3.3 0.00147176 0 0.00147168 0 0.00147178 3.3 0.0014716999999999998 3.3 0.0014717999999999999 0 0.00147172 0 0.00147182 3.3 0.0014717399999999998 3.3 0.0014718399999999999 0 0.00147176 0 0.00147186 3.3 0.00147178 3.3 0.00147188 0 0.0014717999999999999 0 0.0014719 3.3 0.00147182 3.3 0.00147192 0 0.0014718399999999999 0 0.00147194 3.3 0.00147186 3.3 0.00147196 0 0.0014718799999999998 0 0.00147198 3.3 0.0014719 3.3 0.001472 0 0.0014719199999999998 0 0.0014720199999999999 3.3 0.00147194 3.3 0.00147204 0 0.00147196 0 0.00147206 3.3 0.00147198 3.3 0.00147208 0 0.001472 0 0.0014721 3.3 0.0014720199999999999 3.3 0.00147212 0 0.00147204 0 0.00147214 3.3 0.0014720599999999999 3.3 0.00147216 0 0.00147208 0 0.00147218 3.3 0.0014720999999999998 3.3 0.0014722 0 0.00147212 0 0.00147222 3.3 0.0014721399999999998 3.3 0.0014722399999999999 0 0.00147216 0 0.00147226 3.3 0.00147218 3.3 0.00147228 0 0.0014722 0 0.0014723 3.3 0.00147222 3.3 0.00147232 0 0.0014722399999999999 0 0.00147234 3.3 0.00147226 3.3 0.00147236 0 0.0014722799999999999 0 0.00147238 3.3 0.0014723 3.3 0.0014724 0 0.0014723199999999998 0 0.00147242 3.3 0.00147234 3.3 0.00147244 0 0.0014723599999999998 0 0.0014724599999999999 3.3 0.00147238 3.3 0.00147248 0 0.0014724 0 0.0014725 3.3 0.00147242 3.3 0.00147252 0 0.00147244 0 0.00147254 3.3 0.0014724599999999999 3.3 0.00147256 0 0.00147248 0 0.00147258 3.3 0.0014724999999999999 3.3 0.0014726 0 0.00147252 0 0.00147262 3.3 0.0014725399999999998 3.3 0.0014726399999999999 0 0.00147256 0 0.00147266 3.3 0.0014725799999999998 3.3 0.0014726799999999999 0 0.0014726 0 0.0014727 3.3 0.00147262 3.3 0.00147272 0 0.0014726399999999999 0 0.00147274 3.3 0.00147266 3.3 0.00147276 0 0.0014726799999999999 0 0.00147278 3.3 0.0014727 3.3 0.0014728 0 0.0014727199999999998 0 0.00147282 3.3 0.00147274 3.3 0.00147284 0 0.0014727599999999998 0 0.0014728599999999999 3.3 0.00147278 3.3 0.00147288 0 0.0014728 0 0.0014729 3.3 0.00147282 3.3 0.00147292 0 0.00147284 0 0.00147294 3.3 0.0014728599999999999 3.3 0.00147296 0 0.00147288 0 0.00147298 3.3 0.0014728999999999999 3.3 0.001473 0 0.00147292 0 0.00147302 3.3 0.0014729399999999998 3.3 0.00147304 0 0.00147296 0 0.00147306 3.3 0.0014729799999999998 3.3 0.0014730799999999999 0 0.001473 0 0.0014731 3.3 0.00147302 3.3 0.00147312 0 0.00147304 0 0.00147314 3.3 0.00147306 3.3 0.00147316 0 0.0014730799999999999 0 0.00147318 3.3 0.0014731 3.3 0.0014732 0 0.0014731199999999999 0 0.00147322 3.3 0.00147314 3.3 0.00147324 0 0.0014731599999999998 0 0.0014732599999999999 3.3 0.00147318 3.3 0.00147328 0 0.0014731999999999998 0 0.0014732999999999999 3.3 0.00147322 3.3 0.00147332 0 0.00147324 0 0.00147334 3.3 0.0014732599999999999 3.3 0.00147336 0 0.00147328 0 0.00147338 3.3 0.0014732999999999999 3.3 0.0014734 0 0.00147332 0 0.00147342 3.3 0.0014733399999999998 3.3 0.00147344 0 0.00147336 0 0.00147346 3.3 0.0014733799999999998 3.3 0.0014734799999999999 0 0.0014734 0 0.0014735 3.3 0.0014734199999999998 3.3 0.0014735199999999999 0 0.00147344 0 0.00147354 3.3 0.00147346 3.3 0.00147356 0 0.0014734799999999999 0 0.00147358 3.3 0.0014735 3.3 0.0014736 0 0.0014735199999999999 0 0.00147362 3.3 0.00147354 3.3 0.00147364 0 0.0014735599999999998 0 0.00147366 3.3 0.00147358 3.3 0.00147368 0 0.0014735999999999998 0 0.0014736999999999999 3.3 0.00147362 3.3 0.00147372 0 0.00147364 0 0.00147374 3.3 0.00147366 3.3 0.00147376 0 0.00147368 0 0.00147378 3.3 0.0014736999999999999 3.3 0.0014738 0 0.00147372 0 0.00147382 3.3 0.0014737399999999999 3.3 0.00147384 0 0.00147376 0 0.00147386 3.3 0.0014737799999999998 3.3 0.00147388 0 0.0014738 0 0.0014739 3.3 0.0014738199999999998 3.3 0.0014739199999999999 0 0.00147384 0 0.00147394 3.3 0.00147386 3.3 0.00147396 0 0.00147388 0 0.00147398 3.3 0.0014739 3.3 0.001474 0 0.0014739199999999999 0 0.00147402 3.3 0.00147394 3.3 0.00147404 0 0.0014739599999999999 0 0.00147406 3.3 0.00147398 3.3 0.00147408 0 0.0014739999999999998 0 0.0014740999999999999 3.3 0.00147402 3.3 0.00147412 0 0.0014740399999999998 0 0.0014741399999999999 3.3 0.00147406 3.3 0.00147416 0 0.00147408 0 0.00147418 3.3 0.0014740999999999999 3.3 0.0014742 0 0.00147412 0 0.00147422 3.3 0.0014741399999999999 3.3 0.00147424 0 0.00147416 0 0.00147426 3.3 0.0014741799999999998 3.3 0.00147428 0 0.0014742 0 0.0014743 3.3 0.0014742199999999998 3.3 0.0014743199999999999 0 0.00147424 0 0.00147434 3.3 0.0014742599999999998 3.3 0.0014743599999999999 0 0.00147428 0 0.00147438 3.3 0.0014743 3.3 0.0014744 0 0.0014743199999999999 0 0.00147442 3.3 0.00147434 3.3 0.00147444 0 0.0014743599999999999 0 0.00147446 3.3 0.00147438 3.3 0.00147448 0 0.0014743999999999998 0 0.0014745 3.3 0.00147442 3.3 0.00147452 0 0.0014744399999999998 0 0.0014745399999999999 3.3 0.00147446 3.3 0.00147456 0 0.00147448 0 0.00147458 3.3 0.0014745 3.3 0.0014746 0 0.00147452 0 0.00147462 3.3 0.0014745399999999999 3.3 0.00147464 0 0.00147456 0 0.00147466 3.3 0.0014745799999999999 3.3 0.00147468 0 0.0014746 0 0.0014747 3.3 0.0014746199999999998 3.3 0.00147472 0 0.00147464 0 0.00147474 3.3 0.0014746599999999998 3.3 0.0014747599999999999 0 0.00147468 0 0.00147478 3.3 0.0014747 3.3 0.0014748 0 0.00147472 0 0.00147482 3.3 0.00147474 3.3 0.00147484 0 0.0014747599999999999 0 0.00147486 3.3 0.00147478 3.3 0.00147488 0 0.0014747999999999999 0 0.0014749 3.3 0.00147482 3.3 0.00147492 0 0.0014748399999999998 0 0.0014749399999999999 3.3 0.00147486 3.3 0.00147496 0 0.0014748799999999998 0 0.0014749799999999999 3.3 0.0014749 3.3 0.001475 0 0.00147492 0 0.00147502 3.3 0.0014749399999999999 3.3 0.00147504 0 0.00147496 0 0.00147506 3.3 0.0014749799999999999 3.3 0.00147508 0 0.001475 0 0.0014751 3.3 0.0014750199999999998 3.3 0.00147512 0 0.00147504 0 0.00147514 3.3 0.0014750599999999998 3.3 0.0014751599999999999 0 0.00147508 0 0.00147518 3.3 0.0014750999999999998 3.3 0.0014751999999999999 0 0.00147512 0 0.00147522 3.3 0.00147514 3.3 0.00147524 0 0.0014751599999999999 0 0.00147526 3.3 0.00147518 3.3 0.00147528 0 0.0014751999999999999 0 0.0014753 3.3 0.00147522 3.3 0.00147532 0 0.0014752399999999998 0 0.00147534 3.3 0.00147526 3.3 0.00147536 0 0.0014752799999999998 0 0.0014753799999999999 3.3 0.0014753 3.3 0.0014754 0 0.00147532 0 0.00147542 3.3 0.00147534 3.3 0.00147544 0 0.00147536 0 0.00147546 3.3 0.0014753799999999999 3.3 0.00147548 0 0.0014754 0 0.0014755 3.3 0.0014754199999999999 3.3 0.00147552 0 0.00147544 0 0.00147554 3.3 0.0014754599999999998 3.3 0.00147556 0 0.00147548 0 0.00147558 3.3 0.0014754999999999998 3.3 0.0014755999999999999 0 0.00147552 0 0.00147562 3.3 0.00147554 3.3 0.00147564 0 0.00147556 0 0.00147566 3.3 0.00147558 3.3 0.00147568 0 0.0014755999999999999 0 0.0014757 3.3 0.00147562 3.3 0.00147572 0 0.0014756399999999999 0 0.00147574 3.3 0.00147566 3.3 0.00147576 0 0.0014756799999999998 0 0.0014757799999999999 3.3 0.0014757 3.3 0.0014758 0 0.0014757199999999998 0 0.0014758199999999999 3.3 0.00147574 3.3 0.00147584 0 0.00147576 0 0.00147586 3.3 0.0014757799999999999 3.3 0.00147588 0 0.0014758 0 0.0014759 3.3 0.0014758199999999999 3.3 0.00147592 0 0.00147584 0 0.00147594 3.3 0.0014758599999999998 3.3 0.00147596 0 0.00147588 0 0.00147598 3.3 0.0014758999999999998 3.3 0.0014759999999999999 0 0.00147592 0 0.00147602 3.3 0.00147594 3.3 0.00147604 0 0.00147596 0 0.00147606 3.3 0.00147598 3.3 0.00147608 0 0.0014759999999999999 0 0.0014761 3.3 0.00147602 3.3 0.00147612 0 0.0014760399999999999 0 0.00147614 3.3 0.00147606 3.3 0.00147616 0 0.0014760799999999998 0 0.00147618 3.3 0.0014761 3.3 0.0014762 0 0.0014761199999999998 0 0.0014762199999999999 3.3 0.00147614 3.3 0.00147624 0 0.00147616 0 0.00147626 3.3 0.00147618 3.3 0.00147628 0 0.0014762 0 0.0014763 3.3 0.0014762199999999999 3.3 0.00147632 0 0.00147624 0 0.00147634 3.3 0.0014762599999999999 3.3 0.00147636 0 0.00147628 0 0.00147638 3.3 0.0014762999999999998 3.3 0.0014763999999999999 0 0.00147632 0 0.00147642 3.3 0.0014763399999999998 3.3 0.0014764399999999999 0 0.00147636 0 0.00147646 3.3 0.00147638 3.3 0.00147648 0 0.0014763999999999999 0 0.0014765 3.3 0.00147642 3.3 0.00147652 0 0.0014764399999999999 0 0.00147654 3.3 0.00147646 3.3 0.00147656 0 0.0014764799999999998 0 0.00147658 3.3 0.0014765 3.3 0.0014766 0 0.0014765199999999998 0 0.0014766199999999999 3.3 0.00147654 3.3 0.00147664 0 0.0014765599999999998 0 0.0014766599999999999 3.3 0.00147658 3.3 0.00147668 0 0.0014766 0 0.0014767 3.3 0.0014766199999999999 3.3 0.00147672 0 0.00147664 0 0.00147674 3.3 0.0014766599999999999 3.3 0.00147676 0 0.00147668 0 0.00147678 3.3 0.0014766999999999998 3.3 0.0014768 0 0.00147672 0 0.00147682 3.3 0.0014767399999999998 3.3 0.0014768399999999999 0 0.00147676 0 0.00147686 3.3 0.00147678 3.3 0.00147688 0 0.0014768 0 0.0014769 3.3 0.00147682 3.3 0.00147692 0 0.0014768399999999999 0 0.00147694 3.3 0.00147686 3.3 0.00147696 0 0.0014768799999999999 0 0.00147698 3.3 0.0014769 3.3 0.001477 0 0.0014769199999999998 0 0.00147702 3.3 0.00147694 3.3 0.00147704 0 0.0014769599999999998 0 0.0014770599999999999 3.3 0.00147698 3.3 0.00147708 0 0.001477 0 0.0014771 3.3 0.00147702 3.3 0.00147712 0 0.00147704 0 0.00147714 3.3 0.0014770599999999999 3.3 0.00147716 0 0.00147708 0 0.00147718 3.3 0.0014770999999999999 3.3 0.0014772 0 0.00147712 0 0.00147722 3.3 0.0014771399999999998 3.3 0.0014772399999999999 0 0.00147716 0 0.00147726 3.3 0.0014771799999999998 3.3 0.0014772799999999999 0 0.0014772 0 0.0014773 3.3 0.00147722 3.3 0.00147732 0 0.0014772399999999999 0 0.00147734 3.3 0.00147726 3.3 0.00147736 0 0.0014772799999999999 0 0.00147738 3.3 0.0014773 3.3 0.0014774 0 0.0014773199999999998 0 0.00147742 3.3 0.00147734 3.3 0.00147744 0 0.0014773599999999998 0 0.0014774599999999999 3.3 0.00147738 3.3 0.00147748 0 0.0014773999999999998 0 0.0014774999999999999 3.3 0.00147742 3.3 0.00147752 0 0.00147744 0 0.00147754 3.3 0.0014774599999999999 3.3 0.00147756 0 0.00147748 0 0.00147758 3.3 0.0014774999999999999 3.3 0.0014776 0 0.00147752 0 0.00147762 3.3 0.0014775399999999998 3.3 0.00147764 0 0.00147756 0 0.00147766 3.3 0.0014775799999999998 3.3 0.0014776799999999999 0 0.0014776 0 0.0014777 3.3 0.00147762 3.3 0.00147772 0 0.00147764 0 0.00147774 3.3 0.00147766 3.3 0.00147776 0 0.0014776799999999999 0 0.00147778 3.3 0.0014777 3.3 0.0014778 0 0.0014777199999999999 0 0.00147782 3.3 0.00147774 3.3 0.00147784 0 0.0014777599999999998 0 0.00147786 3.3 0.00147778 3.3 0.00147788 0 0.0014777999999999998 0 0.0014778999999999999 3.3 0.00147782 3.3 0.00147792 0 0.00147784 0 0.00147794 3.3 0.00147786 3.3 0.00147796 0 0.00147788 0 0.00147798 3.3 0.0014778999999999999 3.3 0.001478 0 0.00147792 0 0.00147802 3.3 0.0014779399999999999 3.3 0.00147804 0 0.00147796 0 0.00147806 3.3 0.0014779799999999998 3.3 0.0014780799999999999 0 0.001478 0 0.0014781 3.3 0.0014780199999999998 3.3 0.0014781199999999999 0 0.00147804 0 0.00147814 3.3 0.00147806 3.3 0.00147816 0 0.0014780799999999999 0 0.00147818 3.3 0.0014781 3.3 0.0014782 0 0.0014781199999999999 0 0.00147822 3.3 0.00147814 3.3 0.00147824 0 0.0014781599999999998 0 0.00147826 3.3 0.00147818 3.3 0.00147828 0 0.0014781999999999998 0 0.0014782999999999999 3.3 0.00147822 3.3 0.00147832 0 0.0014782399999999998 0 0.0014783399999999999 3.3 0.00147826 3.3 0.00147836 0 0.00147828 0 0.00147838 3.3 0.0014782999999999999 3.3 0.0014784 0 0.00147832 0 0.00147842 3.3 0.0014783399999999999 3.3 0.00147844 0 0.00147836 0 0.00147846 3.3 0.0014783799999999998 3.3 0.00147848 0 0.0014784 0 0.0014785 3.3 0.0014784199999999998 3.3 0.0014785199999999999 0 0.00147844 0 0.00147854 3.3 0.00147846 3.3 0.00147856 0 0.00147848 0 0.00147858 3.3 0.0014785 3.3 0.0014786 0 0.0014785199999999999 0 0.00147862 3.3 0.00147854 3.3 0.00147864 0 0.0014785599999999999 0 0.00147866 3.3 0.00147858 3.3 0.00147868 0 0.0014785999999999998 0 0.0014787 3.3 0.00147862 3.3 0.00147872 0 0.0014786399999999998 0 0.0014787399999999999 3.3 0.00147866 3.3 0.00147876 0 0.00147868 0 0.00147878 3.3 0.0014787 3.3 0.0014788 0 0.00147872 0 0.00147882 3.3 0.0014787399999999999 3.3 0.00147884 0 0.00147876 0 0.00147886 3.3 0.0014787799999999999 3.3 0.00147888 0 0.0014788 0 0.0014789 3.3 0.0014788199999999998 3.3 0.0014789199999999999 0 0.00147884 0 0.00147894 3.3 0.0014788599999999998 3.3 0.0014789599999999999 0 0.00147888 0 0.00147898 3.3 0.0014789 3.3 0.001479 0 0.0014789199999999999 0 0.00147902 3.3 0.00147894 3.3 0.00147904 0 0.0014789599999999999 0 0.00147906 3.3 0.00147898 3.3 0.00147908 0 0.0014789999999999998 0 0.0014791 3.3 0.00147902 3.3 0.00147912 0 0.0014790399999999998 0 0.0014791399999999999 3.3 0.00147906 3.3 0.00147916 0 0.00147908 0 0.00147918 3.3 0.0014791 3.3 0.0014792 0 0.00147912 0 0.00147922 3.3 0.0014791399999999999 3.3 0.00147924 0 0.00147916 0 0.00147926 3.3 0.0014791799999999999 3.3 0.00147928 0 0.0014792 0 0.0014793 3.3 0.0014792199999999998 3.3 0.00147932 0 0.00147924 0 0.00147934 3.3 0.0014792599999999998 3.3 0.0014793599999999999 0 0.00147928 0 0.00147938 3.3 0.0014793 3.3 0.0014794 0 0.00147932 0 0.00147942 3.3 0.00147934 3.3 0.00147944 0 0.0014793599999999999 0 0.00147946 3.3 0.00147938 3.3 0.00147948 0 0.0014793999999999999 0 0.0014795 3.3 0.00147942 3.3 0.00147952 0 0.0014794399999999998 0 0.00147954 3.3 0.00147946 3.3 0.00147956 0 0.0014794799999999998 0 0.0014795799999999999 3.3 0.0014795 3.3 0.0014796 0 0.00147952 0 0.00147962 3.3 0.00147954 3.3 0.00147964 0 0.00147956 0 0.00147966 3.3 0.0014795799999999999 3.3 0.00147968 0 0.0014796 0 0.0014797 3.3 0.0014796199999999999 3.3 0.00147972 0 0.00147964 0 0.00147974 3.3 0.0014796599999999998 3.3 0.0014797599999999999 0 0.00147968 0 0.00147978 3.3 0.0014796999999999998 3.3 0.0014797999999999999 0 0.00147972 0 0.00147982 3.3 0.00147974 3.3 0.00147984 0 0.0014797599999999999 0 0.00147986 3.3 0.00147978 3.3 0.00147988 0 0.0014797999999999999 0 0.0014799 3.3 0.00147982 3.3 0.00147992 0 0.0014798399999999998 0 0.00147994 3.3 0.00147986 3.3 0.00147996 0 0.0014798799999999998 0 0.0014799799999999999 3.3 0.0014799 3.3 0.00148 0 0.00147992 0 0.00148002 3.3 0.00147994 3.3 0.00148004 0 0.00147996 0 0.00148006 3.3 0.0014799799999999999 3.3 0.00148008 0 0.00148 0 0.0014801 3.3 0.0014800199999999999 3.3 0.00148012 0 0.00148004 0 0.00148014 3.3 0.0014800599999999998 3.3 0.00148016 0 0.00148008 0 0.00148018 3.3 0.0014800999999999998 3.3 0.0014801999999999999 0 0.00148012 0 0.00148022 3.3 0.00148014 3.3 0.00148024 0 0.00148016 0 0.00148026 3.3 0.00148018 3.3 0.00148028 0 0.0014801999999999999 0 0.0014803 3.3 0.00148022 3.3 0.00148032 0 0.0014802399999999999 0 0.00148034 3.3 0.00148026 3.3 0.00148036 0 0.0014802799999999998 0 0.0014803799999999999 3.3 0.0014803 3.3 0.0014804 0 0.0014803199999999998 0 0.0014804199999999999 3.3 0.00148034 3.3 0.00148044 0 0.00148036 0 0.00148046 3.3 0.0014803799999999999 3.3 0.00148048 0 0.0014804 0 0.0014805 3.3 0.0014804199999999999 3.3 0.00148052 0 0.00148044 0 0.00148054 3.3 0.0014804599999999998 3.3 0.00148056 0 0.00148048 0 0.00148058 3.3 0.0014804999999999998 3.3 0.0014805999999999999 0 0.00148052 0 0.00148062 3.3 0.0014805399999999998 3.3 0.0014806399999999999 0 0.00148056 0 0.00148066 3.3 0.00148058 3.3 0.00148068 0 0.0014805999999999999 0 0.0014807 3.3 0.00148062 3.3 0.00148072 0 0.0014806399999999999 0 0.00148074 3.3 0.00148066 3.3 0.00148076 0 0.0014806799999999998 0 0.00148078 3.3 0.0014807 3.3 0.0014808 0 0.0014807199999999998 0 0.0014808199999999999 3.3 0.00148074 3.3 0.00148084 0 0.00148076 0 0.00148086 3.3 0.00148078 3.3 0.00148088 0 0.0014808 0 0.0014809 3.3 0.0014808199999999999 3.3 0.00148092 0 0.00148084 0 0.00148094 3.3 0.0014808599999999999 3.3 0.00148096 0 0.00148088 0 0.00148098 3.3 0.0014808999999999998 3.3 0.001481 0 0.00148092 0 0.00148102 3.3 0.0014809399999999998 3.3 0.0014810399999999999 0 0.00148096 0 0.00148106 3.3 0.00148098 3.3 0.00148108 0 0.001481 0 0.0014811 3.3 0.00148102 3.3 0.00148112 0 0.0014810399999999999 0 0.00148114 3.3 0.00148106 3.3 0.00148116 0 0.0014810799999999999 0 0.00148118 3.3 0.0014811 3.3 0.0014812 0 0.0014811199999999998 0 0.0014812199999999999 3.3 0.00148114 3.3 0.00148124 0 0.0014811599999999998 0 0.0014812599999999999 3.3 0.00148118 3.3 0.00148128 0 0.0014812 0 0.0014813 3.3 0.0014812199999999999 3.3 0.00148132 0 0.00148124 0 0.00148134 3.3 0.0014812599999999999 3.3 0.00148136 0 0.00148128 0 0.00148138 3.3 0.0014812999999999998 3.3 0.0014814 0 0.00148132 0 0.00148142 3.3 0.0014813399999999998 3.3 0.0014814399999999999 0 0.00148136 0 0.00148146 3.3 0.0014813799999999998 3.3 0.0014814799999999999 0 0.0014814 0 0.0014815 3.3 0.00148142 3.3 0.00148152 0 0.0014814399999999999 0 0.00148154 3.3 0.00148146 3.3 0.00148156 0 0.0014814799999999999 0 0.00148158 3.3 0.0014815 3.3 0.0014816 0 0.0014815199999999998 0 0.00148162 3.3 0.00148154 3.3 0.00148164 0 0.0014815599999999998 0 0.0014816599999999999 3.3 0.00148158 3.3 0.00148168 0 0.0014816 0 0.0014817 3.3 0.00148162 3.3 0.00148172 0 0.00148164 0 0.00148174 3.3 0.0014816599999999999 3.3 0.00148176 0 0.00148168 0 0.00148178 3.3 0.0014816999999999999 3.3 0.0014818 0 0.00148172 0 0.00148182 3.3 0.0014817399999999998 3.3 0.00148184 0 0.00148176 0 0.00148186 3.3 0.0014817799999999998 3.3 0.0014818799999999999 0 0.0014818 0 0.0014819 3.3 0.00148182 3.3 0.00148192 0 0.00148184 0 0.00148194 3.3 0.00148186 3.3 0.00148196 0 0.0014818799999999999 0 0.00148198 3.3 0.0014819 3.3 0.001482 0 0.0014819199999999999 0 0.00148202 3.3 0.00148194 3.3 0.00148204 0 0.0014819599999999998 0 0.0014820599999999999 3.3 0.00148198 3.3 0.00148208 0 0.0014819999999999998 0 0.0014820999999999999 3.3 0.00148202 3.3 0.00148212 0 0.00148204 0 0.00148214 3.3 0.0014820599999999999 3.3 0.00148216 0 0.00148208 0 0.00148218 3.3 0.0014820999999999999 3.3 0.0014822 0 0.00148212 0 0.00148222 3.3 0.0014821399999999998 3.3 0.00148224 0 0.00148216 0 0.00148226 3.3 0.0014821799999999998 3.3 0.0014822799999999999 0 0.0014822 0 0.0014823 3.3 0.00148222 3.3 0.00148232 0 0.00148224 0 0.00148234 3.3 0.00148226 3.3 0.00148236 0 0.0014822799999999999 0 0.00148238 3.3 0.0014823 3.3 0.0014824 0 0.0014823199999999999 0 0.00148242 3.3 0.00148234 3.3 0.00148244 0 0.0014823599999999998 0 0.00148246 3.3 0.00148238 3.3 0.00148248 0 0.0014823999999999998 0 0.0014824999999999999 3.3 0.00148242 3.3 0.00148252 0 0.00148244 0 0.00148254 3.3 0.00148246 3.3 0.00148256 0 0.00148248 0 0.00148258 3.3 0.0014824999999999999 3.3 0.0014826 0 0.00148252 0 0.00148262 3.3 0.0014825399999999999 3.3 0.00148264 0 0.00148256 0 0.00148266 3.3 0.0014825799999999998 3.3 0.00148268 0 0.0014826 0 0.0014827 3.3 0.0014826199999999998 3.3 0.0014827199999999999 0 0.00148264 0 0.00148274 3.3 0.00148266 3.3 0.00148276 0 0.00148268 0 0.00148278 3.3 0.0014827 3.3 0.0014828 0 0.0014827199999999999 0 0.00148282 3.3 0.00148274 3.3 0.00148284 0 0.0014827599999999999 0 0.00148286 3.3 0.00148278 3.3 0.00148288 0 0.0014827999999999998 0 0.0014828999999999999 3.3 0.00148282 3.3 0.00148292 0 0.0014828399999999998 0 0.0014829399999999999 3.3 0.00148286 3.3 0.00148296 0 0.00148288 0 0.00148298 3.3 0.0014828999999999999 3.3 0.001483 0 0.00148292 0 0.00148302 3.3 0.0014829399999999999 3.3 0.00148304 0 0.00148296 0 0.00148306 3.3 0.0014829799999999998 3.3 0.00148308 0 0.001483 0 0.0014831 3.3 0.0014830199999999998 3.3 0.0014831199999999999 0 0.00148304 0 0.00148314 3.3 0.00148306 3.3 0.00148316 0 0.00148308 0 0.00148318 3.3 0.0014831 3.3 0.0014832 0 0.0014831199999999999 0 0.00148322 3.3 0.00148314 3.3 0.00148324 0 0.0014831599999999999 0 0.00148326 3.3 0.00148318 3.3 0.00148328 0 0.0014831999999999998 0 0.0014833 3.3 0.00148322 3.3 0.00148332 0 0.0014832399999999998 0 0.0014833399999999999 3.3 0.00148326 3.3 0.00148336 0 0.00148328 0 0.00148338 3.3 0.0014833 3.3 0.0014834 0 0.00148332 0 0.00148342 3.3 0.0014833399999999999 3.3 0.00148344 0 0.00148336 0 0.00148346 3.3 0.0014833799999999999 3.3 0.00148348 0 0.0014834 0 0.0014835 3.3 0.0014834199999999998 3.3 0.0014835199999999999 0 0.00148344 0 0.00148354 3.3 0.0014834599999999998 3.3 0.0014835599999999999 0 0.00148348 0 0.00148358 3.3 0.0014835 3.3 0.0014836 0 0.0014835199999999999 0 0.00148362 3.3 0.00148354 3.3 0.00148364 0 0.0014835599999999999 0 0.00148366 3.3 0.00148358 3.3 0.00148368 0 0.0014835999999999998 0 0.0014837 3.3 0.00148362 3.3 0.00148372 0 0.0014836399999999998 0 0.0014837399999999999 3.3 0.00148366 3.3 0.00148376 0 0.0014836799999999998 0 0.0014837799999999999 3.3 0.0014837 3.3 0.0014838 0 0.00148372 0 0.00148382 3.3 0.0014837399999999999 3.3 0.00148384 0 0.00148376 0 0.00148386 3.3 0.0014837799999999999 3.3 0.00148388 0 0.0014838 0 0.0014839 3.3 0.0014838199999999998 3.3 0.00148392 0 0.00148384 0 0.00148394 3.3 0.0014838599999999998 3.3 0.0014839599999999999 0 0.00148388 0 0.00148398 3.3 0.0014839 3.3 0.001484 0 0.00148392 0 0.00148402 3.3 0.00148394 3.3 0.00148404 0 0.0014839599999999999 0 0.00148406 3.3 0.00148398 3.3 0.00148408 0 0.0014839999999999999 0 0.0014841 3.3 0.00148402 3.3 0.00148412 0 0.0014840399999999998 0 0.00148414 3.3 0.00148406 3.3 0.00148416 0 0.0014840799999999998 0 0.0014841799999999999 3.3 0.0014841 3.3 0.0014842 0 0.00148412 0 0.00148422 3.3 0.00148414 3.3 0.00148424 0 0.00148416 0 0.00148426 3.3 0.0014841799999999999 3.3 0.00148428 0 0.0014842 0 0.0014843 3.3 0.0014842199999999999 3.3 0.00148432 0 0.00148424 0 0.00148434 3.3 0.0014842599999999998 3.3 0.0014843599999999999 0 0.00148428 0 0.00148438 3.3 0.0014842999999999998 3.3 0.0014843999999999999 0 0.00148432 0 0.00148442 3.3 0.00148434 3.3 0.00148444 0 0.0014843599999999999 0 0.00148446 3.3 0.00148438 3.3 0.00148448 0 0.0014843999999999999 0 0.0014845 3.3 0.00148442 3.3 0.00148452 0 0.0014844399999999998 0 0.00148454 3.3 0.00148446 3.3 0.00148456 0 0.0014844799999999998 0 0.0014845799999999999 3.3 0.0014845 3.3 0.0014846 0 0.0014845199999999998 0 0.0014846199999999999 3.3 0.00148454 3.3 0.00148464 0 0.00148456 0 0.00148466 3.3 0.0014845799999999999 3.3 0.00148468 0 0.0014846 0 0.0014847 3.3 0.0014846199999999999 3.3 0.00148472 0 0.00148464 0 0.00148474 3.3 0.0014846599999999998 3.3 0.00148476 0 0.00148468 0 0.00148478 3.3 0.0014846999999999998 3.3 0.0014847999999999999 0 0.00148472 0 0.00148482 3.3 0.00148474 3.3 0.00148484 0 0.00148476 0 0.00148486 3.3 0.00148478 3.3 0.00148488 0 0.0014847999999999999 0 0.0014849 3.3 0.00148482 3.3 0.00148492 0 0.0014848399999999999 0 0.00148494 3.3 0.00148486 3.3 0.00148496 0 0.0014848799999999998 0 0.00148498 3.3 0.0014849 3.3 0.001485 0 0.0014849199999999998 0 0.0014850199999999999 3.3 0.00148494 3.3 0.00148504 0 0.00148496 0 0.00148506 3.3 0.00148498 3.3 0.00148508 0 0.001485 0 0.0014851 3.3 0.0014850199999999999 3.3 0.00148512 0 0.00148504 0 0.00148514 3.3 0.0014850599999999999 3.3 0.00148516 0 0.00148508 0 0.00148518 3.3 0.0014850999999999998 3.3 0.0014851999999999999 0 0.00148512 0 0.00148522 3.3 0.0014851399999999998 3.3 0.0014852399999999999 0 0.00148516 0 0.00148526 3.3 0.00148518 3.3 0.00148528 0 0.0014851999999999999 0 0.0014853 3.3 0.00148522 3.3 0.00148532 0 0.0014852399999999999 0 0.00148534 3.3 0.00148526 3.3 0.00148536 0 0.0014852799999999998 0 0.00148538 3.3 0.0014853 3.3 0.0014854 0 0.0014853199999999998 0 0.0014854199999999999 3.3 0.00148534 3.3 0.00148544 0 0.0014853599999999998 0 0.0014854599999999999 3.3 0.00148538 3.3 0.00148548 0 0.0014854 0 0.0014855 3.3 0.0014854199999999999 3.3 0.00148552 0 0.00148544 0 0.00148554 3.3 0.0014854599999999999 3.3 0.00148556 0 0.00148548 0 0.00148558 3.3 0.0014854999999999998 3.3 0.0014856 0 0.00148552 0 0.00148562 3.3 0.0014855399999999998 3.3 0.0014856399999999999 0 0.00148556 0 0.00148566 3.3 0.00148558 3.3 0.00148568 0 0.0014856 0 0.0014857 3.3 0.00148562 3.3 0.00148572 0 0.0014856399999999999 0 0.00148574 3.3 0.00148566 3.3 0.00148576 0 0.0014856799999999999 0 0.00148578 3.3 0.0014857 3.3 0.0014858 0 0.0014857199999999998 0 0.00148582 3.3 0.00148574 3.3 0.00148584 0 0.0014857599999999998 0 0.0014858599999999999 3.3 0.00148578 3.3 0.00148588 0 0.0014858 0 0.0014859 3.3 0.00148582 3.3 0.00148592 0 0.00148584 0 0.00148594 3.3 0.0014858599999999999 3.3 0.00148596 0 0.00148588 0 0.00148598 3.3 0.0014858999999999999 3.3 0.001486 0 0.00148592 0 0.00148602 3.3 0.0014859399999999998 3.3 0.0014860399999999999 0 0.00148596 0 0.00148606 3.3 0.0014859799999999998 3.3 0.0014860799999999999 0 0.001486 0 0.0014861 3.3 0.00148602 3.3 0.00148612 0 0.0014860399999999999 0 0.00148614 3.3 0.00148606 3.3 0.00148616 0 0.0014860799999999999 0 0.00148618 3.3 0.0014861 3.3 0.0014862 0 0.0014861199999999998 0 0.00148622 3.3 0.00148614 3.3 0.00148624 0 0.0014861599999999998 0 0.0014862599999999999 3.3 0.00148618 3.3 0.00148628 0 0.0014862 0 0.0014863 3.3 0.00148622 3.3 0.00148632 0 0.00148624 0 0.00148634 3.3 0.0014862599999999999 3.3 0.00148636 0 0.00148628 0 0.00148638 3.3 0.0014862999999999999 3.3 0.0014864 0 0.00148632 0 0.00148642 3.3 0.0014863399999999998 3.3 0.00148644 0 0.00148636 0 0.00148646 3.3 0.0014863799999999998 3.3 0.0014864799999999999 0 0.0014864 0 0.0014865 3.3 0.00148642 3.3 0.00148652 0 0.00148644 0 0.00148654 3.3 0.00148646 3.3 0.00148656 0 0.0014864799999999999 0 0.00148658 3.3 0.0014865 3.3 0.0014866 0 0.0014865199999999999 0 0.00148662 3.3 0.00148654 3.3 0.00148664 0 0.0014865599999999998 0 0.0014866599999999999 3.3 0.00148658 3.3 0.00148668 0 0.0014865999999999998 0 0.0014866999999999999 3.3 0.00148662 3.3 0.00148672 0 0.00148664 0 0.00148674 3.3 0.0014866599999999999 3.3 0.00148676 0 0.00148668 0 0.00148678 3.3 0.0014866999999999999 3.3 0.0014868 0 0.00148672 0 0.00148682 3.3 0.0014867399999999998 3.3 0.00148684 0 0.00148676 0 0.00148686 3.3 0.0014867799999999998 3.3 0.0014868799999999999 0 0.0014868 0 0.0014869 3.3 0.0014868199999999998 3.3 0.0014869199999999999 0 0.00148684 0 0.00148694 3.3 0.00148686 3.3 0.00148696 0 0.0014868799999999999 0 0.00148698 3.3 0.0014869 3.3 0.001487 0 0.0014869199999999999 0 0.00148702 3.3 0.00148694 3.3 0.00148704 0 0.0014869599999999998 0 0.00148706 3.3 0.00148698 3.3 0.00148708 0 0.0014869999999999998 0 0.0014870999999999999 3.3 0.00148702 3.3 0.00148712 0 0.00148704 0 0.00148714 3.3 0.00148706 3.3 0.00148716 0 0.00148708 0 0.00148718 3.3 0.0014870999999999999 3.3 0.0014872 0 0.00148712 0 0.00148722 3.3 0.0014871399999999999 3.3 0.00148724 0 0.00148716 0 0.00148726 3.3 0.0014871799999999998 3.3 0.00148728 0 0.0014872 0 0.0014873 3.3 0.0014872199999999998 3.3 0.0014873199999999999 0 0.00148724 0 0.00148734 3.3 0.00148726 3.3 0.00148736 0 0.00148728 0 0.00148738 3.3 0.0014873 3.3 0.0014874 0 0.0014873199999999999 0 0.00148742 3.3 0.00148734 3.3 0.00148744 0 0.0014873599999999999 0 0.00148746 3.3 0.00148738 3.3 0.00148748 0 0.0014873999999999998 0 0.0014874999999999999 3.3 0.00148742 3.3 0.00148752 0 0.0014874399999999998 0 0.0014875399999999999 3.3 0.00148746 3.3 0.00148756 0 0.00148748 0 0.00148758 3.3 0.0014874999999999999 3.3 0.0014876 0 0.00148752 0 0.00148762 3.3 0.0014875399999999999 3.3 0.00148764 0 0.00148756 0 0.00148766 3.3 0.0014875799999999998 3.3 0.00148768 0 0.0014876 0 0.0014877 3.3 0.0014876199999999998 3.3 0.0014877199999999999 0 0.00148764 0 0.00148774 3.3 0.0014876599999999998 3.3 0.0014877599999999999 0 0.00148768 0 0.00148778 3.3 0.0014877 3.3 0.0014878 0 0.0014877199999999999 0 0.00148782 3.3 0.00148774 3.3 0.00148784 0 0.0014877599999999999 0 0.00148786 3.3 0.00148778 3.3 0.00148788 0 0.0014877999999999998 0 0.0014879 3.3 0.00148782 3.3 0.00148792 0 0.0014878399999999998 0 0.0014879399999999999 3.3 0.00148786 3.3 0.00148796 0 0.00148788 0 0.00148798 3.3 0.0014879 3.3 0.001488 0 0.00148792 0 0.00148802 3.3 0.0014879399999999999 3.3 0.00148804 0 0.00148796 0 0.00148806 3.3 0.0014879799999999999 3.3 0.00148808 0 0.001488 0 0.0014881 3.3 0.0014880199999999998 3.3 0.00148812 0 0.00148804 0 0.00148814 3.3 0.0014880599999999998 3.3 0.0014881599999999999 0 0.00148808 0 0.00148818 3.3 0.0014881 3.3 0.0014882 0 0.00148812 0 0.00148822 3.3 0.00148814 3.3 0.00148824 0 0.0014881599999999999 0 0.00148826 3.3 0.00148818 3.3 0.00148828 0 0.0014881999999999999 0 0.0014883 3.3 0.00148822 3.3 0.00148832 0 0.0014882399999999998 0 0.0014883399999999999 3.3 0.00148826 3.3 0.00148836 0 0.0014882799999999998 0 0.0014883799999999999 3.3 0.0014883 3.3 0.0014884 0 0.00148832 0 0.00148842 3.3 0.0014883399999999999 3.3 0.00148844 0 0.00148836 0 0.00148846 3.3 0.0014883799999999999 3.3 0.00148848 0 0.0014884 0 0.0014885 3.3 0.0014884199999999998 3.3 0.00148852 0 0.00148844 0 0.00148854 3.3 0.0014884599999999998 3.3 0.0014885599999999999 0 0.00148848 0 0.00148858 3.3 0.0014884999999999998 3.3 0.0014885999999999999 0 0.00148852 0 0.00148862 3.3 0.00148854 3.3 0.00148864 0 0.0014885599999999999 0 0.00148866 3.3 0.00148858 3.3 0.00148868 0 0.0014885999999999999 0 0.0014887 3.3 0.00148862 3.3 0.00148872 0 0.0014886399999999998 0 0.00148874 3.3 0.00148866 3.3 0.00148876 0 0.0014886799999999998 0 0.0014887799999999999 3.3 0.0014887 3.3 0.0014888 0 0.00148872 0 0.00148882 3.3 0.00148874 3.3 0.00148884 0 0.00148876 0 0.00148886 3.3 0.0014887799999999999 3.3 0.00148888 0 0.0014888 0 0.0014889 3.3 0.0014888199999999999 3.3 0.00148892 0 0.00148884 0 0.00148894 3.3 0.0014888599999999998 3.3 0.00148896 0 0.00148888 0 0.00148898 3.3 0.0014888999999999998 3.3 0.0014889999999999999 0 0.00148892 0 0.00148902 3.3 0.00148894 3.3 0.00148904 0 0.00148896 0 0.00148906 3.3 0.00148898 3.3 0.00148908 0 0.0014889999999999999 0 0.0014891 3.3 0.00148902 3.3 0.00148912 0 0.0014890399999999999 0 0.00148914 3.3 0.00148906 3.3 0.00148916 0 0.0014890799999999998 0 0.0014891799999999999 3.3 0.0014891 3.3 0.0014892 0 0.0014891199999999998 0 0.0014892199999999999 3.3 0.00148914 3.3 0.00148924 0 0.00148916 0 0.00148926 3.3 0.0014891799999999999 3.3 0.00148928 0 0.0014892 0 0.0014893 3.3 0.0014892199999999999 3.3 0.00148932 0 0.00148924 0 0.00148934 3.3 0.0014892599999999998 3.3 0.00148936 0 0.00148928 0 0.00148938 3.3 0.0014892999999999998 3.3 0.0014893999999999999 0 0.00148932 0 0.00148942 3.3 0.00148934 3.3 0.00148944 0 0.00148936 0 0.00148946 3.3 0.00148938 3.3 0.00148948 0 0.0014893999999999999 0 0.0014895 3.3 0.00148942 3.3 0.00148952 0 0.0014894399999999999 0 0.00148954 3.3 0.00148946 3.3 0.00148956 0 0.0014894799999999998 0 0.00148958 3.3 0.0014895 3.3 0.0014896 0 0.0014895199999999998 0 0.0014896199999999999 3.3 0.00148954 3.3 0.00148964 0 0.00148956 0 0.00148966 3.3 0.00148958 3.3 0.00148968 0 0.0014896 0 0.0014897 3.3 0.0014896199999999999 3.3 0.00148972 0 0.00148964 0 0.00148974 3.3 0.0014896599999999999 3.3 0.00148976 0 0.00148968 0 0.00148978 3.3 0.0014896999999999998 3.3 0.0014898 0 0.00148972 0 0.00148982 3.3 0.0014897399999999998 3.3 0.0014898399999999999 0 0.00148976 0 0.00148986 3.3 0.00148978 3.3 0.00148988 0 0.0014898 0 0.0014899 3.3 0.00148982 3.3 0.00148992 0 0.0014898399999999999 0 0.00148994 3.3 0.00148986 3.3 0.00148996 0 0.0014898799999999999 0 0.00148998 3.3 0.0014899 3.3 0.00149 0 0.0014899199999999998 0 0.0014900199999999999 3.3 0.00148994 3.3 0.00149004 0 0.0014899599999999998 0 0.0014900599999999999 3.3 0.00148998 3.3 0.00149008 0 0.00149 0 0.0014901 3.3 0.0014900199999999999 3.3 0.00149012 0 0.00149004 0 0.00149014 3.3 0.0014900599999999999 3.3 0.00149016 0 0.00149008 0 0.00149018 3.3 0.0014900999999999998 3.3 0.0014902 0 0.00149012 0 0.00149022 3.3 0.0014901399999999998 3.3 0.0014902399999999999 0 0.00149016 0 0.00149026 3.3 0.00149018 3.3 0.00149028 0 0.0014902 0 0.0014903 3.3 0.00149022 3.3 0.00149032 0 0.0014902399999999999 0 0.00149034 3.3 0.00149026 3.3 0.00149036 0 0.0014902799999999999 0 0.00149038 3.3 0.0014903 3.3 0.0014904 0 0.0014903199999999998 0 0.00149042 3.3 0.00149034 3.3 0.00149044 0 0.0014903599999999998 0 0.0014904599999999999 3.3 0.00149038 3.3 0.00149048 0 0.0014904 0 0.0014905 3.3 0.00149042 3.3 0.00149052 0 0.00149044 0 0.00149054 3.3 0.0014904599999999999 3.3 0.00149056 0 0.00149048 0 0.00149058 3.3 0.0014904999999999999 3.3 0.0014906 0 0.00149052 0 0.00149062 3.3 0.0014905399999999998 3.3 0.0014906399999999999 0 0.00149056 0 0.00149066 3.3 0.0014905799999999998 3.3 0.0014906799999999999 0 0.0014906 0 0.0014907 3.3 0.00149062 3.3 0.00149072 0 0.0014906399999999999 0 0.00149074 3.3 0.00149066 3.3 0.00149076 0 0.0014906799999999999 0 0.00149078 3.3 0.0014907 3.3 0.0014908 0 0.0014907199999999998 0 0.00149082 3.3 0.00149074 3.3 0.00149084 0 0.0014907599999999998 0 0.0014908599999999999 3.3 0.00149078 3.3 0.00149088 0 0.0014907999999999998 0 0.0014908999999999999 3.3 0.00149082 3.3 0.00149092 0 0.00149084 0 0.00149094 3.3 0.0014908599999999999 3.3 0.00149096 0 0.00149088 0 0.00149098 3.3 0.0014908999999999999 3.3 0.001491 0 0.00149092 0 0.00149102 3.3 0.0014909399999999998 3.3 0.00149104 0 0.00149096 0 0.00149106 3.3 0.0014909799999999998 3.3 0.0014910799999999999 0 0.001491 0 0.0014911 3.3 0.00149102 3.3 0.00149112 0 0.00149104 0 0.00149114 3.3 0.00149106 3.3 0.00149116 0 0.0014910799999999999 0 0.00149118 3.3 0.0014911 3.3 0.0014912 0 0.0014911199999999999 0 0.00149122 3.3 0.00149114 3.3 0.00149124 0 0.0014911599999999998 0 0.00149126 3.3 0.00149118 3.3 0.00149128 0 0.0014911999999999998 0 0.0014912999999999999 3.3 0.00149122 3.3 0.00149132 0 0.00149124 0 0.00149134 3.3 0.00149126 3.3 0.00149136 0 0.00149128 0 0.00149138 3.3 0.0014912999999999999 3.3 0.0014914 0 0.00149132 0 0.00149142 3.3 0.0014913399999999999 3.3 0.00149144 0 0.00149136 0 0.00149146 3.3 0.0014913799999999998 3.3 0.0014914799999999999 0 0.0014914 0 0.0014915 3.3 0.0014914199999999998 3.3 0.0014915199999999999 0 0.00149144 0 0.00149154 3.3 0.00149146 3.3 0.00149156 0 0.0014914799999999999 0 0.00149158 3.3 0.0014915 3.3 0.0014916 0 0.0014915199999999999 0 0.00149162 3.3 0.00149154 3.3 0.00149164 0 0.0014915599999999998 0 0.00149166 3.3 0.00149158 3.3 0.00149168 0 0.0014915999999999998 0 0.0014916999999999999 3.3 0.00149162 3.3 0.00149172 0 0.0014916399999999998 0 0.0014917399999999999 3.3 0.00149166 3.3 0.00149176 0 0.00149168 0 0.00149178 3.3 0.0014916999999999999 3.3 0.0014918 0 0.00149172 0 0.00149182 3.3 0.0014917399999999999 3.3 0.00149184 0 0.00149176 0 0.00149186 3.3 0.0014917799999999998 3.3 0.00149188 0 0.0014918 0 0.0014919 3.3 0.0014918199999999998 3.3 0.0014919199999999999 0 0.00149184 0 0.00149194 3.3 0.00149186 3.3 0.00149196 0 0.00149188 0 0.00149198 3.3 0.0014919 3.3 0.001492 0 0.0014919199999999999 0 0.00149202 3.3 0.00149194 3.3 0.00149204 0 0.0014919599999999999 0 0.00149206 3.3 0.00149198 3.3 0.00149208 0 0.0014919999999999998 0 0.0014921 3.3 0.00149202 3.3 0.00149212 0 0.0014920399999999998 0 0.0014921399999999999 3.3 0.00149206 3.3 0.00149216 0 0.00149208 0 0.00149218 3.3 0.0014921 3.3 0.0014922 0 0.00149212 0 0.00149222 3.3 0.0014921399999999999 3.3 0.00149224 0 0.00149216 0 0.00149226 3.3 0.0014921799999999999 3.3 0.00149228 0 0.0014922 0 0.0014923 3.3 0.0014922199999999998 3.3 0.0014923199999999999 0 0.00149224 0 0.00149234 3.3 0.0014922599999999998 3.3 0.0014923599999999999 0 0.00149228 0 0.00149238 3.3 0.0014923 3.3 0.0014924 0 0.0014923199999999999 0 0.00149242 3.3 0.00149234 3.3 0.00149244 0 0.0014923599999999999 0 0.00149246 3.3 0.00149238 3.3 0.00149248 0 0.0014923999999999998 0 0.0014925 3.3 0.00149242 3.3 0.00149252 0 0.0014924399999999998 0 0.0014925399999999999 3.3 0.00149246 3.3 0.00149256 0 0.0014924799999999998 0 0.0014925799999999999 3.3 0.0014925 3.3 0.0014926 0 0.00149252 0 0.00149262 3.3 0.0014925399999999999 3.3 0.00149264 0 0.00149256 0 0.00149266 3.3 0.0014925799999999999 3.3 0.00149268 0 0.0014926 0 0.0014927 3.3 0.0014926199999999998 3.3 0.00149272 0 0.00149264 0 0.00149274 3.3 0.0014926599999999998 3.3 0.0014927599999999999 0 0.00149268 0 0.00149278 3.3 0.0014927 3.3 0.0014928 0 0.00149272 0 0.00149282 3.3 0.00149274 3.3 0.00149284 0 0.0014927599999999999 0 0.00149286 3.3 0.00149278 3.3 0.00149288 0 0.0014927999999999999 0 0.0014929 3.3 0.00149282 3.3 0.00149292 0 0.0014928399999999998 0 0.00149294 3.3 0.00149286 3.3 0.00149296 0 0.0014928799999999998 0 0.0014929799999999999 3.3 0.0014929 3.3 0.001493 0 0.00149292 0 0.00149302 3.3 0.00149294 3.3 0.00149304 0 0.00149296 0 0.00149306 3.3 0.0014929799999999999 3.3 0.00149308 0 0.001493 0 0.0014931 3.3 0.0014930199999999999 3.3 0.00149312 0 0.00149304 0 0.00149314 3.3 0.0014930599999999998 3.3 0.0014931599999999999 0 0.00149308 0 0.00149318 3.3 0.0014930999999999998 3.3 0.0014931999999999999 0 0.00149312 0 0.00149322 3.3 0.00149314 3.3 0.00149324 0 0.0014931599999999999 0 0.00149326 3.3 0.00149318 3.3 0.00149328 0 0.0014931999999999999 0 0.0014933 3.3 0.00149322 3.3 0.00149332 0 0.0014932399999999998 0 0.00149334 3.3 0.00149326 3.3 0.00149336 0 0.0014932799999999998 0 0.0014933799999999999 3.3 0.0014933 3.3 0.0014934 0 0.00149332 0 0.00149342 3.3 0.00149334 3.3 0.00149344 0 0.00149336 0 0.00149346 3.3 0.0014933799999999999 3.3 0.00149348 0 0.0014934 0 0.0014935 3.3 0.0014934199999999999 3.3 0.00149352 0 0.00149344 0 0.00149354 3.3 0.0014934599999999998 3.3 0.00149356 0 0.00149348 0 0.00149358 3.3 0.0014934999999999998 3.3 0.0014935999999999999 0 0.00149352 0 0.00149362 3.3 0.00149354 3.3 0.00149364 0 0.00149356 0 0.00149366 3.3 0.00149358 3.3 0.00149368 0 0.0014935999999999999 0 0.0014937 3.3 0.00149362 3.3 0.00149372 0 0.0014936399999999999 0 0.00149374 3.3 0.00149366 3.3 0.00149376 0 0.0014936799999999998 0 0.0014937799999999999 3.3 0.0014937 3.3 0.0014938 0 0.0014937199999999998 0 0.0014938199999999999 3.3 0.00149374 3.3 0.00149384 0 0.00149376 0 0.00149386 3.3 0.0014937799999999999 3.3 0.00149388 0 0.0014938 0 0.0014939 3.3 0.0014938199999999999 3.3 0.00149392 0 0.00149384 0 0.00149394 3.3 0.0014938599999999998 3.3 0.00149396 0 0.00149388 0 0.00149398 3.3 0.0014938999999999998 3.3 0.0014939999999999999 0 0.00149392 0 0.00149402 3.3 0.0014939399999999998 3.3 0.0014940399999999999 0 0.00149396 0 0.00149406 3.3 0.00149398 3.3 0.00149408 0 0.0014939999999999999 0 0.0014941 3.3 0.00149402 3.3 0.00149412 0 0.0014940399999999999 0 0.00149414 3.3 0.00149406 3.3 0.00149416 0 0.0014940799999999998 0 0.00149418 3.3 0.0014941 3.3 0.0014942 0 0.0014941199999999998 0 0.0014942199999999999 3.3 0.00149414 3.3 0.00149424 0 0.00149416 0 0.00149426 3.3 0.00149418 3.3 0.00149428 0 0.0014942 0 0.0014943 3.3 0.0014942199999999999 3.3 0.00149432 0 0.00149424 0 0.00149434 3.3 0.0014942599999999999 3.3 0.00149436 0 0.00149428 0 0.00149438 3.3 0.0014942999999999998 3.3 0.0014944 0 0.00149432 0 0.00149442 3.3 0.0014943399999999998 3.3 0.0014944399999999999 0 0.00149436 0 0.00149446 3.3 0.00149438 3.3 0.00149448 0 0.0014944 0 0.0014945 3.3 0.00149442 3.3 0.00149452 0 0.0014944399999999999 0 0.00149454 3.3 0.00149446 3.3 0.00149456 0 0.0014944799999999999 0 0.00149458 3.3 0.0014945 3.3 0.0014946 0 0.0014945199999999998 0 0.0014946199999999999 3.3 0.00149454 3.3 0.00149464 0 0.0014945599999999998 0 0.0014946599999999999 3.3 0.00149458 3.3 0.00149468 0 0.0014946 0 0.0014947 3.3 0.0014946199999999999 3.3 0.00149472 0 0.00149464 0 0.00149474 3.3 0.0014946599999999999 3.3 0.00149476 0 0.00149468 0 0.00149478 3.3 0.0014946999999999998 3.3 0.0014948 0 0.00149472 0 0.00149482 3.3 0.0014947399999999998 3.3 0.0014948399999999999 0 0.00149476 0 0.00149486 3.3 0.0014947799999999998 3.3 0.0014948799999999999 0 0.0014948 0 0.0014949 3.3 0.00149482 3.3 0.00149492 0 0.0014948399999999999 0 0.00149494 3.3 0.00149486 3.3 0.00149496 0 0.0014948799999999999 0 0.00149498 3.3 0.0014949 3.3 0.001495 0 0.0014949199999999998 0 0.00149502 3.3 0.00149494 3.3 0.00149504 0 0.0014949599999999998 0 0.0014950599999999999 3.3 0.00149498 3.3 0.00149508 0 0.001495 0 0.0014951 3.3 0.00149502 3.3 0.00149512 0 0.00149504 0 0.00149514 3.3 0.0014950599999999999 3.3 0.00149516 0 0.00149508 0 0.00149518 3.3 0.0014950999999999999 3.3 0.0014952 0 0.00149512 0 0.00149522 3.3 0.0014951399999999998 3.3 0.00149524 0 0.00149516 0 0.00149526 3.3 0.0014951799999999998 3.3 0.0014952799999999999 0 0.0014952 0 0.0014953 3.3 0.00149522 3.3 0.00149532 0 0.00149524 0 0.00149534 3.3 0.00149526 3.3 0.00149536 0 0.0014952799999999999 0 0.00149538 3.3 0.0014953 3.3 0.0014954 0 0.0014953199999999999 0 0.00149542 3.3 0.00149534 3.3 0.00149544 0 0.0014953599999999998 0 0.0014954599999999999 3.3 0.00149538 3.3 0.00149548 0 0.0014953999999999998 0 0.0014954999999999999 3.3 0.00149542 3.3 0.00149552 0 0.00149544 0 0.00149554 3.3 0.0014954599999999999 3.3 0.00149556 0 0.00149548 0 0.00149558 3.3 0.0014954999999999999 3.3 0.0014956 0 0.00149552 0 0.00149562 3.3 0.0014955399999999998 3.3 0.00149564 0 0.00149556 0 0.00149566 3.3 0.0014955799999999998 3.3 0.0014956799999999999 0 0.0014956 0 0.0014957 3.3 0.0014956199999999998 3.3 0.0014957199999999999 0 0.00149564 0 0.00149574 3.3 0.00149566 3.3 0.00149576 0 0.0014956799999999999 0 0.00149578 3.3 0.0014957 3.3 0.0014958 0 0.0014957199999999999 0 0.00149582 3.3 0.00149574 3.3 0.00149584 0 0.0014957599999999998 0 0.00149586 3.3 0.00149578 3.3 0.00149588 0 0.0014957999999999998 0 0.0014958999999999999 3.3 0.00149582 3.3 0.00149592 0 0.00149584 0 0.00149594 3.3 0.00149586 3.3 0.00149596 0 0.00149588 0 0.00149598 3.3 0.0014958999999999999 3.3 0.001496 0 0.00149592 0 0.00149602 3.3 0.0014959399999999999 3.3 0.00149604 0 0.00149596 0 0.00149606 3.3 0.0014959799999999998 3.3 0.00149608 0 0.001496 0 0.0014961 3.3 0.0014960199999999998 3.3 0.0014961199999999999 0 0.00149604 0 0.00149614 3.3 0.00149606 3.3 0.00149616 0 0.00149608 0 0.00149618 3.3 0.0014961 3.3 0.0014962 0 0.0014961199999999999 0 0.00149622 3.3 0.00149614 3.3 0.00149624 0 0.0014961599999999999 0 0.00149626 3.3 0.00149618 3.3 0.00149628 0 0.0014961999999999998 0 0.0014962999999999999 3.3 0.00149622 3.3 0.00149632 0 0.0014962399999999998 0 0.0014963399999999999 3.3 0.00149626 3.3 0.00149636 0 0.00149628 0 0.00149638 3.3 0.0014962999999999999 3.3 0.0014964 0 0.00149632 0 0.00149642 3.3 0.0014963399999999999 3.3 0.00149644 0 0.00149636 0 0.00149646 3.3 0.0014963799999999998 3.3 0.00149648 0 0.0014964 0 0.0014965 3.3 0.0014964199999999998 3.3 0.0014965199999999999 0 0.00149644 0 0.00149654 3.3 0.00149646 3.3 0.00149656 0 0.00149648 0 0.00149658 3.3 0.0014965 3.3 0.0014966 0 0.0014965199999999999 0 0.00149662 3.3 0.00149654 3.3 0.00149664 0 0.0014965599999999999 0 0.00149666 3.3 0.00149658 3.3 0.00149668 0 0.0014965999999999998 0 0.0014967 3.3 0.00149662 3.3 0.00149672 0 0.0014966399999999998 0 0.0014967399999999999 3.3 0.00149666 3.3 0.00149676 0 0.00149668 0 0.00149678 3.3 0.0014967 3.3 0.0014968 0 0.00149672 0 0.00149682 3.3 0.0014967399999999999 3.3 0.00149684 0 0.00149676 0 0.00149686 3.3 0.0014967799999999999 3.3 0.00149688 0 0.0014968 0 0.0014969 3.3 0.0014968199999999998 3.3 0.0014969199999999999 0 0.00149684 0 0.00149694 3.3 0.0014968599999999998 3.3 0.0014969599999999999 0 0.00149688 0 0.00149698 3.3 0.0014969 3.3 0.001497 0 0.0014969199999999999 0 0.00149702 3.3 0.00149694 3.3 0.00149704 0 0.0014969599999999999 0 0.00149706 3.3 0.00149698 3.3 0.00149708 0 0.0014969999999999998 0 0.0014971 3.3 0.00149702 3.3 0.00149712 0 0.0014970399999999998 0 0.0014971399999999999 3.3 0.00149706 3.3 0.00149716 0 0.0014970799999999998 0 0.0014971799999999999 3.3 0.0014971 3.3 0.0014972 0 0.00149712 0 0.00149722 3.3 0.0014971399999999999 3.3 0.00149724 0 0.00149716 0 0.00149726 3.3 0.0014971799999999999 3.3 0.00149728 0 0.0014972 0 0.0014973 3.3 0.0014972199999999998 3.3 0.00149732 0 0.00149724 0 0.00149734 3.3 0.0014972599999999998 3.3 0.0014973599999999999 0 0.00149728 0 0.00149738 3.3 0.0014973 3.3 0.0014974 0 0.00149732 0 0.00149742 3.3 0.00149734 3.3 0.00149744 0 0.0014973599999999999 0 0.00149746 3.3 0.00149738 3.3 0.00149748 0 0.0014973999999999999 0 0.0014975 3.3 0.00149742 3.3 0.00149752 0 0.0014974399999999998 0 0.00149754 3.3 0.00149746 3.3 0.00149756 0 0.0014974799999999998 0 0.0014975799999999999 3.3 0.0014975 3.3 0.0014976 0 0.00149752 0 0.00149762 3.3 0.00149754 3.3 0.00149764 0 0.00149756 0 0.00149766 3.3 0.0014975799999999999 3.3 0.00149768 0 0.0014976 0 0.0014977 3.3 0.0014976199999999999 3.3 0.00149772 0 0.00149764 0 0.00149774 3.3 0.0014976599999999998 3.3 0.0014977599999999999 0 0.00149768 0 0.00149778 3.3 0.0014976999999999998 3.3 0.0014977999999999999 0 0.00149772 0 0.00149782 3.3 0.00149774 3.3 0.00149784 0 0.0014977599999999999 0 0.00149786 3.3 0.00149778 3.3 0.00149788 0 0.0014977999999999999 0 0.0014979 3.3 0.00149782 3.3 0.00149792 0 0.0014978399999999998 0 0.00149794 3.3 0.00149786 3.3 0.00149796 0 0.0014978799999999998 0 0.0014979799999999999 3.3 0.0014979 3.3 0.001498 0 0.0014979199999999998 0 0.0014980199999999999 3.3 0.00149794 3.3 0.00149804 0 0.00149796 0 0.00149806 3.3 0.0014979799999999999 3.3 0.00149808 0 0.001498 0 0.0014981 3.3 0.0014980199999999999 3.3 0.00149812 0 0.00149804 0 0.00149814 3.3 0.0014980599999999998 3.3 0.00149816 0 0.00149808 0 0.00149818 3.3 0.0014980999999999998 3.3 0.0014981999999999999 0 0.00149812 0 0.00149822 3.3 0.00149814 3.3 0.00149824 0 0.00149816 0 0.00149826 3.3 0.00149818 3.3 0.00149828 0 0.0014981999999999999 0 0.0014983 3.3 0.00149822 3.3 0.00149832 0 0.0014982399999999999 0 0.00149834 3.3 0.00149826 3.3 0.00149836 0 0.0014982799999999998 0 0.00149838 3.3 0.0014983 3.3 0.0014984 0 0.0014983199999999998 0 0.0014984199999999999 3.3 0.00149834 3.3 0.00149844 0 0.00149836 0 0.00149846 3.3 0.00149838 3.3 0.00149848 0 0.0014984 0 0.0014985 3.3 0.0014984199999999999 3.3 0.00149852 0 0.00149844 0 0.00149854 3.3 0.0014984599999999999 3.3 0.00149856 0 0.00149848 0 0.00149858 3.3 0.0014984999999999998 3.3 0.0014985999999999999 0 0.00149852 0 0.00149862 3.3 0.0014985399999999998 3.3 0.0014986399999999999 0 0.00149856 0 0.00149866 3.3 0.00149858 3.3 0.00149868 0 0.0014985999999999999 0 0.0014987 3.3 0.00149862 3.3 0.00149872 0 0.0014986399999999999 0 0.00149874 3.3 0.00149866 3.3 0.00149876 0 0.0014986799999999998 0 0.00149878 3.3 0.0014987 3.3 0.0014988 0 0.0014987199999999998 0 0.0014988199999999999 3.3 0.00149874 3.3 0.00149884 0 0.0014987599999999998 0 0.0014988599999999999 3.3 0.00149878 3.3 0.00149888 0 0.0014988 0 0.0014989 3.3 0.0014988199999999999 3.3 0.00149892 0 0.00149884 0 0.00149894 3.3 0.0014988599999999999 3.3 0.00149896 0 0.00149888 0 0.00149898 3.3 0.0014988999999999998 3.3 0.001499 0 0.00149892 0 0.00149902 3.3 0.0014989399999999998 3.3 0.0014990399999999999 0 0.00149896 0 0.00149906 3.3 0.00149898 3.3 0.00149908 0 0.001499 0 0.0014991 3.3 0.00149902 3.3 0.00149912 0 0.0014990399999999999 0 0.00149914 3.3 0.00149906 3.3 0.00149916 0 0.0014990799999999999 0 0.00149918 3.3 0.0014991 3.3 0.0014992 0 0.0014991199999999998 0 0.00149922 3.3 0.00149914 3.3 0.00149924 0 0.0014991599999999998 0 0.0014992599999999999 3.3 0.00149918 3.3 0.00149928 0 0.0014992 0 0.0014993 3.3 0.00149922 3.3 0.00149932 0 0.00149924 0 0.00149934 3.3 0.0014992599999999999 3.3 0.00149936 0 0.00149928 0 0.00149938 3.3 0.0014992999999999999 3.3 0.0014994 0 0.00149932 0 0.00149942 3.3 0.0014993399999999998 3.3 0.0014994399999999999 0 0.00149936 0 0.00149946 3.3 0.0014993799999999998 3.3 0.0014994799999999999 0 0.0014994 0 0.0014995 3.3 0.00149942 3.3 0.00149952 0 0.0014994399999999999 0 0.00149954 3.3 0.00149946 3.3 0.00149956 0 0.0014994799999999999 0 0.00149958 3.3 0.0014995 3.3 0.0014996 0 0.0014995199999999998 0 0.00149962 3.3 0.00149954 3.3 0.00149964 0 0.0014995599999999998 0 0.0014996599999999999 3.3 0.00149958 3.3 0.00149968 0 0.0014996 0 0.0014997 3.3 0.00149962 3.3 0.00149972 0 0.00149964 0 0.00149974 3.3 0.0014996599999999999 3.3 0.00149976 0 0.00149968 0 0.00149978 3.3 0.0014996999999999999 3.3 0.0014998 0 0.00149972 0 0.00149982 3.3 0.0014997399999999998 3.3 0.00149984 0 0.00149976 0 0.00149986 3.3 0.0014997799999999998 3.3 0.0014998799999999999 0 0.0014998 0 0.0014999 3.3 0.00149982 3.3 0.00149992 0 0.00149984 0 0.00149994 3.3 0.00149986 3.3 0.00149996 0 0.0014998799999999999 0 0.00149998 3.3 0.0014999 3.3 0.0015 0 0.0014999199999999999 0 0.00150002 3.3 0.00149994 3.3 0.00150004 0 0.0014999599999999998 0 0.00150006 3.3 0.00149998 3.3 0.00150008 0 0.0014999999999999998 0 0.0015000999999999999 3.3 0.00150002 3.3 0.00150012 0 0.00150004 0 0.00150014 3.3 0.00150006 3.3 0.00150016 0 0.00150008 0 0.00150018 3.3 0.0015000999999999999 3.3 0.0015002 0 0.00150012 0 0.00150022 3.3 0.0015001399999999999 3.3 0.00150024 0 0.00150016 0 0.00150026 3.3 0.0015001799999999998 3.3 0.0015002799999999999 0 0.0015002 0 0.0015003 3.3 0.0015002199999999998 3.3 0.0015003199999999999 0 0.00150024 0 0.00150034 3.3 0.00150026 3.3 0.00150036 0 0.0015002799999999999 0 0.00150038 3.3 0.0015003 3.3 0.0015004 0 0.0015003199999999999 0 0.00150042 3.3 0.00150034 3.3 0.00150044 0 0.0015003599999999998 0 0.00150046 3.3 0.00150038 3.3 0.00150048 0 0.0015003999999999998 0 0.0015004999999999999 3.3 0.00150042 3.3 0.00150052 0 0.00150044 0 0.00150054 3.3 0.00150046 3.3 0.00150056 0 0.00150048 0 0.00150058 3.3 0.0015004999999999999 3.3 0.0015006 0 0.00150052 0 0.00150062 3.3 0.0015005399999999999 3.3 0.00150064 0 0.00150056 0 0.00150066 3.3 0.0015005799999999998 3.3 0.00150068 0 0.0015006 0 0.0015007 3.3 0.0015006199999999998 3.3 0.0015007199999999999 0 0.00150064 0 0.00150074 3.3 0.00150066 3.3 0.00150076 0 0.00150068 0 0.00150078 3.3 0.0015007 3.3 0.0015008 0 0.0015007199999999999 0 0.00150082 3.3 0.00150074 3.3 0.00150084 0 0.0015007599999999999 0 0.00150086 3.3 0.00150078 3.3 0.00150088 0 0.0015007999999999998 0 0.0015008999999999999 3.3 0.00150082 3.3 0.00150092 0 0.0015008399999999998 0 0.0015009399999999999 3.3 0.00150086 3.3 0.00150096 0 0.00150088 0 0.00150098 3.3 0.0015008999999999999 3.3 0.001501 0 0.00150092 0 0.00150102 3.3 0.0015009399999999999 3.3 0.00150104 0 0.00150096 0 0.00150106 3.3 0.0015009799999999998 3.3 0.00150108 0 0.001501 0 0.0015011 3.3 0.0015010199999999998 3.3 0.0015011199999999999 0 0.00150104 0 0.00150114 3.3 0.0015010599999999998 3.3 0.0015011599999999999 0 0.00150108 0 0.00150118 3.3 0.0015011 3.3 0.0015012 0 0.0015011199999999999 0 0.00150122 3.3 0.00150114 3.3 0.00150124 0 0.0015011599999999999 0 0.00150126 3.3 0.00150118 3.3 0.00150128 0 0.0015011999999999998 0 0.0015013 3.3 0.00150122 3.3 0.00150132 0 0.0015012399999999998 0 0.0015013399999999999 3.3 0.00150126 3.3 0.00150136 0 0.00150128 0 0.00150138 3.3 0.0015013 3.3 0.0015014 0 0.00150132 0 0.00150142 3.3 0.0015013399999999999 3.3 0.00150144 0 0.00150136 0 0.00150146 3.3 0.0015013799999999999 3.3 0.00150148 0 0.0015014 0 0.0015015 3.3 0.0015014199999999998 3.3 0.00150152 0 0.00150144 0 0.00150154 3.3 0.0015014599999999998 3.3 0.0015015599999999999 0 0.00150148 0 0.00150158 3.3 0.0015015 3.3 0.0015016 0 0.00150152 0 0.00150162 3.3 0.00150154 3.3 0.00150164 0 0.0015015599999999999 0 0.00150166 3.3 0.00150158 3.3 0.00150168 0 0.0015015999999999999 0 0.0015017 3.3 0.00150162 3.3 0.00150172 0 0.0015016399999999998 0 0.0015017399999999999 3.3 0.00150166 3.3 0.00150176 0 0.0015016799999999998 0 0.0015017799999999999 3.3 0.0015017 3.3 0.0015018 0 0.00150172 0 0.00150182 3.3 0.0015017399999999999 3.3 0.00150184 0 0.00150176 0 0.00150186 3.3 0.0015017799999999999 3.3 0.00150188 0 0.0015018 0 0.0015019 3.3 0.0015018199999999998 3.3 0.00150192 0 0.00150184 0 0.00150194 3.3 0.0015018599999999998 3.3 0.0015019599999999999 0 0.00150188 0 0.00150198 3.3 0.0015018999999999998 3.3 0.0015019999999999999 0 0.00150192 0 0.00150202 3.3 0.00150194 3.3 0.00150204 0 0.0015019599999999999 0 0.00150206 3.3 0.00150198 3.3 0.00150208 0 0.0015019999999999999 0 0.0015021 3.3 0.00150202 3.3 0.00150212 0 0.0015020399999999998 0 0.00150214 3.3 0.00150206 3.3 0.00150216 0 0.0015020799999999998 0 0.0015021799999999999 3.3 0.0015021 3.3 0.0015022 0 0.00150212 0 0.00150222 3.3 0.00150214 3.3 0.00150224 0 0.00150216 0 0.00150226 3.3 0.0015021799999999999 3.3 0.00150228 0 0.0015022 0 0.0015023 3.3 0.0015022199999999999 3.3 0.00150232 0 0.00150224 0 0.00150234 3.3 0.0015022599999999998 3.3 0.00150236 0 0.00150228 0 0.00150238 3.3 0.0015022999999999998 3.3 0.0015023999999999999 0 0.00150232 0 0.00150242 3.3 0.00150234 3.3 0.00150244 0 0.00150236 0 0.00150246 3.3 0.00150238 3.3 0.00150248 0 0.0015023999999999999 0 0.0015025 3.3 0.00150242 3.3 0.00150252 0 0.0015024399999999999 0 0.00150254 3.3 0.00150246 3.3 0.00150256 0 0.0015024799999999998 0 0.0015025799999999999 3.3 0.0015025 3.3 0.0015026 0 0.0015025199999999998 0 0.0015026199999999999 3.3 0.00150254 3.3 0.00150264 0 0.00150256 0 0.00150266 3.3 0.0015025799999999999 3.3 0.00150268 0 0.0015026 0 0.0015027 3.3 0.0015026199999999999 3.3 0.00150272 0 0.00150264 0 0.00150274 3.3 0.0015026599999999998 3.3 0.00150276 0 0.00150268 0 0.00150278 3.3 0.0015026999999999998 3.3 0.0015027999999999999 0 0.00150272 0 0.00150282 3.3 0.0015027399999999998 3.3 0.0015028399999999999 0 0.00150276 0 0.00150286 3.3 0.00150278 3.3 0.00150288 0 0.0015027999999999999 0 0.0015029 3.3 0.00150282 3.3 0.00150292 0 0.0015028399999999999 0 0.00150294 3.3 0.00150286 3.3 0.00150296 0 0.0015028799999999998 0 0.00150298 3.3 0.0015029 3.3 0.001503 0 0.0015029199999999998 0 0.0015030199999999999 3.3 0.00150294 3.3 0.00150304 0 0.00150296 0 0.00150306 3.3 0.00150298 3.3 0.00150308 0 0.001503 0 0.0015031 3.3 0.0015030199999999999 3.3 0.00150312 0 0.00150304 0 0.00150314 3.3 0.0015030599999999999 3.3 0.00150316 0 0.00150308 0 0.00150318 3.3 0.0015030999999999998 3.3 0.0015032 0 0.00150312 0 0.00150322 3.3 0.0015031399999999998 3.3 0.0015032399999999999 0 0.00150316 0 0.00150326 3.3 0.00150318 3.3 0.00150328 0 0.0015032 0 0.0015033 3.3 0.00150322 3.3 0.00150332 0 0.0015032399999999999 0 0.00150334 3.3 0.00150326 3.3 0.00150336 0 0.0015032799999999999 0 0.00150338 3.3 0.0015033 3.3 0.0015034 0 0.0015033199999999998 0 0.0015034199999999999 3.3 0.00150334 3.3 0.00150344 0 0.0015033599999999998 0 0.0015034599999999999 3.3 0.00150338 3.3 0.00150348 0 0.0015034 0 0.0015035 3.3 0.0015034199999999999 3.3 0.00150352 0 0.00150344 0 0.00150354 3.3 0.0015034599999999999 3.3 0.00150356 0 0.00150348 0 0.00150358 3.3 0.0015034999999999998 3.3 0.0015036 0 0.00150352 0 0.00150362 3.3 0.0015035399999999998 3.3 0.0015036399999999999 0 0.00150356 0 0.00150366 3.3 0.00150358 3.3 0.00150368 0 0.0015036 0 0.0015037 3.3 0.00150362 3.3 0.00150372 0 0.0015036399999999999 0 0.00150374 3.3 0.00150366 3.3 0.00150376 0 0.0015036799999999999 0 0.00150378 3.3 0.0015037 3.3 0.0015038 0 0.0015037199999999998 0 0.00150382 3.3 0.00150374 3.3 0.00150384 0 0.0015037599999999998 0 0.0015038599999999999 3.3 0.00150378 3.3 0.00150388 0 0.0015038 0 0.0015039 3.3 0.00150382 3.3 0.00150392 0 0.00150384 0 0.00150394 3.3 0.0015038599999999999 3.3 0.00150396 0 0.00150388 0 0.00150398 3.3 0.0015038999999999999 3.3 0.001504 0 0.00150392 0 0.00150402 3.3 0.0015039399999999998 3.3 0.0015040399999999999 0 0.00150396 0 0.00150406 3.3 0.0015039799999999998 3.3 0.0015040799999999999 0 0.001504 0 0.0015041 3.3 0.00150402 3.3 0.00150412 0 0.0015040399999999999 0 0.00150414 3.3 0.00150406 3.3 0.00150416 0 0.0015040799999999999 0 0.00150418 3.3 0.0015041 3.3 0.0015042 0 0.0015041199999999998 0 0.00150422 3.3 0.00150414 3.3 0.00150424 0 0.0015041599999999998 0 0.0015042599999999999 3.3 0.00150418 3.3 0.00150428 0 0.0015041999999999998 0 0.0015042999999999999 3.3 0.00150422 3.3 0.00150432 0 0.00150424 0 0.00150434 3.3 0.0015042599999999999 3.3 0.00150436 0 0.00150428 0 0.00150438 3.3 0.0015042999999999999 3.3 0.0015044 0 0.00150432 0 0.00150442 3.3 0.0015043399999999998 3.3 0.00150444 0 0.00150436 0 0.00150446 3.3 0.0015043799999999998 3.3 0.0015044799999999999 0 0.0015044 0 0.0015045 3.3 0.00150442 3.3 0.00150452 0 0.00150444 0 0.00150454 3.3 0.00150446 3.3 0.00150456 0 0.0015044799999999999 0 0.00150458 3.3 0.0015045 3.3 0.0015046 0 0.0015045199999999999 0 0.00150462 3.3 0.00150454 3.3 0.00150464 0 0.0015045599999999998 0 0.00150466 3.3 0.00150458 3.3 0.00150468 0 0.0015045999999999998 0 0.0015046999999999999 3.3 0.00150462 3.3 0.00150472 0 0.00150464 0 0.00150474 3.3 0.00150466 3.3 0.00150476 0 0.00150468 0 0.00150478 3.3 0.0015046999999999999 3.3 0.0015048 0 0.00150472 0 0.00150482 3.3 0.0015047399999999999 3.3 0.00150484 0 0.00150476 0 0.00150486 3.3 0.0015047799999999998 3.3 0.0015048799999999999 0 0.0015048 0 0.0015049 3.3 0.0015048199999999998 3.3 0.0015049199999999999 0 0.00150484 0 0.00150494 3.3 0.00150486 3.3 0.00150496 0 0.0015048799999999999 0 0.00150498 3.3 0.0015049 3.3 0.001505 0 0.0015049199999999999 0 0.00150502 3.3 0.00150494 3.3 0.00150504 0 0.0015049599999999998 0 0.00150506 3.3 0.00150498 3.3 0.00150508 0 0.0015049999999999998 0 0.0015050999999999999 3.3 0.00150502 3.3 0.00150512 0 0.0015050399999999998 0 0.0015051399999999999 3.3 0.00150506 3.3 0.00150516 0 0.00150508 0 0.00150518 3.3 0.0015050999999999999 3.3 0.0015052 0 0.00150512 0 0.00150522 3.3 0.0015051399999999999 3.3 0.00150524 0 0.00150516 0 0.00150526 3.3 0.0015051799999999998 3.3 0.00150528 0 0.0015052 0 0.0015053 3.3 0.0015052199999999998 3.3 0.0015053199999999999 0 0.00150524 0 0.00150534 3.3 0.00150526 3.3 0.00150536 0 0.00150528 0 0.00150538 3.3 0.0015053 3.3 0.0015054 0 0.0015053199999999999 0 0.00150542 3.3 0.00150534 3.3 0.00150544 0 0.0015053599999999999 0 0.00150546 3.3 0.00150538 3.3 0.00150548 0 0.0015053999999999998 0 0.0015055 3.3 0.00150542 3.3 0.00150552 0 0.0015054399999999998 0 0.0015055399999999999 3.3 0.00150546 3.3 0.00150556 0 0.00150548 0 0.00150558 3.3 0.0015055 3.3 0.0015056 0 0.00150552 0 0.00150562 3.3 0.0015055399999999999 3.3 0.00150564 0 0.00150556 0 0.00150566 3.3 0.0015055799999999999 3.3 0.00150568 0 0.0015056 0 0.0015057 3.3 0.0015056199999999998 3.3 0.0015057199999999999 0 0.00150564 0 0.00150574 3.3 0.0015056599999999998 3.3 0.0015057599999999999 0 0.00150568 0 0.00150578 3.3 0.0015057 3.3 0.0015058 0 0.0015057199999999999 0 0.00150582 3.3 0.00150574 3.3 0.00150584 0 0.0015057599999999999 0 0.00150586 3.3 0.00150578 3.3 0.00150588 0 0.0015057999999999998 0 0.0015059 3.3 0.00150582 3.3 0.00150592 0 0.0015058399999999998 0 0.0015059399999999999 3.3 0.00150586 3.3 0.00150596 0 0.0015058799999999998 0 0.0015059799999999999 3.3 0.0015059 3.3 0.001506 0 0.00150592 0 0.00150602 3.3 0.0015059399999999999 3.3 0.00150604 0 0.00150596 0 0.00150606 3.3 0.0015059799999999999 3.3 0.00150608 0 0.001506 0 0.0015061 3.3 0.0015060199999999998 3.3 0.00150612 0 0.00150604 0 0.00150614 3.3 0.0015060599999999998 3.3 0.0015061599999999999 0 0.00150608 0 0.00150618 3.3 0.0015061 3.3 0.0015062 0 0.00150612 0 0.00150622 3.3 0.00150614 3.3 0.00150624 0 0.0015061599999999999 0 0.00150626 3.3 0.00150618 3.3 0.00150628 0 0.0015061999999999999 0 0.0015063 3.3 0.00150622 3.3 0.00150632 0 0.0015062399999999998 0 0.00150634 3.3 0.00150626 3.3 0.00150636 0 0.0015062799999999998 0 0.0015063799999999999 3.3 0.0015063 3.3 0.0015064 0 0.00150632 0 0.00150642 3.3 0.00150634 3.3 0.00150644 0 0.00150636 0 0.00150646 3.3 0.0015063799999999999 3.3 0.00150648 0 0.0015064 0 0.0015065 3.3 0.0015064199999999999 3.3 0.00150652 0 0.00150644 0 0.00150654 3.3 0.0015064599999999998 3.3 0.0015065599999999999 0 0.00150648 0 0.00150658 3.3 0.0015064999999999998 3.3 0.0015065999999999999 0 0.00150652 0 0.00150662 3.3 0.00150654 3.3 0.00150664 0 0.0015065599999999999 0 0.00150666 3.3 0.00150658 3.3 0.00150668 0 0.0015065999999999999 0 0.0015067 3.3 0.00150662 3.3 0.00150672 0 0.0015066399999999998 0 0.00150674 3.3 0.00150666 3.3 0.00150676 0 0.0015066799999999998 0 0.0015067799999999999 3.3 0.0015067 3.3 0.0015068 0 0.00150672 0 0.00150682 3.3 0.00150674 3.3 0.00150684 0 0.00150676 0 0.00150686 3.3 0.0015067799999999999 3.3 0.00150688 0 0.0015068 0 0.0015069 3.3 0.0015068199999999999 3.3 0.00150692 0 0.00150684 0 0.00150694 3.3 0.0015068599999999998 3.3 0.00150696 0 0.00150688 0 0.00150698 3.3 0.0015068999999999998 3.3 0.0015069999999999999 0 0.00150692 0 0.00150702 3.3 0.00150694 3.3 0.00150704 0 0.00150696 0 0.00150706 3.3 0.00150698 3.3 0.00150708 0 0.0015069999999999999 0 0.0015071 3.3 0.00150702 3.3 0.00150712 0 0.0015070399999999999 0 0.00150714 3.3 0.00150706 3.3 0.00150716 0 0.0015070799999999998 0 0.0015071799999999999 3.3 0.0015071 3.3 0.0015072 0 0.0015071199999999998 0 0.0015072199999999999 3.3 0.00150714 3.3 0.00150724 0 0.00150716 0 0.00150726 3.3 0.0015071799999999999 3.3 0.00150728 0 0.0015072 0 0.0015073 3.3 0.0015072199999999999 3.3 0.00150732 0 0.00150724 0 0.00150734 3.3 0.0015072599999999998 3.3 0.00150736 0 0.00150728 0 0.00150738 3.3 0.0015072999999999998 3.3 0.0015073999999999999 0 0.00150732 0 0.00150742 3.3 0.0015073399999999998 3.3 0.0015074399999999999 0 0.00150736 0 0.00150746 3.3 0.00150738 3.3 0.00150748 0 0.0015073999999999999 0 0.0015075 3.3 0.00150742 3.3 0.00150752 0 0.0015074399999999999 0 0.00150754 3.3 0.00150746 3.3 0.00150756 0 0.0015074799999999998 0 0.00150758 3.3 0.0015075 3.3 0.0015076 0 0.0015075199999999998 0 0.0015076199999999999 3.3 0.00150754 3.3 0.00150764 0 0.00150756 0 0.00150766 3.3 0.00150758 3.3 0.00150768 0 0.0015076 0 0.0015077 3.3 0.0015076199999999999 3.3 0.00150772 0 0.00150764 0 0.00150774 3.3 0.0015076599999999999 3.3 0.00150776 0 0.00150768 0 0.00150778 3.3 0.0015076999999999998 3.3 0.0015078 0 0.00150772 0 0.00150782 3.3 0.0015077399999999998 3.3 0.0015078399999999999 0 0.00150776 0 0.00150786 3.3 0.00150778 3.3 0.00150788 0 0.0015078 0 0.0015079 3.3 0.00150782 3.3 0.00150792 0 0.0015078399999999999 0 0.00150794 3.3 0.00150786 3.3 0.00150796 0 0.0015078799999999999 0 0.00150798 3.3 0.0015079 3.3 0.001508 0 0.0015079199999999998 0 0.0015080199999999999 3.3 0.00150794 3.3 0.00150804 0 0.0015079599999999998 0 0.0015080599999999999 3.3 0.00150798 3.3 0.00150808 0 0.001508 0 0.0015081 3.3 0.0015080199999999999 3.3 0.00150812 0 0.00150804 0 0.00150814 3.3 0.0015080599999999999 3.3 0.00150816 0 0.00150808 0 0.00150818 3.3 0.0015080999999999998 3.3 0.0015082 0 0.00150812 0 0.00150822 3.3 0.0015081399999999998 3.3 0.0015082399999999999 0 0.00150816 0 0.00150826 3.3 0.0015081799999999998 3.3 0.0015082799999999999 0 0.0015082 0 0.0015083 3.3 0.00150822 3.3 0.00150832 0 0.0015082399999999999 0 0.00150834 3.3 0.00150826 3.3 0.00150836 0 0.0015082799999999999 0 0.00150838 3.3 0.0015083 3.3 0.0015084 0 0.0015083199999999998 0 0.00150842 3.3 0.00150834 3.3 0.00150844 0 0.0015083599999999998 0 0.0015084599999999999 3.3 0.00150838 3.3 0.00150848 0 0.0015084 0 0.0015085 3.3 0.00150842 3.3 0.00150852 0 0.00150844 0 0.00150854 3.3 0.0015084599999999999 3.3 0.00150856 0 0.00150848 0 0.00150858 3.3 0.0015084999999999999 3.3 0.0015086 0 0.00150852 0 0.00150862 3.3 0.0015085399999999998 3.3 0.00150864 0 0.00150856 0 0.00150866 3.3 0.0015085799999999998 3.3 0.0015086799999999999 0 0.0015086 0 0.0015087 3.3 0.00150862 3.3 0.00150872 0 0.00150864 0 0.00150874 3.3 0.00150866 3.3 0.00150876 0 0.0015086799999999999 0 0.00150878 3.3 0.0015087 3.3 0.0015088 0 0.0015087199999999999 0 0.00150882 3.3 0.00150874 3.3 0.00150884 0 0.0015087599999999998 0 0.0015088599999999999 3.3 0.00150878 3.3 0.00150888 0 0.0015087999999999998 0 0.0015088999999999999 3.3 0.00150882 3.3 0.00150892 0 0.00150884 0 0.00150894 3.3 0.0015088599999999999 3.3 0.00150896 0 0.00150888 0 0.00150898 3.3 0.0015088999999999999 3.3 0.001509 0 0.00150892 0 0.00150902 3.3 0.0015089399999999998 3.3 0.00150904 0 0.00150896 0 0.00150906 3.3 0.0015089799999999998 3.3 0.0015090799999999999 0 0.001509 0 0.0015091 3.3 0.0015090199999999998 3.3 0.0015091199999999999 0 0.00150904 0 0.00150914 3.3 0.00150906 3.3 0.00150916 0 0.0015090799999999999 0 0.00150918 3.3 0.0015091 3.3 0.0015092 0 0.0015091199999999999 0 0.00150922 3.3 0.00150914 3.3 0.00150924 0 0.0015091599999999998 0 0.00150926 3.3 0.00150918 3.3 0.00150928 0 0.0015091999999999998 0 0.0015092999999999999 3.3 0.00150922 3.3 0.00150932 0 0.00150924 0 0.00150934 3.3 0.00150926 3.3 0.00150936 0 0.00150928 0 0.00150938 3.3 0.0015092999999999999 3.3 0.0015094 0 0.00150932 0 0.00150942 3.3 0.0015093399999999999 3.3 0.00150944 0 0.00150936 0 0.00150946 3.3 0.0015093799999999998 3.3 0.00150948 0 0.0015094 0 0.0015095 3.3 0.0015094199999999998 3.3 0.0015095199999999999 0 0.00150944 0 0.00150954 3.3 0.00150946 3.3 0.00150956 0 0.00150948 0 0.00150958 3.3 0.0015095 3.3 0.0015096 0 0.0015095199999999999 0 0.00150962 3.3 0.00150954 3.3 0.00150964 0 0.0015095599999999999 0 0.00150966 3.3 0.00150958 3.3 0.00150968 0 0.0015095999999999998 0 0.0015096999999999999 3.3 0.00150962 3.3 0.00150972 0 0.0015096399999999998 0 0.0015097399999999999 3.3 0.00150966 3.3 0.00150976 0 0.00150968 0 0.00150978 3.3 0.0015096999999999999 3.3 0.0015098 0 0.00150972 0 0.00150982 3.3 0.0015097399999999999 3.3 0.00150984 0 0.00150976 0 0.00150986 3.3 0.0015097799999999998 3.3 0.00150988 0 0.0015098 0 0.0015099 3.3 0.0015098199999999998 3.3 0.0015099199999999999 0 0.00150984 0 0.00150994 3.3 0.0015098599999999998 3.3 0.0015099599999999999 0 0.00150988 0 0.00150998 3.3 0.0015099 3.3 0.00151 0 0.0015099199999999999 0 0.00151002 3.3 0.00150994 3.3 0.00151004 0 0.0015099599999999999 0 0.00151006 3.3 0.00150998 3.3 0.00151008 0 0.0015099999999999998 0 0.0015101 3.3 0.00151002 3.3 0.00151012 0 0.0015100399999999998 0 0.0015101399999999999 3.3 0.00151006 3.3 0.00151016 0 0.00151008 0 0.00151018 3.3 0.0015101 3.3 0.0015102 0 0.00151012 0 0.00151022 3.3 0.0015101399999999999 3.3 0.00151024 0 0.00151016 0 0.00151026 3.3 0.0015101799999999999 3.3 0.00151028 0 0.0015102 0 0.0015103 3.3 0.0015102199999999998 3.3 0.00151032 0 0.00151024 0 0.00151034 3.3 0.0015102599999999998 3.3 0.0015103599999999999 0 0.00151028 0 0.00151038 3.3 0.0015103 3.3 0.0015104 0 0.00151032 0 0.00151042 3.3 0.00151034 3.3 0.00151044 0 0.0015103599999999999 0 0.00151046 3.3 0.00151038 3.3 0.00151048 0 0.0015103999999999999 0 0.0015105 3.3 0.00151042 3.3 0.00151052 0 0.0015104399999999998 0 0.0015105399999999999 3.3 0.00151046 3.3 0.00151056 0 0.0015104799999999998 0 0.0015105799999999999 3.3 0.0015105 3.3 0.0015106 0 0.00151052 0 0.00151062 3.3 0.0015105399999999999 3.3 0.00151064 0 0.00151056 0 0.00151066 3.3 0.0015105799999999999 3.3 0.00151068 0 0.0015106 0 0.0015107 3.3 0.0015106199999999998 3.3 0.00151072 0 0.00151064 0 0.00151074 3.3 0.0015106599999999998 3.3 0.0015107599999999999 0 0.00151068 0 0.00151078 3.3 0.0015107 3.3 0.0015108 0 0.00151072 0 0.00151082 3.3 0.00151074 3.3 0.00151084 0 0.0015107599999999999 0 0.00151086 3.3 0.00151078 3.3 0.00151088 0 0.0015107999999999999 0 0.0015109 3.3 0.00151082 3.3 0.00151092 0 0.0015108399999999998 0 0.00151094 3.3 0.00151086 3.3 0.00151096 0 0.0015108799999999998 0 0.0015109799999999999 3.3 0.0015109 3.3 0.001511 0 0.00151092 0 0.00151102 3.3 0.00151094 3.3 0.00151104 0 0.00151096 0 0.00151106 3.3 0.0015109799999999999 3.3 0.00151108 0 0.001511 0 0.0015111 3.3 0.0015110199999999999 3.3 0.00151112 0 0.00151104 0 0.00151114 3.3 0.0015110599999999998 3.3 0.0015111599999999999 0 0.00151108 0 0.00151118 3.3 0.0015110999999999998 3.3 0.0015111999999999999 0 0.00151112 0 0.00151122 3.3 0.00151114 3.3 0.00151124 0 0.0015111599999999999 0 0.00151126 3.3 0.00151118 3.3 0.00151128 0 0.0015111999999999999 0 0.0015113 3.3 0.00151122 3.3 0.00151132 0 0.0015112399999999998 0 0.00151134 3.3 0.00151126 3.3 0.00151136 0 0.0015112799999999998 0 0.0015113799999999999 3.3 0.0015113 3.3 0.0015114 0 0.0015113199999999998 0 0.0015114199999999999 3.3 0.00151134 3.3 0.00151144 0 0.00151136 0 0.00151146 3.3 0.0015113799999999999 3.3 0.00151148 0 0.0015114 0 0.0015115 3.3 0.0015114199999999999 3.3 0.00151152 0 0.00151144 0 0.00151154 3.3 0.0015114599999999998 3.3 0.00151156 0 0.00151148 0 0.00151158 3.3 0.0015114999999999998 3.3 0.0015115999999999999 0 0.00151152 0 0.00151162 3.3 0.00151154 3.3 0.00151164 0 0.00151156 0 0.00151166 3.3 0.00151158 3.3 0.00151168 0 0.0015115999999999999 0 0.0015117 3.3 0.00151162 3.3 0.00151172 0 0.0015116399999999999 0 0.00151174 3.3 0.00151166 3.3 0.00151176 0 0.0015116799999999998 0 0.00151178 3.3 0.0015117 3.3 0.0015118 0 0.0015117199999999998 0 0.0015118199999999999 3.3 0.00151174 3.3 0.00151184 0 0.00151176 0 0.00151186 3.3 0.00151178 3.3 0.00151188 0 0.0015118 0 0.0015119 3.3 0.0015118199999999999 3.3 0.00151192 0 0.00151184 0 0.00151194 3.3 0.0015118599999999999 3.3 0.00151196 0 0.00151188 0 0.00151198 3.3 0.0015118999999999998 3.3 0.0015119999999999999 0 0.00151192 0 0.00151202 3.3 0.0015119399999999998 3.3 0.0015120399999999999 0 0.00151196 0 0.00151206 3.3 0.00151198 3.3 0.00151208 0 0.0015119999999999999 0 0.0015121 3.3 0.00151202 3.3 0.00151212 0 0.0015120399999999999 0 0.00151214 3.3 0.00151206 3.3 0.00151216 0 0.0015120799999999998 0 0.00151218 3.3 0.0015121 3.3 0.0015122 0 0.0015121199999999998 0 0.0015122199999999999 3.3 0.00151214 3.3 0.00151224 0 0.0015121599999999998 0 0.0015122599999999999 3.3 0.00151218 3.3 0.00151228 0 0.0015122 0 0.0015123 3.3 0.0015122199999999999 3.3 0.00151232 0 0.00151224 0 0.00151234 3.3 0.0015122599999999999 3.3 0.00151236 0 0.00151228 0 0.00151238 3.3 0.0015122999999999998 3.3 0.0015124 0 0.00151232 0 0.00151242 3.3 0.0015123399999999998 3.3 0.0015124399999999999 0 0.00151236 0 0.00151246 3.3 0.00151238 3.3 0.00151248 0 0.0015124 0 0.0015125 3.3 0.00151242 3.3 0.00151252 0 0.0015124399999999999 0 0.00151254 3.3 0.00151246 3.3 0.00151256 0 0.0015124799999999999 0 0.00151258 3.3 0.0015125 3.3 0.0015126 0 0.0015125199999999998 0 0.00151262 3.3 0.00151254 3.3 0.00151264 0 0.0015125599999999998 0 0.0015126599999999999 3.3 0.00151258 3.3 0.00151268 0 0.0015126 0 0.0015127 3.3 0.00151262 3.3 0.00151272 0 0.00151264 0 0.00151274 3.3 0.0015126599999999999 3.3 0.00151276 0 0.00151268 0 0.00151278 3.3 0.0015126999999999999 3.3 0.0015128 0 0.00151272 0 0.00151282 3.3 0.0015127399999999998 3.3 0.0015128399999999999 0 0.00151276 0 0.00151286 3.3 0.0015127799999999998 3.3 0.0015128799999999999 0 0.0015128 0 0.0015129 3.3 0.00151282 3.3 0.00151292 0 0.0015128399999999999 0 0.00151294 3.3 0.00151286 3.3 0.00151296 0 0.0015128799999999999 0 0.00151298 3.3 0.0015129 3.3 0.001513 0 0.0015129199999999998 0 0.00151302 3.3 0.00151294 3.3 0.00151304 0 0.0015129599999999998 0 0.0015130599999999999 3.3 0.00151298 3.3 0.00151308 0 0.0015129999999999998 0 0.0015130999999999999 3.3 0.00151302 3.3 0.00151312 0 0.00151304 0 0.00151314 3.3 0.0015130599999999999 3.3 0.00151316 0 0.00151308 0 0.00151318 3.3 0.0015130999999999999 3.3 0.0015132 0 0.00151312 0 0.00151322 3.3 0.0015131399999999998 3.3 0.00151324 0 0.00151316 0 0.00151326 3.3 0.0015131799999999998 3.3 0.0015132799999999999 0 0.0015132 0 0.0015133 3.3 0.00151322 3.3 0.00151332 0 0.00151324 0 0.00151334 3.3 0.00151326 3.3 0.00151336 0 0.0015132799999999999 0 0.00151338 3.3 0.0015133 3.3 0.0015134 0 0.0015133199999999999 0 0.00151342 3.3 0.00151334 3.3 0.00151344 0 0.0015133599999999998 0 0.00151346 3.3 0.00151338 3.3 0.00151348 0 0.0015133999999999998 0 0.0015134999999999999 3.3 0.00151342 3.3 0.00151352 0 0.00151344 0 0.00151354 3.3 0.00151346 3.3 0.00151356 0 0.00151348 0 0.00151358 3.3 0.0015134999999999999 3.3 0.0015136 0 0.00151352 0 0.00151362 3.3 0.0015135399999999999 3.3 0.00151364 0 0.00151356 0 0.00151366 3.3 0.0015135799999999998 3.3 0.0015136799999999999 0 0.0015136 0 0.0015137 3.3 0.0015136199999999998 3.3 0.0015137199999999999 0 0.00151364 0 0.00151374 3.3 0.00151366 3.3 0.00151376 0 0.0015136799999999999 0 0.00151378 3.3 0.0015137 3.3 0.0015138 0 0.0015137199999999999 0 0.00151382 3.3 0.00151374 3.3 0.00151384 0 0.0015137599999999998 0 0.00151386 3.3 0.00151378 3.3 0.00151388 0 0.0015137999999999998 0 0.0015138999999999999 3.3 0.00151382 3.3 0.00151392 0 0.00151384 0 0.00151394 3.3 0.00151386 3.3 0.00151396 0 0.00151388 0 0.00151398 3.3 0.0015138999999999999 3.3 0.001514 0 0.00151392 0 0.00151402 3.3 0.0015139399999999999 3.3 0.00151404 0 0.00151396 0 0.00151406 3.3 0.0015139799999999998 3.3 0.00151408 0 0.001514 0 0.0015141 3.3 0.0015140199999999998 3.3 0.0015141199999999999 0 0.00151404 0 0.00151414 3.3 0.00151406 3.3 0.00151416 0 0.00151408 0 0.00151418 3.3 0.0015141 3.3 0.0015142 0 0.0015141199999999999 0 0.00151422 3.3 0.00151414 3.3 0.00151424 0 0.0015141599999999999 0 0.00151426 3.3 0.00151418 3.3 0.00151428 0 0.0015141999999999998 0 0.0015142999999999999 3.3 0.00151422 3.3 0.00151432 0 0.0015142399999999998 0 0.0015143399999999999 3.3 0.00151426 3.3 0.00151436 0 0.00151428 0 0.00151438 3.3 0.0015142999999999999 3.3 0.0015144 0 0.00151432 0 0.00151442 3.3 0.0015143399999999999 3.3 0.00151444 0 0.00151436 0 0.00151446 3.3 0.0015143799999999998 3.3 0.00151448 0 0.0015144 0 0.0015145 3.3 0.0015144199999999998 3.3 0.0015145199999999999 0 0.00151444 0 0.00151454 3.3 0.0015144599999999998 3.3 0.0015145599999999999 0 0.00151448 0 0.00151458 3.3 0.0015145 3.3 0.0015146 0 0.0015145199999999999 0 0.00151462 3.3 0.00151454 3.3 0.00151464 0 0.0015145599999999999 0 0.00151466 3.3 0.00151458 3.3 0.00151468 0 0.0015145999999999998 0 0.0015147 3.3 0.00151462 3.3 0.00151472 0 0.0015146399999999998 0 0.0015147399999999999 3.3 0.00151466 3.3 0.00151476 0 0.00151468 0 0.00151478 3.3 0.0015147 3.3 0.0015148 0 0.00151472 0 0.00151482 3.3 0.0015147399999999999 3.3 0.00151484 0 0.00151476 0 0.00151486 3.3 0.0015147799999999999 3.3 0.00151488 0 0.0015148 0 0.0015149 3.3 0.0015148199999999998 3.3 0.00151492 0 0.00151484 0 0.00151494 3.3 0.0015148599999999998 3.3 0.0015149599999999999 0 0.00151488 0 0.00151498 3.3 0.0015149 3.3 0.001515 0 0.00151492 0 0.00151502 3.3 0.00151494 3.3 0.00151504 0 0.0015149599999999999 0 0.00151506 3.3 0.00151498 3.3 0.00151508 0 0.0015149999999999999 0 0.0015151 3.3 0.00151502 3.3 0.00151512 0 0.0015150399999999998 0 0.0015151399999999999 3.3 0.00151506 3.3 0.00151516 0 0.0015150799999999998 0 0.0015151799999999999 3.3 0.0015151 3.3 0.0015152 0 0.00151512 0 0.00151522 3.3 0.0015151399999999999 3.3 0.00151524 0 0.00151516 0 0.00151526 3.3 0.0015151799999999999 3.3 0.00151528 0 0.0015152 0 0.0015153 3.3 0.0015152199999999998 3.3 0.00151532 0 0.00151524 0 0.00151534 3.3 0.0015152599999999998 3.3 0.0015153599999999999 0 0.00151528 0 0.00151538 3.3 0.0015152999999999998 3.3 0.0015153999999999999 0 0.00151532 0 0.00151542 3.3 0.00151534 3.3 0.00151544 0 0.0015153599999999999 0 0.00151546 3.3 0.00151538 3.3 0.00151548 0 0.0015153999999999999 0 0.0015155 3.3 0.00151542 3.3 0.00151552 0 0.0015154399999999998 0 0.00151554 3.3 0.00151546 3.3 0.00151556 0 0.0015154799999999998 0 0.0015155799999999999 3.3 0.0015155 3.3 0.0015156 0 0.00151552 0 0.00151562 3.3 0.00151554 3.3 0.00151564 0 0.00151556 0 0.00151566 3.3 0.0015155799999999999 3.3 0.00151568 0 0.0015156 0 0.0015157 3.3 0.0015156199999999999 3.3 0.00151572 0 0.00151564 0 0.00151574 3.3 0.0015156599999999998 3.3 0.00151576 0 0.00151568 0 0.00151578 3.3 0.0015156999999999998 3.3 0.0015157999999999999 0 0.00151572 0 0.00151582 3.3 0.00151574 3.3 0.00151584 0 0.00151576 0 0.00151586 3.3 0.00151578 3.3 0.00151588 0 0.0015157999999999999 0 0.0015159 3.3 0.00151582 3.3 0.00151592 0 0.0015158399999999999 0 0.00151594 3.3 0.00151586 3.3 0.00151596 0 0.0015158799999999998 0 0.0015159799999999999 3.3 0.0015159 3.3 0.001516 0 0.0015159199999999998 0 0.0015160199999999999 3.3 0.00151594 3.3 0.00151604 0 0.00151596 0 0.00151606 3.3 0.0015159799999999999 3.3 0.00151608 0 0.001516 0 0.0015161 3.3 0.0015160199999999999 3.3 0.00151612 0 0.00151604 0 0.00151614 3.3 0.0015160599999999998 3.3 0.00151616 0 0.00151608 0 0.00151618 3.3 0.0015160999999999998 3.3 0.0015161999999999999 0 0.00151612 0 0.00151622 3.3 0.0015161399999999998 3.3 0.0015162399999999999 0 0.00151616 0 0.00151626 3.3 0.00151618 3.3 0.00151628 0 0.0015161999999999999 0 0.0015163 3.3 0.00151622 3.3 0.00151632 0 0.0015162399999999999 0 0.00151634 3.3 0.00151626 3.3 0.00151636 0 0.0015162799999999998 0 0.00151638 3.3 0.0015163 3.3 0.0015164 0 0.0015163199999999998 0 0.0015164199999999999 3.3 0.00151634 3.3 0.00151644 0 0.00151636 0 0.00151646 3.3 0.00151638 3.3 0.00151648 0 0.0015164 0 0.0015165 3.3 0.0015164199999999999 3.3 0.00151652 0 0.00151644 0 0.00151654 3.3 0.0015164599999999999 3.3 0.00151656 0 0.00151648 0 0.00151658 3.3 0.0015164999999999998 3.3 0.0015166 0 0.00151652 0 0.00151662 3.3 0.0015165399999999998 3.3 0.0015166399999999999 0 0.00151656 0 0.00151666 3.3 0.00151658 3.3 0.00151668 0 0.0015166 0 0.0015167 3.3 0.00151662 3.3 0.00151672 0 0.0015166399999999999 0 0.00151674 3.3 0.00151666 3.3 0.00151676 0 0.0015166799999999999 0 0.00151678 3.3 0.0015167 3.3 0.0015168 0 0.0015167199999999998 0 0.0015168199999999999 3.3 0.00151674 3.3 0.00151684 0 0.0015167599999999998 0 0.0015168599999999999 3.3 0.00151678 3.3 0.00151688 0 0.0015168 0 0.0015169 3.3 0.0015168199999999999 3.3 0.00151692 0 0.00151684 0 0.00151694 3.3 0.0015168599999999999 3.3 0.00151696 0 0.00151688 0 0.00151698 3.3 0.0015168999999999998 3.3 0.001517 0 0.00151692 0 0.00151702 3.3 0.0015169399999999998 3.3 0.0015170399999999999 0 0.00151696 0 0.00151706 3.3 0.00151698 3.3 0.00151708 0 0.001517 0 0.0015171 3.3 0.00151702 3.3 0.00151712 0 0.0015170399999999999 0 0.00151714 3.3 0.00151706 3.3 0.00151716 0 0.0015170799999999999 0 0.00151718 3.3 0.0015171 3.3 0.0015172 0 0.0015171199999999998 0 0.00151722 3.3 0.00151714 3.3 0.00151724 0 0.0015171599999999998 0 0.0015172599999999999 3.3 0.00151718 3.3 0.00151728 0 0.0015172 0 0.0015173 3.3 0.00151722 3.3 0.00151732 0 0.00151724 0 0.00151734 3.3 0.0015172599999999999 3.3 0.00151736 0 0.00151728 0 0.00151738 3.3 0.0015172999999999999 3.3 0.0015174 0 0.00151732 0 0.00151742 3.3 0.0015173399999999998 3.3 0.0015174399999999999 0 0.00151736 0 0.00151746 3.3 0.0015173799999999998 3.3 0.0015174799999999999 0 0.0015174 0 0.0015175 3.3 0.00151742 3.3 0.00151752 0 0.0015174399999999999 0 0.00151754 3.3 0.00151746 3.3 0.00151756 0 0.0015174799999999999 0 0.00151758 3.3 0.0015175 3.3 0.0015176 0 0.0015175199999999998 0 0.00151762 3.3 0.00151754 3.3 0.00151764 0 0.0015175599999999998 0 0.0015176599999999999 3.3 0.00151758 3.3 0.00151768 0 0.0015175999999999998 0 0.0015176999999999999 3.3 0.00151762 3.3 0.00151772 0 0.00151764 0 0.00151774 3.3 0.0015176599999999999 3.3 0.00151776 0 0.00151768 0 0.00151778 3.3 0.0015176999999999999 3.3 0.0015178 0 0.00151772 0 0.00151782 3.3 0.0015177399999999998 3.3 0.00151784 0 0.00151776 0 0.00151786 3.3 0.0015177799999999998 3.3 0.0015178799999999999 0 0.0015178 0 0.0015179 3.3 0.00151782 3.3 0.00151792 0 0.00151784 0 0.00151794 3.3 0.00151786 3.3 0.00151796 0 0.0015178799999999999 0 0.00151798 3.3 0.0015179 3.3 0.001518 0 0.0015179199999999999 0 0.00151802 3.3 0.00151794 3.3 0.00151804 0 0.0015179599999999998 0 0.00151806 3.3 0.00151798 3.3 0.00151808 0 0.0015179999999999998 0 0.0015180999999999999 3.3 0.00151802 3.3 0.00151812 0 0.00151804 0 0.00151814 3.3 0.00151806 3.3 0.00151816 0 0.00151808 0 0.00151818 3.3 0.0015180999999999999 3.3 0.0015182 0 0.00151812 0 0.00151822 3.3 0.0015181399999999999 3.3 0.00151824 0 0.00151816 0 0.00151826 3.3 0.0015181799999999998 3.3 0.0015182799999999999 0 0.0015182 0 0.0015183 3.3 0.0015182199999999998 3.3 0.0015183199999999999 0 0.00151824 0 0.00151834 3.3 0.00151826 3.3 0.00151836 0 0.0015182799999999999 0 0.00151838 3.3 0.0015183 3.3 0.0015184 0 0.0015183199999999999 0 0.00151842 3.3 0.00151834 3.3 0.00151844 0 0.0015183599999999998 0 0.00151846 3.3 0.00151838 3.3 0.00151848 0 0.0015183999999999998 0 0.0015184999999999999 3.3 0.00151842 3.3 0.00151852 0 0.0015184399999999998 0 0.0015185399999999999 3.3 0.00151846 3.3 0.00151856 0 0.00151848 0 0.00151858 3.3 0.0015184999999999999 3.3 0.0015186 0 0.00151852 0 0.00151862 3.3 0.0015185399999999999 3.3 0.00151864 0 0.00151856 0 0.00151866 3.3 0.0015185799999999998 3.3 0.00151868 0 0.0015186 0 0.0015187 3.3 0.0015186199999999998 3.3 0.0015187199999999999 0 0.00151864 0 0.00151874 3.3 0.00151866 3.3 0.00151876 0 0.00151868 0 0.00151878 3.3 0.0015187 3.3 0.0015188 0 0.0015187199999999999 0 0.00151882 3.3 0.00151874 3.3 0.00151884 0 0.0015187599999999999 0 0.00151886 3.3 0.00151878 3.3 0.00151888 0 0.0015187999999999998 0 0.0015189 3.3 0.00151882 3.3 0.00151892 0 0.0015188399999999998 0 0.0015189399999999999 3.3 0.00151886 3.3 0.00151896 0 0.00151888 0 0.00151898 3.3 0.0015189 3.3 0.001519 0 0.00151892 0 0.00151902 3.3 0.0015189399999999999 3.3 0.00151904 0 0.00151896 0 0.00151906 3.3 0.0015189799999999999 3.3 0.00151908 0 0.001519 0 0.0015191 3.3 0.0015190199999999998 3.3 0.0015191199999999999 0 0.00151904 0 0.00151914 3.3 0.0015190599999999998 3.3 0.0015191599999999999 0 0.00151908 0 0.00151918 3.3 0.0015191 3.3 0.0015192 0 0.0015191199999999999 0 0.00151922 3.3 0.00151914 3.3 0.00151924 0 0.0015191599999999999 0 0.00151926 3.3 0.00151918 3.3 0.00151928 0 0.0015191999999999998 0 0.0015193 3.3 0.00151922 3.3 0.00151932 0 0.0015192399999999998 0 0.0015193399999999999 3.3 0.00151926 3.3 0.00151936 0 0.0015192799999999998 0 0.0015193799999999999 3.3 0.0015193 3.3 0.0015194 0 0.00151932 0 0.00151942 3.3 0.0015193399999999999 3.3 0.00151944 0 0.00151936 0 0.00151946 3.3 0.0015193799999999999 3.3 0.00151948 0 0.0015194 0 0.0015195 3.3 0.0015194199999999998 3.3 0.00151952 0 0.00151944 0 0.00151954 3.3 0.0015194599999999998 3.3 0.0015195599999999999 0 0.00151948 0 0.00151958 3.3 0.0015195 3.3 0.0015196 0 0.00151952 0 0.00151962 3.3 0.00151954 3.3 0.00151964 0 0.0015195599999999999 0 0.00151966 3.3 0.00151958 3.3 0.00151968 0 0.0015195999999999999 0 0.0015197 3.3 0.00151962 3.3 0.00151972 0 0.0015196399999999998 0 0.00151974 3.3 0.00151966 3.3 0.00151976 0 0.0015196799999999998 0 0.0015197799999999999 3.3 0.0015197 3.3 0.0015198 0 0.00151972 0 0.00151982 3.3 0.00151974 3.3 0.00151984 0 0.00151976 0 0.00151986 3.3 0.0015197799999999999 3.3 0.00151988 0 0.0015198 0 0.0015199 3.3 0.0015198199999999999 3.3 0.00151992 0 0.00151984 0 0.00151994 3.3 0.0015198599999999998 3.3 0.0015199599999999999 0 0.00151988 0 0.00151998 3.3 0.0015198999999999998 3.3 0.0015199999999999999 0 0.00151992 0 0.00152002 3.3 0.00151994 3.3 0.00152004 0 0.0015199599999999999 0 0.00152006 3.3 0.00151998 3.3 0.00152008 0 0.0015199999999999999 0 0.0015201 3.3 0.00152002 3.3 0.00152012 0 0.0015200399999999998 0 0.00152014 3.3 0.00152006 3.3 0.00152016 0 0.0015200799999999998 0 0.0015201799999999999 3.3 0.0015201 3.3 0.0015202 0 0.0015201199999999998 0 0.0015202199999999999 3.3 0.00152014 3.3 0.00152024 0 0.00152016 0 0.00152026 3.3 0.0015201799999999999 3.3 0.00152028 0 0.0015202 0 0.0015203 3.3 0.0015202199999999999 3.3 0.00152032 0 0.00152024 0 0.00152034 3.3 0.0015202599999999998 3.3 0.00152036 0 0.00152028 0 0.00152038 3.3 0.0015202999999999998 3.3 0.0015203999999999999 0 0.00152032 0 0.00152042 3.3 0.00152034 3.3 0.00152044 0 0.00152036 0 0.00152046 3.3 0.00152038 3.3 0.00152048 0 0.0015203999999999999 0 0.0015205 3.3 0.00152042 3.3 0.00152052 0 0.0015204399999999999 0 0.00152054 3.3 0.00152046 3.3 0.00152056 0 0.0015204799999999998 0 0.00152058 3.3 0.0015205 3.3 0.0015206 0 0.0015205199999999998 0 0.0015206199999999999 3.3 0.00152054 3.3 0.00152064 0 0.00152056 0 0.00152066 3.3 0.00152058 3.3 0.00152068 0 0.0015206 0 0.0015207 3.3 0.0015206199999999999 3.3 0.00152072 0 0.00152064 0 0.00152074 3.3 0.0015206599999999999 3.3 0.00152076 0 0.00152068 0 0.00152078 3.3 0.0015206999999999998 3.3 0.0015207999999999999 0 0.00152072 0 0.00152082 3.3 0.0015207399999999998 3.3 0.0015208399999999999 0 0.00152076 0 0.00152086 3.3 0.00152078 3.3 0.00152088 0 0.0015207999999999999 0 0.0015209 3.3 0.00152082 3.3 0.00152092 0 0.0015208399999999999 0 0.00152094 3.3 0.00152086 3.3 0.00152096 0 0.0015208799999999998 0 0.00152098 3.3 0.0015209 3.3 0.001521 0 0.0015209199999999998 0 0.0015210199999999999 3.3 0.00152094 3.3 0.00152104 0 0.00152096 0 0.00152106 3.3 0.00152098 3.3 0.00152108 0 0.001521 0 0.0015211 3.3 0.0015210199999999999 3.3 0.00152112 0 0.00152104 0 0.00152114 3.3 0.0015210599999999999 3.3 0.00152116 0 0.00152108 0 0.00152118 3.3 0.0015210999999999998 3.3 0.0015212 0 0.00152112 0 0.00152122 3.3 0.0015211399999999998 3.3 0.0015212399999999999 0 0.00152116 0 0.00152126 3.3 0.00152118 3.3 0.00152128 0 0.0015212 0 0.0015213 3.3 0.00152122 3.3 0.00152132 0 0.0015212399999999999 0 0.00152134 3.3 0.00152126 3.3 0.00152136 0 0.0015212799999999999 0 0.00152138 3.3 0.0015213 3.3 0.0015214 0 0.0015213199999999998 0 0.0015214199999999999 3.3 0.00152134 3.3 0.00152144 0 0.0015213599999999998 0 0.0015214599999999999 3.3 0.00152138 3.3 0.00152148 0 0.0015214 0 0.0015215 3.3 0.0015214199999999999 3.3 0.00152152 0 0.00152144 0 0.00152154 3.3 0.0015214599999999999 3.3 0.00152156 0 0.00152148 0 0.00152158 3.3 0.0015214999999999998 3.3 0.0015216 0 0.00152152 0 0.00152162 3.3 0.0015215399999999998 3.3 0.0015216399999999999 0 0.00152156 0 0.00152166 3.3 0.0015215799999999998 3.3 0.0015216799999999999 0 0.0015216 0 0.0015217 3.3 0.00152162 3.3 0.00152172 0 0.0015216399999999999 0 0.00152174 3.3 0.00152166 3.3 0.00152176 0 0.0015216799999999999 0 0.00152178 3.3 0.0015217 3.3 0.0015218 0 0.0015217199999999998 0 0.00152182 3.3 0.00152174 3.3 0.00152184 0 0.0015217599999999998 0 0.0015218599999999999 3.3 0.00152178 3.3 0.00152188 0 0.0015218 0 0.0015219 3.3 0.00152182 3.3 0.00152192 0 0.00152184 0 0.00152194 3.3 0.0015218599999999999 3.3 0.00152196 0 0.00152188 0 0.00152198 3.3 0.0015218999999999999 3.3 0.001522 0 0.00152192 0 0.00152202 3.3 0.0015219399999999998 3.3 0.00152204 0 0.00152196 0 0.00152206 3.3 0.0015219799999999998 3.3 0.0015220799999999999 0 0.001522 0 0.0015221 3.3 0.00152202 3.3 0.00152212 0 0.00152204 0 0.00152214 3.3 0.00152206 3.3 0.00152216 0 0.0015220799999999999 0 0.00152218 3.3 0.0015221 3.3 0.0015222 0 0.0015221199999999999 0 0.00152222 3.3 0.00152214 3.3 0.00152224 0 0.0015221599999999998 0 0.0015222599999999999 3.3 0.00152218 3.3 0.00152228 0 0.0015221999999999998 0 0.0015222999999999999 3.3 0.00152222 3.3 0.00152232 0 0.00152224 0 0.00152234 3.3 0.0015222599999999999 3.3 0.00152236 0 0.00152228 0 0.00152238 3.3 0.0015222999999999999 3.3 0.0015224 0 0.00152232 0 0.00152242 3.3 0.0015223399999999998 3.3 0.00152244 0 0.00152236 0 0.00152246 3.3 0.0015223799999999998 3.3 0.0015224799999999999 0 0.0015224 0 0.0015225 3.3 0.0015224199999999998 3.3 0.0015225199999999999 0 0.00152244 0 0.00152254 3.3 0.00152246 3.3 0.00152256 0 0.0015224799999999999 0 0.00152258 3.3 0.0015225 3.3 0.0015226 0 0.0015225199999999999 0 0.00152262 3.3 0.00152254 3.3 0.00152264 0 0.0015225599999999998 0 0.00152266 3.3 0.00152258 3.3 0.00152268 0 0.0015225999999999998 0 0.0015226999999999999 3.3 0.00152262 3.3 0.00152272 0 0.00152264 0 0.00152274 3.3 0.00152266 3.3 0.00152276 0 0.00152268 0 0.00152278 3.3 0.0015226999999999999 3.3 0.0015228 0 0.00152272 0 0.00152282 3.3 0.0015227399999999999 3.3 0.00152284 0 0.00152276 0 0.00152286 3.3 0.0015227799999999998 3.3 0.00152288 0 0.0015228 0 0.0015229 3.3 0.0015228199999999998 3.3 0.0015229199999999999 0 0.00152284 0 0.00152294 3.3 0.00152286 3.3 0.00152296 0 0.00152288 0 0.00152298 3.3 0.0015229 3.3 0.001523 0 0.0015229199999999999 0 0.00152302 3.3 0.00152294 3.3 0.00152304 0 0.0015229599999999999 0 0.00152306 3.3 0.00152298 3.3 0.00152308 0 0.0015229999999999998 0 0.0015230999999999999 3.3 0.00152302 3.3 0.00152312 0 0.0015230399999999998 0 0.0015231399999999999 3.3 0.00152306 3.3 0.00152316 0 0.00152308 0 0.00152318 3.3 0.0015230999999999999 3.3 0.0015232 0 0.00152312 0 0.00152322 3.3 0.0015231399999999999 3.3 0.00152324 0 0.00152316 0 0.00152326 3.3 0.0015231799999999998 3.3 0.00152328 0 0.0015232 0 0.0015233 3.3 0.0015232199999999998 3.3 0.0015233199999999999 0 0.00152324 0 0.00152334 3.3 0.0015232599999999998 3.3 0.0015233599999999999 0 0.00152328 0 0.00152338 3.3 0.0015233 3.3 0.0015234 0 0.0015233199999999999 0 0.00152342 3.3 0.00152334 3.3 0.00152344 0 0.0015233599999999999 0 0.00152346 3.3 0.00152338 3.3 0.00152348 0 0.0015233999999999998 0 0.0015235 3.3 0.00152342 3.3 0.00152352 0 0.0015234399999999998 0 0.0015235399999999999 3.3 0.00152346 3.3 0.00152356 0 0.00152348 0 0.00152358 3.3 0.0015235 3.3 0.0015236 0 0.00152352 0 0.00152362 3.3 0.0015235399999999999 3.3 0.00152364 0 0.00152356 0 0.00152366 3.3 0.0015235799999999999 3.3 0.00152368 0 0.0015236 0 0.0015237 3.3 0.0015236199999999998 3.3 0.00152372 0 0.00152364 0 0.00152374 3.3 0.0015236599999999998 3.3 0.0015237599999999999 0 0.00152368 0 0.00152378 3.3 0.0015237 3.3 0.0015238 0 0.00152372 0 0.00152382 3.3 0.00152374 3.3 0.00152384 0 0.0015237599999999999 0 0.00152386 3.3 0.00152378 3.3 0.00152388 0 0.0015237999999999999 0 0.0015239 3.3 0.00152382 3.3 0.00152392 0 0.0015238399999999998 0 0.0015239399999999999 3.3 0.00152386 3.3 0.00152396 0 0.0015238799999999998 0 0.0015239799999999999 3.3 0.0015239 3.3 0.001524 0 0.00152392 0 0.00152402 3.3 0.0015239399999999999 3.3 0.00152404 0 0.00152396 0 0.00152406 3.3 0.0015239799999999999 3.3 0.00152408 0 0.001524 0 0.0015241 3.3 0.0015240199999999998 3.3 0.00152412 0 0.00152404 0 0.00152414 3.3 0.0015240599999999998 3.3 0.0015241599999999999 0 0.00152408 0 0.00152418 3.3 0.0015241 3.3 0.0015242 0 0.00152412 0 0.00152422 3.3 0.00152414 3.3 0.00152424 0 0.0015241599999999999 0 0.00152426 3.3 0.00152418 3.3 0.00152428 0 0.0015241999999999999 0 0.0015243 3.3 0.00152422 3.3 0.00152432 0 0.0015242399999999998 0 0.00152434 3.3 0.00152426 3.3 0.00152436 0 0.0015242799999999998 0 0.0015243799999999999 3.3 0.0015243 3.3 0.0015244 0 0.00152432 0 0.00152442 3.3 0.00152434 3.3 0.00152444 0 0.00152436 0 0.00152446 3.3 0.0015243799999999999 3.3 0.00152448 0 0.0015244 0 0.0015245 3.3 0.0015244199999999999 3.3 0.00152452 0 0.00152444 0 0.00152454 3.3 0.0015244599999999998 3.3 0.0015245599999999999 0 0.00152448 0 0.00152458 3.3 0.0015244999999999998 3.3 0.0015245999999999999 0 0.00152452 0 0.00152462 3.3 0.00152454 3.3 0.00152464 0 0.0015245599999999999 0 0.00152466 3.3 0.00152458 3.3 0.00152468 0 0.0015245999999999999 0 0.0015247 3.3 0.00152462 3.3 0.00152472 0 0.0015246399999999998 0 0.00152474 3.3 0.00152466 3.3 0.00152476 0 0.0015246799999999998 0 0.0015247799999999999 3.3 0.0015247 3.3 0.0015248 0 0.0015247199999999998 0 0.0015248199999999999 3.3 0.00152474 3.3 0.00152484 0 0.00152476 0 0.00152486 3.3 0.0015247799999999999 3.3 0.00152488 0 0.0015248 0 0.0015249 3.3 0.0015248199999999999 3.3 0.00152492 0 0.00152484 0 0.00152494 3.3 0.0015248599999999998 3.3 0.00152496 0 0.00152488 0 0.00152498 3.3 0.0015248999999999998 3.3 0.0015249999999999999 0 0.00152492 0 0.00152502 3.3 0.00152494 3.3 0.00152504 0 0.00152496 0 0.00152506 3.3 0.00152498 3.3 0.00152508 0 0.0015249999999999999 0 0.0015251 3.3 0.00152502 3.3 0.00152512 0 0.0015250399999999999 0 0.00152514 3.3 0.00152506 3.3 0.00152516 0 0.0015250799999999998 0 0.00152518 3.3 0.0015251 3.3 0.0015252 0 0.0015251199999999998 0 0.0015252199999999999 3.3 0.00152514 3.3 0.00152524 0 0.00152516 0 0.00152526 3.3 0.00152518 3.3 0.00152528 0 0.0015252 0 0.0015253 3.3 0.0015252199999999999 3.3 0.00152532 0 0.00152524 0 0.00152534 3.3 0.0015252599999999999 3.3 0.00152536 0 0.00152528 0 0.00152538 3.3 0.0015252999999999998 3.3 0.0015253999999999999 0 0.00152532 0 0.00152542 3.3 0.0015253399999999998 3.3 0.0015254399999999999 0 0.00152536 0 0.00152546 3.3 0.00152538 3.3 0.00152548 0 0.0015253999999999999 0 0.0015255 3.3 0.00152542 3.3 0.00152552 0 0.0015254399999999999 0 0.00152554 3.3 0.00152546 3.3 0.00152556 0 0.0015254799999999998 0 0.00152558 3.3 0.0015255 3.3 0.0015256 0 0.0015255199999999998 0 0.0015256199999999999 3.3 0.00152554 3.3 0.00152564 0 0.0015255599999999998 0 0.0015256599999999999 3.3 0.00152558 3.3 0.00152568 0 0.0015256 0 0.0015257 3.3 0.0015256199999999999 3.3 0.00152572 0 0.00152564 0 0.00152574 3.3 0.0015256599999999999 3.3 0.00152576 0 0.00152568 0 0.00152578 3.3 0.0015256999999999998 3.3 0.0015258 0 0.00152572 0 0.00152582 3.3 0.0015257399999999998 3.3 0.0015258399999999999 0 0.00152576 0 0.00152586 3.3 0.00152578 3.3 0.00152588 0 0.0015258 0 0.0015259 3.3 0.00152582 3.3 0.00152592 0 0.0015258399999999999 0 0.00152594 3.3 0.00152586 3.3 0.00152596 0 0.0015258799999999999 0 0.00152598 3.3 0.0015259 3.3 0.001526 0 0.0015259199999999998 0 0.00152602 3.3 0.00152594 3.3 0.00152604 0 0.0015259599999999998 0 0.0015260599999999999 3.3 0.00152598 3.3 0.00152608 0 0.001526 0 0.0015261 3.3 0.00152602 3.3 0.00152612 0 0.00152604 0 0.00152614 3.3 0.0015260599999999999 3.3 0.00152616 0 0.00152608 0 0.00152618 3.3 0.0015260999999999999 3.3 0.0015262 0 0.00152612 0 0.00152622 3.3 0.0015261399999999998 3.3 0.0015262399999999999 0 0.00152616 0 0.00152626 3.3 0.0015261799999999998 3.3 0.0015262799999999999 0 0.0015262 0 0.0015263 3.3 0.00152622 3.3 0.00152632 0 0.0015262399999999999 0 0.00152634 3.3 0.00152626 3.3 0.00152636 0 0.0015262799999999999 0 0.00152638 3.3 0.0015263 3.3 0.0015264 0 0.0015263199999999998 0 0.00152642 3.3 0.00152634 3.3 0.00152644 0 0.0015263599999999998 0 0.0015264599999999999 3.3 0.00152638 3.3 0.00152648 0 0.0015263999999999998 0 0.0015264999999999999 3.3 0.00152642 3.3 0.00152652 0 0.00152644 0 0.00152654 3.3 0.0015264599999999999 3.3 0.00152656 0 0.00152648 0 0.00152658 3.3 0.0015264999999999999 3.3 0.0015266 0 0.00152652 0 0.00152662 3.3 0.0015265399999999998 3.3 0.00152664 0 0.00152656 0 0.00152666 3.3 0.0015265799999999998 3.3 0.0015266799999999999 0 0.0015266 0 0.0015267 3.3 0.00152662 3.3 0.00152672 0 0.00152664 0 0.00152674 3.3 0.00152666 3.3 0.00152676 0 0.0015266799999999999 0 0.00152678 3.3 0.0015267 3.3 0.0015268 0 0.0015267199999999999 0 0.00152682 3.3 0.00152674 3.3 0.00152684 0 0.0015267599999999998 0 0.00152686 3.3 0.00152678 3.3 0.00152688 0 0.0015267999999999998 0 0.0015268999999999999 3.3 0.00152682 3.3 0.00152692 0 0.00152684 0 0.00152694 3.3 0.00152686 3.3 0.00152696 0 0.00152688 0 0.00152698 3.3 0.0015268999999999999 3.3 0.001527 0 0.00152692 0 0.00152702 3.3 0.0015269399999999999 3.3 0.00152704 0 0.00152696 0 0.00152706 3.3 0.0015269799999999998 3.3 0.0015270799999999999 0 0.001527 0 0.0015271 3.3 0.0015270199999999998 3.3 0.0015271199999999999 0 0.00152704 0 0.00152714 3.3 0.00152706 3.3 0.00152716 0 0.0015270799999999999 0 0.00152718 3.3 0.0015271 3.3 0.0015272 0 0.0015271199999999999 0 0.00152722 3.3 0.00152714 3.3 0.00152724 0 0.0015271599999999998 0 0.00152726 3.3 0.00152718 3.3 0.00152728 0 0.0015271999999999998 0 0.0015272999999999999 3.3 0.00152722 3.3 0.00152732 0 0.0015272399999999998 0 0.0015273399999999999 3.3 0.00152726 3.3 0.00152736 0 0.00152728 0 0.00152738 3.3 0.0015272999999999999 3.3 0.0015274 0 0.00152732 0 0.00152742 3.3 0.0015273399999999999 3.3 0.00152744 0 0.00152736 0 0.00152746 3.3 0.0015273799999999998 3.3 0.00152748 0 0.0015274 0 0.0015275 3.3 0.0015274199999999998 3.3 0.0015275199999999999 0 0.00152744 0 0.00152754 3.3 0.00152746 3.3 0.00152756 0 0.00152748 0 0.00152758 3.3 0.0015275 3.3 0.0015276 0 0.0015275199999999999 0 0.00152762 3.3 0.00152754 3.3 0.00152764 0 0.0015275599999999999 0 0.00152766 3.3 0.00152758 3.3 0.00152768 0 0.0015275999999999998 0 0.0015276999999999999 3.3 0.00152762 3.3 0.00152772 0 0.0015276399999999998 0 0.0015277399999999999 3.3 0.00152766 3.3 0.00152776 0 0.00152768 0 0.00152778 3.3 0.0015276999999999999 3.3 0.0015278 0 0.00152772 0 0.00152782 3.3 0.0015277399999999999 3.3 0.00152784 0 0.00152776 0 0.00152786 3.3 0.0015277799999999998 3.3 0.00152788 0 0.0015278 0 0.0015279 3.3 0.0015278199999999998 3.3 0.0015279199999999999 0 0.00152784 0 0.00152794 3.3 0.0015278599999999998 3.3 0.0015279599999999999 0 0.00152788 0 0.00152798 3.3 0.0015279 3.3 0.001528 0 0.0015279199999999999 0 0.00152802 3.3 0.00152794 3.3 0.00152804 0 0.0015279599999999999 0 0.00152806 3.3 0.00152798 3.3 0.00152808 0 0.0015279999999999998 0 0.0015281 3.3 0.00152802 3.3 0.00152812 0 0.0015280399999999998 0 0.0015281399999999999 3.3 0.00152806 3.3 0.00152816 0 0.00152808 0 0.00152818 3.3 0.0015281 3.3 0.0015282 0 0.00152812 0 0.00152822 3.3 0.0015281399999999999 3.3 0.00152824 0 0.00152816 0 0.00152826 3.3 0.0015281799999999999 3.3 0.00152828 0 0.0015282 0 0.0015283 3.3 0.0015282199999999998 3.3 0.00152832 0 0.00152824 0 0.00152834 3.3 0.0015282599999999998 3.3 0.0015283599999999999 0 0.00152828 0 0.00152838 3.3 0.0015283 3.3 0.0015284 0 0.00152832 0 0.00152842 3.3 0.00152834 3.3 0.00152844 0 0.0015283599999999999 0 0.00152846 3.3 0.00152838 3.3 0.00152848 0 0.0015283999999999999 0 0.0015285 3.3 0.00152842 3.3 0.00152852 0 0.0015284399999999998 0 0.0015285399999999999 3.3 0.00152846 3.3 0.00152856 0 0.0015284799999999998 0 0.0015285799999999999 3.3 0.0015285 3.3 0.0015286 0 0.00152852 0 0.00152862 3.3 0.0015285399999999999 3.3 0.00152864 0 0.00152856 0 0.00152866 3.3 0.0015285799999999999 3.3 0.00152868 0 0.0015286 0 0.0015287 3.3 0.0015286199999999998 3.3 0.00152872 0 0.00152864 0 0.00152874 3.3 0.0015286599999999998 3.3 0.0015287599999999999 0 0.00152868 0 0.00152878 3.3 0.0015286999999999998 3.3 0.0015287999999999999 0 0.00152872 0 0.00152882 3.3 0.00152874 3.3 0.00152884 0 0.0015287599999999999 0 0.00152886 3.3 0.00152878 3.3 0.00152888 0 0.0015287999999999999 0 0.0015289 3.3 0.00152882 3.3 0.00152892 0 0.0015288399999999998 0 0.00152894 3.3 0.00152886 3.3 0.00152896 0 0.0015288799999999998 0 0.0015289799999999999 3.3 0.0015289 3.3 0.001529 0 0.00152892 0 0.00152902 3.3 0.00152894 3.3 0.00152904 0 0.00152896 0 0.00152906 3.3 0.0015289799999999999 3.3 0.00152908 0 0.001529 0 0.0015291 3.3 0.0015290199999999999 3.3 0.00152912 0 0.00152904 0 0.00152914 3.3 0.0015290599999999998 3.3 0.00152916 0 0.00152908 0 0.00152918 3.3 0.0015290999999999998 3.3 0.0015291999999999999 0 0.00152912 0 0.00152922 3.3 0.00152914 3.3 0.00152924 0 0.00152916 0 0.00152926 3.3 0.00152918 3.3 0.00152928 0 0.0015291999999999999 0 0.0015293 3.3 0.00152922 3.3 0.00152932 0 0.0015292399999999999 0 0.00152934 3.3 0.00152926 3.3 0.00152936 0 0.0015292799999999998 0 0.0015293799999999999 3.3 0.0015293 3.3 0.0015294 0 0.0015293199999999998 0 0.0015294199999999999 3.3 0.00152934 3.3 0.00152944 0 0.00152936 0 0.00152946 3.3 0.0015293799999999999 3.3 0.00152948 0 0.0015294 0 0.0015295 3.3 0.0015294199999999999 3.3 0.00152952 0 0.00152944 0 0.00152954 3.3 0.0015294599999999998 3.3 0.00152956 0 0.00152948 0 0.00152958 3.3 0.0015294999999999998 3.3 0.0015295999999999999 0 0.00152952 0 0.00152962 3.3 0.0015295399999999998 3.3 0.0015296399999999999 0 0.00152956 0 0.00152966 3.3 0.00152958 3.3 0.00152968 0 0.0015295999999999999 0 0.0015297 3.3 0.00152962 3.3 0.00152972 0 0.0015296399999999999 0 0.00152974 3.3 0.00152966 3.3 0.00152976 0 0.0015296799999999998 0 0.00152978 3.3 0.0015297 3.3 0.0015298 0 0.0015297199999999998 0 0.0015298199999999999 3.3 0.00152974 3.3 0.00152984 0 0.00152976 0 0.00152986 3.3 0.00152978 3.3 0.00152988 0 0.0015298 0 0.0015299 3.3 0.0015298199999999999 3.3 0.00152992 0 0.00152984 0 0.00152994 3.3 0.0015298599999999999 3.3 0.00152996 0 0.00152988 0 0.00152998 3.3 0.0015298999999999998 3.3 0.00153 0 0.00152992 0 0.00153002 3.3 0.0015299399999999998 3.3 0.0015300399999999999 0 0.00152996 0 0.00153006 3.3 0.00152998 3.3 0.00153008 0 0.00153 0 0.0015301 3.3 0.00153002 3.3 0.00153012 0 0.0015300399999999999 0 0.00153014 3.3 0.00153006 3.3 0.00153016 0 0.0015300799999999999 0 0.00153018 3.3 0.0015301 3.3 0.0015302 0 0.0015301199999999998 0 0.0015302199999999999 3.3 0.00153014 3.3 0.00153024 0 0.0015301599999999998 0 0.0015302599999999999 3.3 0.00153018 3.3 0.00153028 0 0.0015302 0 0.0015303 3.3 0.0015302199999999999 3.3 0.00153032 0 0.00153024 0 0.00153034 3.3 0.0015302599999999999 3.3 0.00153036 0 0.00153028 0 0.00153038 3.3 0.0015302999999999998 3.3 0.0015304 0 0.00153032 0 0.00153042 3.3 0.0015303399999999998 3.3 0.0015304399999999999 0 0.00153036 0 0.00153046 3.3 0.0015303799999999998 3.3 0.0015304799999999999 0 0.0015304 0 0.0015305 3.3 0.00153042 3.3 0.00153052 0 0.0015304399999999999 0 0.00153054 3.3 0.00153046 3.3 0.00153056 0 0.0015304799999999999 0 0.00153058 3.3 0.0015305 3.3 0.0015306 0 0.0015305199999999998 0 0.00153062 3.3 0.00153054 3.3 0.00153064 0 0.0015305599999999998 0 0.0015306599999999999 3.3 0.00153058 3.3 0.00153068 0 0.0015306 0 0.0015307 3.3 0.00153062 3.3 0.00153072 0 0.00153064 0 0.00153074 3.3 0.0015306599999999999 3.3 0.00153076 0 0.00153068 0 0.00153078 3.3 0.0015306999999999999 3.3 0.0015308 0 0.00153072 0 0.00153082 3.3 0.0015307399999999998 3.3 0.00153084 0 0.00153076 0 0.00153086 3.3 0.0015307799999999998 3.3 0.0015308799999999999 0 0.0015308 0 0.0015309 3.3 0.00153082 3.3 0.00153092 0 0.00153084 0 0.00153094 3.3 0.00153086 3.3 0.00153096 0 0.0015308799999999999 0 0.00153098 3.3 0.0015309 3.3 0.001531 0 0.0015309199999999999 0 0.00153102 3.3 0.00153094 3.3 0.00153104 0 0.0015309599999999998 0 0.0015310599999999999 3.3 0.00153098 3.3 0.00153108 0 0.0015309999999999998 0 0.0015310999999999999 3.3 0.00153102 3.3 0.00153112 0 0.00153104 0 0.00153114 3.3 0.0015310599999999999 3.3 0.00153116 0 0.00153108 0 0.00153118 3.3 0.0015310999999999999 3.3 0.0015312 0 0.00153112 0 0.00153122 3.3 0.0015311399999999998 3.3 0.00153124 0 0.00153116 0 0.00153126 3.3 0.0015311799999999998 3.3 0.0015312799999999999 0 0.0015312 0 0.0015313 3.3 0.00153122 3.3 0.00153132 0 0.00153124 0 0.00153134 3.3 0.00153126 3.3 0.00153136 0 0.0015312799999999999 0 0.00153138 3.3 0.0015313 3.3 0.0015314 0 0.0015313199999999999 0 0.00153142 3.3 0.00153134 3.3 0.00153144 0 0.0015313599999999998 0 0.00153146 3.3 0.00153138 3.3 0.00153148 0 0.0015313999999999998 0 0.0015314999999999999 3.3 0.00153142 3.3 0.00153152 0 0.00153144 0 0.00153154 3.3 0.00153146 3.3 0.00153156 0 0.00153148 0 0.00153158 3.3 0.0015314999999999999 3.3 0.0015316 0 0.00153152 0 0.00153162 3.3 0.0015315399999999999 3.3 0.00153164 0 0.00153156 0 0.00153166 3.3 0.0015315799999999998 3.3 0.0015316799999999999 0 0.0015316 0 0.0015317 3.3 0.0015316199999999998 3.3 0.0015317199999999999 0 0.00153164 0 0.00153174 3.3 0.00153166 3.3 0.00153176 0 0.0015316799999999999 0 0.00153178 3.3 0.0015317 3.3 0.0015318 0 0.0015317199999999999 0 0.00153182 3.3 0.00153174 3.3 0.00153184 0 0.0015317599999999998 0 0.00153186 3.3 0.00153178 3.3 0.00153188 0 0.0015317999999999998 0 0.0015318999999999999 3.3 0.00153182 3.3 0.00153192 0 0.0015318399999999998 0 0.0015319399999999999 3.3 0.00153186 3.3 0.00153196 0 0.00153188 0 0.00153198 3.3 0.0015318999999999999 3.3 0.001532 0 0.00153192 0 0.00153202 3.3 0.0015319399999999999 3.3 0.00153204 0 0.00153196 0 0.00153206 3.3 0.0015319799999999998 3.3 0.00153208 0 0.001532 0 0.0015321 3.3 0.0015320199999999998 3.3 0.0015321199999999999 0 0.00153204 0 0.00153214 3.3 0.00153206 3.3 0.00153216 0 0.00153208 0 0.00153218 3.3 0.0015321 3.3 0.0015322 0 0.0015321199999999999 0 0.00153222 3.3 0.00153214 3.3 0.00153224 0 0.0015321599999999999 0 0.00153226 3.3 0.00153218 3.3 0.00153228 0 0.0015321999999999998 0 0.0015323 3.3 0.00153222 3.3 0.00153232 0 0.0015322399999999998 0 0.0015323399999999999 3.3 0.00153226 3.3 0.00153236 0 0.00153228 0 0.00153238 3.3 0.0015323 3.3 0.0015324 0 0.00153232 0 0.00153242 3.3 0.0015323399999999999 3.3 0.00153244 0 0.00153236 0 0.00153246 3.3 0.0015323799999999999 3.3 0.00153248 0 0.0015324 0 0.0015325 3.3 0.0015324199999999998 3.3 0.0015325199999999999 0 0.00153244 0 0.00153254 3.3 0.0015324599999999998 3.3 0.0015325599999999999 0 0.00153248 0 0.00153258 3.3 0.0015325 3.3 0.0015326 0 0.0015325199999999999 0 0.00153262 3.3 0.00153254 3.3 0.00153264 0 0.0015325599999999999 0 0.00153266 3.3 0.00153258 3.3 0.00153268 0 0.0015325999999999998 0 0.0015327 3.3 0.00153262 3.3 0.00153272 0 0.0015326399999999998 0 0.0015327399999999999 3.3 0.00153266 3.3 0.00153276 0 0.0015326799999999998 0 0.0015327799999999999 3.3 0.0015327 3.3 0.0015328 0 0.00153272 0 0.00153282 3.3 0.0015327399999999999 3.3 0.00153284 0 0.00153276 0 0.00153286 3.3 0.0015327799999999999 3.3 0.00153288 0 0.0015328 0 0.0015329 3.3 0.0015328199999999998 3.3 0.00153292 0 0.00153284 0 0.00153294 3.3 0.0015328599999999998 3.3 0.0015329599999999999 0 0.00153288 0 0.00153298 3.3 0.0015329 3.3 0.001533 0 0.00153292 0 0.00153302 3.3 0.00153294 3.3 0.00153304 0 0.0015329599999999999 0 0.00153306 3.3 0.00153298 3.3 0.00153308 0 0.0015329999999999999 0 0.0015331 3.3 0.00153302 3.3 0.00153312 0 0.0015330399999999998 0 0.00153314 3.3 0.00153306 3.3 0.00153316 0 0.0015330799999999998 0 0.0015331799999999999 3.3 0.0015331 3.3 0.0015332 0 0.00153312 0 0.00153322 3.3 0.00153314 3.3 0.00153324 0 0.00153316 0 0.00153326 3.3 0.0015331799999999999 3.3 0.00153328 0 0.0015332 0 0.0015333 3.3 0.0015332199999999999 3.3 0.00153332 0 0.00153324 0 0.00153334 3.3 0.0015332599999999998 3.3 0.0015333599999999999 0 0.00153328 0 0.00153338 3.3 0.0015332999999999998 3.3 0.0015333999999999999 0 0.00153332 0 0.00153342 3.3 0.00153334 3.3 0.00153344 0 0.0015333599999999999 0 0.00153346 3.3 0.00153338 3.3 0.00153348 0 0.0015333999999999999 0 0.0015335 3.3 0.00153342 3.3 0.00153352 0 0.0015334399999999998 0 0.00153354 3.3 0.00153346 3.3 0.00153356 0 0.0015334799999999998 0 0.0015335799999999999 3.3 0.0015335 3.3 0.0015336 0 0.0015335199999999998 0 0.0015336199999999999 3.3 0.00153354 3.3 0.00153364 0 0.00153356 0 0.00153366 3.3 0.0015335799999999999 3.3 0.00153368 0 0.0015336 0 0.0015337 3.3 0.0015336199999999999 3.3 0.00153372 0 0.00153364 0 0.00153374 3.3 0.0015336599999999998 3.3 0.00153376 0 0.00153368 0 0.00153378 3.3 0.0015336999999999998 3.3 0.0015337999999999999 0 0.00153372 0 0.00153382 3.3 0.00153374 3.3 0.00153384 0 0.00153376 0 0.00153386 3.3 0.00153378 3.3 0.00153388 0 0.0015337999999999999 0 0.0015339 3.3 0.00153382 3.3 0.00153392 0 0.0015338399999999999 0 0.00153394 3.3 0.00153386 3.3 0.00153396 0 0.0015338799999999998 0 0.00153398 3.3 0.0015339 3.3 0.001534 0 0.0015339199999999998 0 0.0015340199999999999 3.3 0.00153394 3.3 0.00153404 0 0.00153396 0 0.00153406 3.3 0.00153398 3.3 0.00153408 0 0.001534 0 0.0015341 3.3 0.0015340199999999999 3.3 0.00153412 0 0.00153404 0 0.00153414 3.3 0.0015340599999999999 3.3 0.00153416 0 0.00153408 0 0.00153418 3.3 0.0015340999999999998 3.3 0.0015341999999999999 0 0.00153412 0 0.00153422 3.3 0.0015341399999999998 3.3 0.0015342399999999999 0 0.00153416 0 0.00153426 3.3 0.00153418 3.3 0.00153428 0 0.0015341999999999999 0 0.0015343 3.3 0.00153422 3.3 0.00153432 0 0.0015342399999999999 0 0.00153434 3.3 0.00153426 3.3 0.00153436 0 0.0015342799999999998 0 0.00153438 3.3 0.0015343 3.3 0.0015344 0 0.0015343199999999998 0 0.0015344199999999999 3.3 0.00153434 3.3 0.00153444 0 0.00153436 0 0.00153446 3.3 0.00153438 3.3 0.00153448 0 0.0015344 0 0.0015345 3.3 0.0015344199999999999 3.3 0.00153452 0 0.00153444 0 0.00153454 3.3 0.0015344599999999999 3.3 0.00153456 0 0.00153448 0 0.00153458 3.3 0.0015344999999999998 3.3 0.0015346 0 0.00153452 0 0.00153462 3.3 0.0015345399999999998 3.3 0.0015346399999999999 0 0.00153456 0 0.00153466 3.3 0.00153458 3.3 0.00153468 0 0.0015346 0 0.0015347 3.3 0.00153462 3.3 0.00153472 0 0.0015346399999999999 0 0.00153474 3.3 0.00153466 3.3 0.00153476 0 0.0015346799999999999 0 0.00153478 3.3 0.0015347 3.3 0.0015348 0 0.0015347199999999998 0 0.0015348199999999999 3.3 0.00153474 3.3 0.00153484 0 0.0015347599999999998 0 0.0015348599999999999 3.3 0.00153478 3.3 0.00153488 0 0.0015348 0 0.0015349 3.3 0.0015348199999999999 3.3 0.00153492 0 0.00153484 0 0.00153494 3.3 0.0015348599999999999 3.3 0.00153496 0 0.00153488 0 0.00153498 3.3 0.0015348999999999998 3.3 0.001535 0 0.00153492 0 0.00153502 3.3 0.0015349399999999998 3.3 0.0015350399999999999 0 0.00153496 0 0.00153506 3.3 0.0015349799999999998 3.3 0.0015350799999999999 0 0.001535 0 0.0015351 3.3 0.00153502 3.3 0.00153512 0 0.0015350399999999999 0 0.00153514 3.3 0.00153506 3.3 0.00153516 0 0.0015350799999999999 0 0.00153518 3.3 0.0015351 3.3 0.0015352 0 0.0015351199999999998 0 0.00153522 3.3 0.00153514 3.3 0.00153524 0 0.0015351599999999998 0 0.0015352599999999999 3.3 0.00153518 3.3 0.00153528 0 0.0015352 0 0.0015353 3.3 0.00153522 3.3 0.00153532 0 0.00153524 0 0.00153534 3.3 0.0015352599999999999 3.3 0.00153536 0 0.00153528 0 0.00153538 3.3 0.0015352999999999999 3.3 0.0015354 0 0.00153532 0 0.00153542 3.3 0.0015353399999999998 3.3 0.00153544 0 0.00153536 0 0.00153546 3.3 0.0015353799999999998 3.3 0.0015354799999999999 0 0.0015354 0 0.0015355 3.3 0.00153542 3.3 0.00153552 0 0.00153544 0 0.00153554 3.3 0.00153546 3.3 0.00153556 0 0.0015354799999999999 0 0.00153558 3.3 0.0015355 3.3 0.0015356 0 0.0015355199999999999 0 0.00153562 3.3 0.00153554 3.3 0.00153564 0 0.0015355599999999998 0 0.0015356599999999999 3.3 0.00153558 3.3 0.00153568 0 0.0015355999999999998 0 0.0015356999999999999 3.3 0.00153562 3.3 0.00153572 0 0.00153564 0 0.00153574 3.3 0.0015356599999999999 3.3 0.00153576 0 0.00153568 0 0.00153578 3.3 0.0015356999999999999 3.3 0.0015358 0 0.00153572 0 0.00153582 3.3 0.0015357399999999998 3.3 0.00153584 0 0.00153576 0 0.00153586 3.3 0.0015357799999999998 3.3 0.0015358799999999999 0 0.0015358 0 0.0015359 3.3 0.0015358199999999998 3.3 0.0015359199999999999 0 0.00153584 0 0.00153594 3.3 0.00153586 3.3 0.00153596 0 0.0015358799999999999 0 0.00153598 3.3 0.0015359 3.3 0.001536 0 0.0015359199999999999 0 0.00153602 3.3 0.00153594 3.3 0.00153604 0 0.0015359599999999998 0 0.00153606 3.3 0.00153598 3.3 0.00153608 0 0.0015359999999999998 0 0.0015360999999999999 3.3 0.00153602 3.3 0.00153612 0 0.00153604 0 0.00153614 3.3 0.00153606 3.3 0.00153616 0 0.00153608 0 0.00153618 3.3 0.0015360999999999999 3.3 0.0015362 0 0.00153612 0 0.00153622 3.3 0.0015361399999999999 3.3 0.00153624 0 0.00153616 0 0.00153626 3.3 0.0015361799999999998 3.3 0.00153628 0 0.0015362 0 0.0015363 3.3 0.0015362199999999998 3.3 0.0015363199999999999 0 0.00153624 0 0.00153634 3.3 0.00153626 3.3 0.00153636 0 0.00153628 0 0.00153638 3.3 0.0015363 3.3 0.0015364 0 0.0015363199999999999 0 0.00153642 3.3 0.00153634 3.3 0.00153644 0 0.0015363599999999999 0 0.00153646 3.3 0.00153638 3.3 0.00153648 0 0.0015363999999999998 0 0.0015364999999999999 3.3 0.00153642 3.3 0.00153652 0 0.0015364399999999998 0 0.0015365399999999999 3.3 0.00153646 3.3 0.00153656 0 0.00153648 0 0.00153658 3.3 0.0015364999999999999 3.3 0.0015366 0 0.00153652 0 0.00153662 3.3 0.0015365399999999999 3.3 0.00153664 0 0.00153656 0 0.00153666 3.3 0.0015365799999999998 3.3 0.00153668 0 0.0015366 0 0.0015367 3.3 0.0015366199999999998 3.3 0.0015367199999999999 0 0.00153664 0 0.00153674 3.3 0.0015366599999999998 3.3 0.0015367599999999999 0 0.00153668 0 0.00153678 3.3 0.0015367 3.3 0.0015368 0 0.0015367199999999999 0 0.00153682 3.3 0.00153674 3.3 0.00153684 0 0.0015367599999999999 0 0.00153686 3.3 0.00153678 3.3 0.00153688 0 0.0015367999999999998 0 0.0015369 3.3 0.00153682 3.3 0.00153692 0 0.0015368399999999998 0 0.0015369399999999999 3.3 0.00153686 3.3 0.00153696 0 0.00153688 0 0.00153698 3.3 0.0015369 3.3 0.001537 0 0.00153692 0 0.00153702 3.3 0.0015369399999999999 3.3 0.00153704 0 0.00153696 0 0.00153706 3.3 0.0015369799999999999 3.3 0.00153708 0 0.001537 0 0.0015371 3.3 0.0015370199999999998 3.3 0.00153712 0 0.00153704 0 0.00153714 3.3 0.0015370599999999998 3.3 0.0015371599999999999 0 0.00153708 0 0.00153718 3.3 0.0015371 3.3 0.0015372 0 0.00153712 0 0.00153722 3.3 0.00153714 3.3 0.00153724 0 0.0015371599999999999 0 0.00153726 3.3 0.00153718 3.3 0.00153728 0 0.0015371999999999999 0 0.0015373 3.3 0.00153722 3.3 0.00153732 0 0.0015372399999999998 0 0.0015373399999999999 3.3 0.00153726 3.3 0.00153736 0 0.0015372799999999998 0 0.0015373799999999999 3.3 0.0015373 3.3 0.0015374 0 0.00153732 0 0.00153742 3.3 0.0015373399999999999 3.3 0.00153744 0 0.00153736 0 0.00153746 3.3 0.0015373799999999999 3.3 0.00153748 0 0.0015374 0 0.0015375 3.3 0.0015374199999999998 3.3 0.00153752 0 0.00153744 0 0.00153754 3.3 0.0015374599999999998 3.3 0.0015375599999999999 0 0.00153748 0 0.00153758 3.3 0.0015374999999999998 3.3 0.0015375999999999999 0 0.00153752 0 0.00153762 3.3 0.00153754 3.3 0.00153764 0 0.0015375599999999999 0 0.00153766 3.3 0.00153758 3.3 0.00153768 0 0.0015375999999999999 0 0.0015377 3.3 0.00153762 3.3 0.00153772 0 0.0015376399999999998 0 0.00153774 3.3 0.00153766 3.3 0.00153776 0 0.0015376799999999998 0 0.0015377799999999999 3.3 0.0015377 3.3 0.0015378 0 0.00153772 0 0.00153782 3.3 0.00153774 3.3 0.00153784 0 0.00153776 0 0.00153786 3.3 0.0015377799999999999 3.3 0.00153788 0 0.0015378 0 0.0015379 3.3 0.0015378199999999999 3.3 0.00153792 0 0.00153784 0 0.00153794 3.3 0.0015378599999999998 3.3 0.0015379599999999999 0 0.00153788 0 0.00153798 3.3 0.0015378999999999998 3.3 0.0015379999999999999 0 0.00153792 0 0.00153802 3.3 0.00153794 3.3 0.00153804 0 0.0015379599999999999 0 0.00153806 3.3 0.00153798 3.3 0.00153808 0 0.0015379999999999999 0 0.0015381 3.3 0.00153802 3.3 0.00153812 0 0.0015380399999999998 0 0.00153814 3.3 0.00153806 3.3 0.00153816 0 0.0015380799999999998 0 0.0015381799999999999 3.3 0.0015381 3.3 0.0015382 0 0.0015381199999999998 0 0.0015382199999999999 3.3 0.00153814 3.3 0.00153824 0 0.00153816 0 0.00153826 3.3 0.0015381799999999999 3.3 0.00153828 0 0.0015382 0 0.0015383 3.3 0.0015382199999999999 3.3 0.00153832 0 0.00153824 0 0.00153834 3.3 0.0015382599999999998 3.3 0.00153836 0 0.00153828 0 0.00153838 3.3 0.0015382999999999998 3.3 0.0015383999999999999 0 0.00153832 0 0.00153842 3.3 0.00153834 3.3 0.00153844 0 0.00153836 0 0.00153846 3.3 0.00153838 3.3 0.00153848 0 0.0015383999999999999 0 0.0015385 3.3 0.00153842 3.3 0.00153852 0 0.0015384399999999999 0 0.00153854 3.3 0.00153846 3.3 0.00153856 0 0.0015384799999999998 0 0.00153858 3.3 0.0015385 3.3 0.0015386 0 0.0015385199999999998 0 0.0015386199999999999 3.3 0.00153854 3.3 0.00153864 0 0.00153856 0 0.00153866 3.3 0.00153858 3.3 0.00153868 0 0.0015386 0 0.0015387 3.3 0.0015386199999999999 3.3 0.00153872 0 0.00153864 0 0.00153874 3.3 0.0015386599999999999 3.3 0.00153876 0 0.00153868 0 0.00153878 3.3 0.0015386999999999998 3.3 0.0015387999999999999 0 0.00153872 0 0.00153882 3.3 0.0015387399999999998 3.3 0.0015388399999999999 0 0.00153876 0 0.00153886 3.3 0.00153878 3.3 0.00153888 0 0.0015387999999999999 0 0.0015389 3.3 0.00153882 3.3 0.00153892 0 0.0015388399999999999 0 0.00153894 3.3 0.00153886 3.3 0.00153896 0 0.0015388799999999998 0 0.00153898 3.3 0.0015389 3.3 0.001539 0 0.0015389199999999998 0 0.0015390199999999999 3.3 0.00153894 3.3 0.00153904 0 0.0015389599999999998 0 0.0015390599999999999 3.3 0.00153898 3.3 0.00153908 0 0.001539 0 0.0015391 3.3 0.0015390199999999999 3.3 0.00153912 0 0.00153904 0 0.00153914 3.3 0.0015390599999999999 3.3 0.00153916 0 0.00153908 0 0.00153918 3.3 0.0015390999999999998 3.3 0.0015392 0 0.00153912 0 0.00153922 3.3 0.0015391399999999998 3.3 0.0015392399999999999 0 0.00153916 0 0.00153926 3.3 0.00153918 3.3 0.00153928 0 0.0015392 0 0.0015393 3.3 0.00153922 3.3 0.00153932 0 0.0015392399999999999 0 0.00153934 3.3 0.00153926 3.3 0.00153936 0 0.0015392799999999999 0 0.00153938 3.3 0.0015393 3.3 0.0015394 0 0.0015393199999999998 0 0.00153942 3.3 0.00153934 3.3 0.00153944 0 0.0015393599999999998 0 0.0015394599999999999 3.3 0.00153938 3.3 0.00153948 0 0.0015394 0 0.0015395 3.3 0.00153942 3.3 0.00153952 0 0.00153944 0 0.00153954 3.3 0.0015394599999999999 3.3 0.00153956 0 0.00153948 0 0.00153958 3.3 0.0015394999999999999 3.3 0.0015396 0 0.00153952 0 0.00153962 3.3 0.0015395399999999998 3.3 0.0015396399999999999 0 0.00153956 0 0.00153966 3.3 0.0015395799999999998 3.3 0.0015396799999999999 0 0.0015396 0 0.0015397 3.3 0.00153962 3.3 0.00153972 0 0.0015396399999999999 0 0.00153974 3.3 0.00153966 3.3 0.00153976 0 0.0015396799999999999 0 0.00153978 3.3 0.0015397 3.3 0.0015398 0 0.0015397199999999998 0 0.00153982 3.3 0.00153974 3.3 0.00153984 0 0.0015397599999999998 0 0.0015398599999999999 3.3 0.00153978 3.3 0.00153988 0 0.0015397999999999998 0 0.0015398999999999999 3.3 0.00153982 3.3 0.00153992 0 0.00153984 0 0.00153994 3.3 0.0015398599999999999 3.3 0.00153996 0 0.00153988 0 0.00153998 3.3 0.0015398999999999999 3.3 0.00154 0 0.00153992 0 0.00154002 3.3 0.0015399399999999998 3.3 0.00154004 0 0.00153996 0 0.00154006 3.3 0.0015399799999999998 3.3 0.0015400799999999999 0 0.00154 0 0.0015401 3.3 0.00154002 3.3 0.00154012 0 0.00154004 0 0.00154014 3.3 0.00154006 3.3 0.00154016 0 0.0015400799999999999 0 0.00154018 3.3 0.0015401 3.3 0.0015402 0 0.0015401199999999999 0 0.00154022 3.3 0.00154014 3.3 0.00154024 0 0.0015401599999999998 0 0.00154026 3.3 0.00154018 3.3 0.00154028 0 0.0015401999999999998 0 0.0015402999999999999 3.3 0.00154022 3.3 0.00154032 0 0.00154024 0 0.00154034 3.3 0.00154026 3.3 0.00154036 0 0.00154028 0 0.00154038 3.3 0.0015402999999999999 3.3 0.0015404 0 0.00154032 0 0.00154042 3.3 0.0015403399999999999 3.3 0.00154044 0 0.00154036 0 0.00154046 3.3 0.0015403799999999998 3.3 0.0015404799999999999 0 0.0015404 0 0.0015405 3.3 0.0015404199999999998 3.3 0.0015405199999999999 0 0.00154044 0 0.00154054 3.3 0.00154046 3.3 0.00154056 0 0.0015404799999999999 0 0.00154058 3.3 0.0015405 3.3 0.0015406 0 0.0015405199999999999 0 0.00154062 3.3 0.00154054 3.3 0.00154064 0 0.0015405599999999998 0 0.00154066 3.3 0.00154058 3.3 0.00154068 0 0.0015405999999999998 0 0.0015406999999999999 3.3 0.00154062 3.3 0.00154072 0 0.0015406399999999998 0 0.0015407399999999999 3.3 0.00154066 3.3 0.00154076 0 0.00154068 0 0.00154078 3.3 0.0015406999999999999 3.3 0.0015408 0 0.00154072 0 0.00154082 3.3 0.0015407399999999999 3.3 0.00154084 0 0.00154076 0 0.00154086 3.3 0.0015407799999999998 3.3 0.00154088 0 0.0015408 0 0.0015409 3.3 0.0015408199999999998 3.3 0.0015409199999999999 0 0.00154084 0 0.00154094 3.3 0.00154086 3.3 0.00154096 0 0.00154088 0 0.00154098 3.3 0.0015409 3.3 0.001541 0 0.0015409199999999999 0 0.00154102 3.3 0.00154094 3.3 0.00154104 0 0.0015409599999999999 0 0.00154106 3.3 0.00154098 3.3 0.00154108 0 0.0015409999999999998 0 0.0015411 3.3 0.00154102 3.3 0.00154112 0 0.0015410399999999998 0 0.0015411399999999999 3.3 0.00154106 3.3 0.00154116 0 0.00154108 0 0.00154118 3.3 0.0015411 3.3 0.0015412 0 0.00154112 0 0.00154122 3.3 0.0015411399999999999 3.3 0.00154124 0 0.00154116 0 0.00154126 3.3 0.0015411799999999999 3.3 0.00154128 0 0.0015412 0 0.0015413 3.3 0.0015412199999999998 3.3 0.0015413199999999999 0 0.00154124 0 0.00154134 3.3 0.0015412599999999998 3.3 0.0015413599999999999 0 0.00154128 0 0.00154138 3.3 0.0015413 3.3 0.0015414 0 0.0015413199999999999 0 0.00154142 3.3 0.00154134 3.3 0.00154144 0 0.0015413599999999999 0 0.00154146 3.3 0.00154138 3.3 0.00154148 0 0.0015413999999999998 0 0.0015415 3.3 0.00154142 3.3 0.00154152 0 0.0015414399999999998 0 0.0015415399999999999 3.3 0.00154146 3.3 0.00154156 0 0.00154148 0 0.00154158 3.3 0.0015415 3.3 0.0015416 0 0.00154152 0 0.00154162 3.3 0.0015415399999999999 3.3 0.00154164 0 0.00154156 0 0.00154166 3.3 0.0015415799999999999 3.3 0.00154168 0 0.0015416 0 0.0015417 3.3 0.0015416199999999998 3.3 0.00154172 0 0.00154164 0 0.00154174 3.3 0.0015416599999999998 3.3 0.0015417599999999999 0 0.00154168 0 0.00154178 3.3 0.0015417 3.3 0.0015418 0 0.00154172 0 0.00154182 3.3 0.00154174 3.3 0.00154184 0 0.0015417599999999999 0 0.00154186 3.3 0.00154178 3.3 0.00154188 0 0.0015417999999999999 0 0.0015419 3.3 0.00154182 3.3 0.00154192 0 0.0015418399999999998 0 0.0015419399999999999 3.3 0.00154186 3.3 0.00154196 0 0.0015418799999999998 0 0.0015419799999999999 3.3 0.0015419 3.3 0.001542 0 0.00154192 0 0.00154202 3.3 0.0015419399999999999 3.3 0.00154204 0 0.00154196 0 0.00154206 3.3 0.0015419799999999999 3.3 0.00154208 0 0.001542 0 0.0015421 3.3 0.0015420199999999998 3.3 0.00154212 0 0.00154204 0 0.00154214 3.3 0.0015420599999999998 3.3 0.0015421599999999999 0 0.00154208 0 0.00154218 3.3 0.0015420999999999998 3.3 0.0015421999999999999 0 0.00154212 0 0.00154222 3.3 0.00154214 3.3 0.00154224 0 0.0015421599999999999 0 0.00154226 3.3 0.00154218 3.3 0.00154228 0 0.0015421999999999999 0 0.0015423 3.3 0.00154222 3.3 0.00154232 0 0.0015422399999999998 0 0.00154234 3.3 0.00154226 3.3 0.00154236 0 0.0015422799999999998 0 0.0015423799999999999 3.3 0.0015423 3.3 0.0015424 0 0.00154232 0 0.00154242 3.3 0.00154234 3.3 0.00154244 0 0.00154236 0 0.00154246 3.3 0.0015423799999999999 3.3 0.00154248 0 0.0015424 0 0.0015425 3.3 0.0015424199999999999 3.3 0.00154252 0 0.00154244 0 0.00154254 3.3 0.0015424599999999998 3.3 0.00154256 0 0.00154248 0 0.00154258 3.3 0.0015424999999999998 3.3 0.0015425999999999999 0 0.00154252 0 0.00154262 3.3 0.00154254 3.3 0.00154264 0 0.00154256 0 0.00154266 3.3 0.00154258 3.3 0.00154268 0 0.0015425999999999999 0 0.0015427 3.3 0.00154262 3.3 0.00154272 0 0.0015426399999999999 0 0.00154274 3.3 0.00154266 3.3 0.00154276 0 0.0015426799999999998 0 0.0015427799999999999 3.3 0.0015427 3.3 0.0015428 0 0.0015427199999999998 0 0.0015428199999999999 3.3 0.00154274 3.3 0.00154284 0 0.00154276 0 0.00154286 3.3 0.0015427799999999999 3.3 0.00154288 0 0.0015428 0 0.0015429 3.3 0.0015428199999999999 3.3 0.00154292 0 0.00154284 0 0.00154294 3.3 0.0015428599999999998 3.3 0.00154296 0 0.00154288 0 0.00154298 3.3 0.0015428999999999998 3.3 0.0015429999999999999 0 0.00154292 0 0.00154302 3.3 0.0015429399999999998 3.3 0.0015430399999999999 0 0.00154296 0 0.00154306 3.3 0.00154298 3.3 0.00154308 0 0.0015429999999999999 0 0.0015431 3.3 0.00154302 3.3 0.00154312 0 0.0015430399999999999 0 0.00154314 3.3 0.00154306 3.3 0.00154316 0 0.0015430799999999998 0 0.00154318 3.3 0.0015431 3.3 0.0015432 0 0.0015431199999999998 0 0.0015432199999999999 3.3 0.00154314 3.3 0.00154324 0 0.00154316 0 0.00154326 3.3 0.00154318 3.3 0.00154328 0 0.0015432 0 0.0015433 3.3 0.0015432199999999999 3.3 0.00154332 0 0.00154324 0 0.00154334 3.3 0.0015432599999999999 3.3 0.00154336 0 0.00154328 0 0.00154338 3.3 0.0015432999999999998 3.3 0.0015434 0 0.00154332 0 0.00154342 3.3 0.0015433399999999998 3.3 0.0015434399999999999 0 0.00154336 0 0.00154346 3.3 0.00154338 3.3 0.00154348 0 0.0015434 0 0.0015435 3.3 0.00154342 3.3 0.00154352 0 0.0015434399999999999 0 0.00154354 3.3 0.00154346 3.3 0.00154356 0 0.0015434799999999999 0 0.00154358 3.3 0.0015435 3.3 0.0015436 0 0.0015435199999999998 0 0.0015436199999999999 3.3 0.00154354 3.3 0.00154364 0 0.0015435599999999998 0 0.0015436599999999999 3.3 0.00154358 3.3 0.00154368 0 0.0015436 0 0.0015437 3.3 0.0015436199999999999 3.3 0.00154372 0 0.00154364 0 0.00154374 3.3 0.0015436599999999999 3.3 0.00154376 0 0.00154368 0 0.00154378 3.3 0.0015436999999999998 3.3 0.0015438 0 0.00154372 0 0.00154382 3.3 0.0015437399999999998 3.3 0.0015438399999999999 0 0.00154376 0 0.00154386 3.3 0.0015437799999999998 3.3 0.0015438799999999999 0 0.0015438 0 0.0015439 3.3 0.00154382 3.3 0.00154392 0 0.0015438399999999999 0 0.00154394 3.3 0.00154386 3.3 0.00154396 0 0.0015438799999999999 0 0.00154398 3.3 0.0015439 3.3 0.001544 0 0.0015439199999999998 0 0.00154402 3.3 0.00154394 3.3 0.00154404 0 0.0015439599999999998 0 0.0015440599999999999 3.3 0.00154398 3.3 0.00154408 0 0.001544 0 0.0015441 3.3 0.00154402 3.3 0.00154412 0 0.00154404 0 0.00154414 3.3 0.0015440599999999999 3.3 0.00154416 0 0.00154408 0 0.00154418 3.3 0.0015440999999999999 3.3 0.0015442 0 0.00154412 0 0.00154422 3.3 0.0015441399999999998 3.3 0.00154424 0 0.00154416 0 0.00154426 3.3 0.0015441799999999998 3.3 0.0015442799999999999 0 0.0015442 0 0.0015443 3.3 0.00154422 3.3 0.00154432 0 0.00154424 0 0.00154434 3.3 0.00154426 3.3 0.00154436 0 0.0015442799999999999 0 0.00154438 3.3 0.0015443 3.3 0.0015444 0 0.0015443199999999999 0 0.00154442 3.3 0.00154434 3.3 0.00154444 0 0.0015443599999999998 0 0.0015444599999999999 3.3 0.00154438 3.3 0.00154448 0 0.0015443999999999998 0 0.0015444999999999999 3.3 0.00154442 3.3 0.00154452 0 0.00154444 0 0.00154454 3.3 0.0015444599999999999 3.3 0.00154456 0 0.00154448 0 0.00154458 3.3 0.0015444999999999999 3.3 0.0015446 0 0.00154452 0 0.00154462 3.3 0.0015445399999999998 3.3 0.00154464 0 0.00154456 0 0.00154466 3.3 0.0015445799999999998 3.3 0.0015446799999999999 0 0.0015446 0 0.0015447 3.3 0.0015446199999999998 3.3 0.0015447199999999999 0 0.00154464 0 0.00154474 3.3 0.00154466 3.3 0.00154476 0 0.0015446799999999999 0 0.00154478 3.3 0.0015447 3.3 0.0015448 0 0.0015447199999999999 0 0.00154482 3.3 0.00154474 3.3 0.00154484 0 0.0015447599999999998 0 0.00154486 3.3 0.00154478 3.3 0.00154488 0 0.0015447999999999998 0 0.0015448999999999999 3.3 0.00154482 3.3 0.00154492 0 0.00154484 0 0.00154494 3.3 0.00154486 3.3 0.00154496 0 0.00154488 0 0.00154498 3.3 0.0015448999999999999 3.3 0.001545 0 0.00154492 0 0.00154502 3.3 0.0015449399999999999 3.3 0.00154504 0 0.00154496 0 0.00154506 3.3 0.0015449799999999998 3.3 0.0015450799999999999 0 0.001545 0 0.0015451 3.3 0.0015450199999999998 3.3 0.0015451199999999999 0 0.00154504 0 0.00154514 3.3 0.00154506 3.3 0.00154516 0 0.0015450799999999999 0 0.00154518 3.3 0.0015451 3.3 0.0015452 0 0.0015451199999999999 0 0.00154522 3.3 0.00154514 3.3 0.00154524 0 0.0015451599999999998 0 0.00154526 3.3 0.00154518 3.3 0.00154528 0 0.0015451999999999998 0 0.0015452999999999999 3.3 0.00154522 3.3 0.00154532 0 0.0015452399999999998 0 0.0015453399999999999 3.3 0.00154526 3.3 0.00154536 0 0.00154528 0 0.00154538 3.3 0.0015452999999999999 3.3 0.0015454 0 0.00154532 0 0.00154542 3.3 0.0015453399999999999 3.3 0.00154544 0 0.00154536 0 0.00154546 3.3 0.0015453799999999998 3.3 0.00154548 0 0.0015454 0 0.0015455 3.3 0.0015454199999999998 3.3 0.0015455199999999999 0 0.00154544 0 0.00154554 3.3 0.00154546 3.3 0.00154556 0 0.00154548 0 0.00154558 3.3 0.0015455 3.3 0.0015456 0 0.0015455199999999999 0 0.00154562 3.3 0.00154554 3.3 0.00154564 0 0.0015455599999999999 0 0.00154566 3.3 0.00154558 3.3 0.00154568 0 0.0015455999999999998 0 0.0015457 3.3 0.00154562 3.3 0.00154572 0 0.0015456399999999998 0 0.0015457399999999999 3.3 0.00154566 3.3 0.00154576 0 0.00154568 0 0.00154578 3.3 0.0015457 3.3 0.0015458 0 0.00154572 0 0.00154582 3.3 0.0015457399999999999 3.3 0.00154584 0 0.00154576 0 0.00154586 3.3 0.0015457799999999999 3.3 0.00154588 0 0.0015458 0 0.0015459 3.3 0.0015458199999999998 3.3 0.0015459199999999999 0 0.00154584 0 0.00154594 3.3 0.0015458599999999998 3.3 0.0015459599999999999 0 0.00154588 0 0.00154598 3.3 0.0015459 3.3 0.001546 0 0.0015459199999999999 0 0.00154602 3.3 0.00154594 3.3 0.00154604 0 0.0015459599999999999 0 0.00154606 3.3 0.00154598 3.3 0.00154608 0 0.0015459999999999998 0 0.0015461 3.3 0.00154602 3.3 0.00154612 0 0.0015460399999999998 0 0.0015461399999999999 3.3 0.00154606 3.3 0.00154616 0 0.0015460799999999998 0 0.0015461799999999999 3.3 0.0015461 3.3 0.0015462 0 0.00154612 0 0.00154622 3.3 0.0015461399999999999 3.3 0.00154624 0 0.00154616 0 0.00154626 3.3 0.0015461799999999999 3.3 0.00154628 0 0.0015462 0 0.0015463 3.3 0.0015462199999999998 3.3 0.00154632 0 0.00154624 0 0.00154634 3.3 0.0015462599999999998 3.3 0.0015463599999999999 0 0.00154628 0 0.00154638 3.3 0.0015463 3.3 0.0015464 0 0.00154632 0 0.00154642 3.3 0.00154634 3.3 0.00154644 0 0.0015463599999999999 0 0.00154646 3.3 0.00154638 3.3 0.00154648 0 0.0015463999999999999 0 0.0015465 3.3 0.00154642 3.3 0.00154652 0 0.0015464399999999998 0 0.00154654 3.3 0.00154646 3.3 0.00154656 0 0.0015464799999999998 0 0.0015465799999999999 3.3 0.0015465 3.3 0.0015466 0 0.00154652 0 0.00154662 3.3 0.00154654 3.3 0.00154664 0 0.00154656 0 0.00154666 3.3 0.0015465799999999999 3.3 0.00154668 0 0.0015466 0 0.0015467 3.3 0.0015466199999999999 3.3 0.00154672 0 0.00154664 0 0.00154674 3.3 0.0015466599999999998 3.3 0.0015467599999999999 0 0.00154668 0 0.00154678 3.3 0.0015466999999999998 3.3 0.0015467999999999999 0 0.00154672 0 0.00154682 3.3 0.00154674 3.3 0.00154684 0 0.0015467599999999999 0 0.00154686 3.3 0.00154678 3.3 0.00154688 0 0.0015467999999999999 0 0.0015469 3.3 0.00154682 3.3 0.00154692 0 0.0015468399999999998 0 0.00154694 3.3 0.00154686 3.3 0.00154696 0 0.0015468799999999998 0 0.0015469799999999999 3.3 0.0015469 3.3 0.001547 0 0.0015469199999999998 0 0.0015470199999999999 3.3 0.00154694 3.3 0.00154704 0 0.00154696 0 0.00154706 3.3 0.0015469799999999999 3.3 0.00154708 0 0.001547 0 0.0015471 3.3 0.0015470199999999999 3.3 0.00154712 0 0.00154704 0 0.00154714 3.3 0.0015470599999999998 3.3 0.00154716 0 0.00154708 0 0.00154718 3.3 0.0015470999999999998 3.3 0.0015471999999999999 0 0.00154712 0 0.00154722 3.3 0.00154714 3.3 0.00154724 0 0.00154716 0 0.00154726 3.3 0.00154718 3.3 0.00154728 0 0.0015471999999999999 0 0.0015473 3.3 0.00154722 3.3 0.00154732 0 0.0015472399999999999 0 0.00154734 3.3 0.00154726 3.3 0.00154736 0 0.0015472799999999998 0 0.00154738 3.3 0.0015473 3.3 0.0015474 0 0.0015473199999999998 0 0.0015474199999999999 3.3 0.00154734 3.3 0.00154744 0 0.00154736 0 0.00154746 3.3 0.00154738 3.3 0.00154748 0 0.0015474 0 0.0015475 3.3 0.0015474199999999999 3.3 0.00154752 0 0.00154744 0 0.00154754 3.3 0.0015474599999999999 3.3 0.00154756 0 0.00154748 0 0.00154758 3.3 0.0015474999999999998 3.3 0.0015475999999999999 0 0.00154752 0 0.00154762 3.3 0.0015475399999999998 3.3 0.0015476399999999999 0 0.00154756 0 0.00154766 3.3 0.00154758 3.3 0.00154768 0 0.0015475999999999999 0 0.0015477 3.3 0.00154762 3.3 0.00154772 0 0.0015476399999999999 0 0.00154774 3.3 0.00154766 3.3 0.00154776 0 0.0015476799999999998 0 0.00154778 3.3 0.0015477 3.3 0.0015478 0 0.0015477199999999998 0 0.0015478199999999999 3.3 0.00154774 3.3 0.00154784 0 0.0015477599999999998 0 0.0015478599999999999 3.3 0.00154778 3.3 0.00154788 0 0.0015478 0 0.0015479 3.3 0.0015478199999999999 3.3 0.00154792 0 0.00154784 0 0.00154794 3.3 0.0015478599999999999 3.3 0.00154796 0 0.00154788 0 0.00154798 3.3 0.0015478999999999998 3.3 0.001548 0 0.00154792 0 0.00154802 3.3 0.0015479399999999998 3.3 0.0015480399999999999 0 0.00154796 0 0.00154806 3.3 0.00154798 3.3 0.00154808 0 0.001548 0 0.0015481 3.3 0.00154802 3.3 0.00154812 0 0.0015480399999999999 0 0.00154814 3.3 0.00154806 3.3 0.00154816 0 0.0015480799999999999 0 0.00154818 3.3 0.0015481 3.3 0.0015482 0 0.0015481199999999998 0 0.0015482199999999999 3.3 0.00154814 3.3 0.00154824 0 0.0015481599999999998 0 0.0015482599999999999 3.3 0.00154818 3.3 0.00154828 0 0.0015482 0 0.0015483 3.3 0.0015482199999999999 3.3 0.00154832 0 0.00154824 0 0.00154834 3.3 0.0015482599999999999 3.3 0.00154836 0 0.00154828 0 0.00154838 3.3 0.0015482999999999998 3.3 0.0015484 0 0.00154832 0 0.00154842 3.3 0.0015483399999999998 3.3 0.0015484399999999999 0 0.00154836 0 0.00154846 3.3 0.0015483799999999998 3.3 0.0015484799999999999 0 0.0015484 0 0.0015485 3.3 0.00154842 3.3 0.00154852 0 0.0015484399999999999 0 0.00154854 3.3 0.00154846 3.3 0.00154856 0 0.0015484799999999999 0 0.00154858 3.3 0.0015485 3.3 0.0015486 0 0.0015485199999999998 0 0.00154862 3.3 0.00154854 3.3 0.00154864 0 0.0015485599999999998 0 0.0015486599999999999 3.3 0.00154858 3.3 0.00154868 0 0.0015486 0 0.0015487 3.3 0.00154862 3.3 0.00154872 0 0.00154864 0 0.00154874 3.3 0.0015486599999999999 3.3 0.00154876 0 0.00154868 0 0.00154878 3.3 0.0015486999999999999 3.3 0.0015488 0 0.00154872 0 0.00154882 3.3 0.0015487399999999998 3.3 0.00154884 0 0.00154876 0 0.00154886 3.3 0.0015487799999999998 3.3 0.0015488799999999999 0 0.0015488 0 0.0015489 3.3 0.00154882 3.3 0.00154892 0 0.00154884 0 0.00154894 3.3 0.00154886 3.3 0.00154896 0 0.0015488799999999999 0 0.00154898 3.3 0.0015489 3.3 0.001549 0 0.0015489199999999999 0 0.00154902 3.3 0.00154894 3.3 0.00154904 0 0.0015489599999999998 0 0.0015490599999999999 3.3 0.00154898 3.3 0.00154908 0 0.0015489999999999998 0 0.0015490999999999999 3.3 0.00154902 3.3 0.00154912 0 0.00154904 0 0.00154914 3.3 0.0015490599999999999 3.3 0.00154916 0 0.00154908 0 0.00154918 3.3 0.0015490999999999999 3.3 0.0015492 0 0.00154912 0 0.00154922 3.3 0.0015491399999999998 3.3 0.00154924 0 0.00154916 0 0.00154926 3.3 0.0015491799999999998 3.3 0.0015492799999999999 0 0.0015492 0 0.0015493 3.3 0.0015492199999999998 3.3 0.0015493199999999999 0 0.00154924 0 0.00154934 3.3 0.00154926 3.3 0.00154936 0 0.0015492799999999999 0 0.00154938 3.3 0.0015493 3.3 0.0015494 0 0.0015493199999999999 0 0.00154942 3.3 0.00154934 3.3 0.00154944 0 0.0015493599999999998 0 0.00154946 3.3 0.00154938 3.3 0.00154948 0 0.0015493999999999998 0 0.0015494999999999999 3.3 0.00154942 3.3 0.00154952 0 0.00154944 0 0.00154954 3.3 0.00154946 3.3 0.00154956 0 0.00154948 0 0.00154958 3.3 0.0015494999999999999 3.3 0.0015496 0 0.00154952 0 0.00154962 3.3 0.0015495399999999999 3.3 0.00154964 0 0.00154956 0 0.00154966 3.3 0.0015495799999999998 3.3 0.00154968 0 0.0015496 0 0.0015497 3.3 0.0015496199999999998 3.3 0.0015497199999999999 0 0.00154964 0 0.00154974 3.3 0.00154966 3.3 0.00154976 0 0.00154968 0 0.00154978 3.3 0.0015497 3.3 0.0015498 0 0.0015497199999999999 0 0.00154982 3.3 0.00154974 3.3 0.00154984 0 0.0015497599999999999 0 0.00154986 3.3 0.00154978 3.3 0.00154988 0 0.0015497999999999998 0 0.0015498999999999999 3.3 0.00154982 3.3 0.00154992 0 0.0015498399999999998 0 0.0015499399999999999 3.3 0.00154986 3.3 0.00154996 0 0.00154988 0 0.00154998 3.3 0.0015498999999999999 3.3 0.00155 0 0.00154992 0 0.00155002 3.3 0.0015499399999999999 3.3 0.00155004 0 0.00154996 0 0.00155006 3.3 0.0015499799999999998 3.3 0.00155008 0 0.00155 0 0.0015501 3.3 0.0015500199999999998 3.3 0.0015501199999999999 0 0.00155004 0 0.00155014 3.3 0.0015500599999999998 3.3 0.0015501599999999999 0 0.00155008 0 0.00155018 3.3 0.0015501 3.3 0.0015502 0 0.0015501199999999999 0 0.00155022 3.3 0.00155014 3.3 0.00155024 0 0.0015501599999999999 0 0.00155026 3.3 0.00155018 3.3 0.00155028 0 0.0015501999999999998 0 0.0015503 3.3 0.00155022 3.3 0.00155032 0 0.0015502399999999998 0 0.0015503399999999999 3.3 0.00155026 3.3 0.00155036 0 0.00155028 0 0.00155038 3.3 0.0015503 3.3 0.0015504 0 0.00155032 0 0.00155042 3.3 0.0015503399999999999 3.3 0.00155044 0 0.00155036 0 0.00155046 3.3 0.0015503799999999999 3.3 0.00155048 0 0.0015504 0 0.0015505 3.3 0.0015504199999999998 3.3 0.00155052 0 0.00155044 0 0.00155054 3.3 0.0015504599999999998 3.3 0.0015505599999999999 0 0.00155048 0 0.00155058 3.3 0.0015505 3.3 0.0015506 0 0.00155052 0 0.00155062 3.3 0.00155054 3.3 0.00155064 0 0.0015505599999999999 0 0.00155066 3.3 0.00155058 3.3 0.00155068 0 0.0015505999999999999 0 0.0015507 3.3 0.00155062 3.3 0.00155072 0 0.0015506399999999998 0 0.0015507399999999999 3.3 0.00155066 3.3 0.00155076 0 0.0015506799999999998 0 0.0015507799999999999 3.3 0.0015507 3.3 0.0015508 0 0.00155072 0 0.00155082 3.3 0.0015507399999999999 3.3 0.00155084 0 0.00155076 0 0.00155086 3.3 0.0015507799999999999 3.3 0.00155088 0 0.0015508 0 0.0015509 3.3 0.0015508199999999998 3.3 0.00155092 0 0.00155084 0 0.00155094 3.3 0.0015508599999999998 3.3 0.0015509599999999999 0 0.00155088 0 0.00155098 3.3 0.0015508999999999998 3.3 0.0015509999999999999 0 0.00155092 0 0.00155102 3.3 0.00155094 3.3 0.00155104 0 0.0015509599999999999 0 0.00155106 3.3 0.00155098 3.3 0.00155108 0 0.0015509999999999999 0 0.0015511 3.3 0.00155102 3.3 0.00155112 0 0.0015510399999999998 0 0.00155114 3.3 0.00155106 3.3 0.00155116 0 0.0015510799999999998 0 0.0015511799999999999 3.3 0.0015511 3.3 0.0015512 0 0.00155112 0 0.00155122 3.3 0.00155114 3.3 0.00155124 0 0.00155116 0 0.00155126 3.3 0.0015511799999999999 3.3 0.00155128 0 0.0015512 0 0.0015513 3.3 0.0015512199999999999 3.3 0.00155132 0 0.00155124 0 0.00155134 3.3 0.0015512599999999998 3.3 0.00155136 0 0.00155128 0 0.00155138 3.3 0.0015512999999999998 3.3 0.0015513999999999999 0 0.00155132 0 0.00155142 3.3 0.00155134 3.3 0.00155144 0 0.00155136 0 0.00155146 3.3 0.00155138 3.3 0.00155148 0 0.0015513999999999999 0 0.0015515 3.3 0.00155142 3.3 0.00155152 0 0.0015514399999999999 0 0.00155154 3.3 0.00155146 3.3 0.00155156 0 0.0015514799999999998 0 0.0015515799999999999 3.3 0.0015515 3.3 0.0015516 0 0.0015515199999999998 0 0.0015516199999999999 3.3 0.00155154 3.3 0.00155164 0 0.00155156 0 0.00155166 3.3 0.0015515799999999999 3.3 0.00155168 0 0.0015516 0 0.0015517 3.3 0.0015516199999999999 3.3 0.00155172 0 0.00155164 0 0.00155174 3.3 0.0015516599999999998 3.3 0.00155176 0 0.00155168 0 0.00155178 3.3 0.0015516999999999998 3.3 0.0015517999999999999 0 0.00155172 0 0.00155182 3.3 0.00155174 3.3 0.00155184 0 0.00155176 0 0.00155186 3.3 0.00155178 3.3 0.00155188 0 0.0015517999999999999 0 0.0015519 3.3 0.00155182 3.3 0.00155192 0 0.0015518399999999999 0 0.00155194 3.3 0.00155186 3.3 0.00155196 0 0.0015518799999999998 0 0.00155198 3.3 0.0015519 3.3 0.001552 0 0.0015519199999999998 0 0.0015520199999999999 3.3 0.00155194 3.3 0.00155204 0 0.00155196 0 0.00155206 3.3 0.00155198 3.3 0.00155208 0 0.001552 0 0.0015521 3.3 0.0015520199999999999 3.3 0.00155212 0 0.00155204 0 0.00155214 3.3 0.0015520599999999999 3.3 0.00155216 0 0.00155208 0 0.00155218 3.3 0.0015520999999999998 3.3 0.0015521999999999999 0 0.00155212 0 0.00155222 3.3 0.0015521399999999998 3.3 0.0015522399999999999 0 0.00155216 0 0.00155226 3.3 0.00155218 3.3 0.00155228 0 0.0015521999999999999 0 0.0015523 3.3 0.00155222 3.3 0.00155232 0 0.0015522399999999999 0 0.00155234 3.3 0.00155226 3.3 0.00155236 0 0.0015522799999999998 0 0.00155238 3.3 0.0015523 3.3 0.0015524 0 0.0015523199999999998 0 0.0015524199999999999 3.3 0.00155234 3.3 0.00155244 0 0.0015523599999999998 0 0.0015524599999999999 3.3 0.00155238 3.3 0.00155248 0 0.0015524 0 0.0015525 3.3 0.0015524199999999999 3.3 0.00155252 0 0.00155244 0 0.00155254 3.3 0.0015524599999999999 3.3 0.00155256 0 0.00155248 0 0.00155258 3.3 0.0015524999999999998 3.3 0.0015526 0 0.00155252 0 0.00155262 3.3 0.0015525399999999998 3.3 0.0015526399999999999 0 0.00155256 0 0.00155266 3.3 0.00155258 3.3 0.00155268 0 0.0015526 0 0.0015527 3.3 0.00155262 3.3 0.00155272 0 0.0015526399999999999 0 0.00155274 3.3 0.00155266 3.3 0.00155276 0 0.0015526799999999999 0 0.00155278 3.3 0.0015527 3.3 0.0015528 0 0.0015527199999999998 0 0.00155282 3.3 0.00155274 3.3 0.00155284 0 0.0015527599999999998 0 0.0015528599999999999 3.3 0.00155278 3.3 0.00155288 0 0.0015528 0 0.0015529 3.3 0.00155282 3.3 0.00155292 0 0.00155284 0 0.00155294 3.3 0.0015528599999999999 3.3 0.00155296 0 0.00155288 0 0.00155298 3.3 0.0015528999999999999 3.3 0.001553 0 0.00155292 0 0.00155302 3.3 0.0015529399999999998 3.3 0.0015530399999999999 0 0.00155296 0 0.00155306 3.3 0.0015529799999999998 3.3 0.0015530799999999999 0 0.001553 0 0.0015531 3.3 0.00155302 3.3 0.00155312 0 0.0015530399999999999 0 0.00155314 3.3 0.00155306 3.3 0.00155316 0 0.0015530799999999999 0 0.00155318 3.3 0.0015531 3.3 0.0015532 0 0.0015531199999999998 0 0.00155322 3.3 0.00155314 3.3 0.00155324 0 0.0015531599999999998 0 0.0015532599999999999 3.3 0.00155318 3.3 0.00155328 0 0.0015531999999999998 0 0.0015532999999999999 3.3 0.00155322 3.3 0.00155332 0 0.00155324 0 0.00155334 3.3 0.0015532599999999999 3.3 0.00155336 0 0.00155328 0 0.00155338 3.3 0.0015532999999999999 3.3 0.0015534 0 0.00155332 0 0.00155342 3.3 0.0015533399999999998 3.3 0.00155344 0 0.00155336 0 0.00155346 3.3 0.0015533799999999998 3.3 0.0015534799999999999 0 0.0015534 0 0.0015535 3.3 0.00155342 3.3 0.00155352 0 0.00155344 0 0.00155354 3.3 0.00155346 3.3 0.00155356 0 0.0015534799999999999 0 0.00155358 3.3 0.0015535 3.3 0.0015536 0 0.0015535199999999999 0 0.00155362 3.3 0.00155354 3.3 0.00155364 0 0.0015535599999999998 0 0.00155366 3.3 0.00155358 3.3 0.00155368 0 0.0015535999999999998 0 0.0015536999999999999 3.3 0.00155362 3.3 0.00155372 0 0.00155364 0 0.00155374 3.3 0.00155366 3.3 0.00155376 0 0.00155368 0 0.00155378 3.3 0.0015536999999999999 3.3 0.0015538 0 0.00155372 0 0.00155382 3.3 0.0015537399999999999 3.3 0.00155384 0 0.00155376 0 0.00155386 3.3 0.0015537799999999998 3.3 0.0015538799999999999 0 0.0015538 0 0.0015539 3.3 0.0015538199999999998 3.3 0.0015539199999999999 0 0.00155384 0 0.00155394 3.3 0.00155386 3.3 0.00155396 0 0.0015538799999999999 0 0.00155398 3.3 0.0015539 3.3 0.001554 0 0.0015539199999999999 0 0.00155402 3.3 0.00155394 3.3 0.00155404 0 0.0015539599999999998 0 0.00155406 3.3 0.00155398 3.3 0.00155408 0 0.0015539999999999998 0 0.0015540999999999999 3.3 0.00155402 3.3 0.00155412 0 0.0015540399999999998 0 0.0015541399999999999 3.3 0.00155406 3.3 0.00155416 0 0.00155408 0 0.00155418 3.3 0.0015540999999999999 3.3 0.0015542 0 0.00155412 0 0.00155422 3.3 0.0015541399999999999 3.3 0.00155424 0 0.00155416 0 0.00155426 3.3 0.0015541799999999998 3.3 0.00155428 0 0.0015542 0 0.0015543 3.3 0.0015542199999999998 3.3 0.0015543199999999999 0 0.00155424 0 0.00155434 3.3 0.00155426 3.3 0.00155436 0 0.00155428 0 0.00155438 3.3 0.0015543 3.3 0.0015544 0 0.0015543199999999999 0 0.00155442 3.3 0.00155434 3.3 0.00155444 0 0.0015543599999999999 0 0.00155446 3.3 0.00155438 3.3 0.00155448 0 0.0015543999999999998 0 0.0015545 3.3 0.00155442 3.3 0.00155452 0 0.0015544399999999998 0 0.0015545399999999999 3.3 0.00155446 3.3 0.00155456 0 0.00155448 0 0.00155458 3.3 0.0015545 3.3 0.0015546 0 0.00155452 0 0.00155462 3.3 0.0015545399999999999 3.3 0.00155464 0 0.00155456 0 0.00155466 3.3 0.0015545799999999999 3.3 0.00155468 0 0.0015546 0 0.0015547 3.3 0.0015546199999999998 3.3 0.0015547199999999999 0 0.00155464 0 0.00155474 3.3 0.0015546599999999998 3.3 0.0015547599999999999 0 0.00155468 0 0.00155478 3.3 0.0015547 3.3 0.0015548 0 0.0015547199999999999 0 0.00155482 3.3 0.00155474 3.3 0.00155484 0 0.0015547599999999999 0 0.00155486 3.3 0.00155478 3.3 0.00155488 0 0.0015547999999999998 0 0.0015549 3.3 0.00155482 3.3 0.00155492 0 0.0015548399999999998 0 0.0015549399999999999 3.3 0.00155486 3.3 0.00155496 0 0.0015548799999999998 0 0.0015549799999999999 3.3 0.0015549 3.3 0.001555 0 0.00155492 0 0.00155502 3.3 0.0015549399999999999 3.3 0.00155504 0 0.00155496 0 0.00155506 3.3 0.0015549799999999999 3.3 0.00155508 0 0.001555 0 0.0015551 3.3 0.0015550199999999998 3.3 0.00155512 0 0.00155504 0 0.00155514 3.3 0.0015550599999999998 3.3 0.0015551599999999999 0 0.00155508 0 0.00155518 3.3 0.0015551 3.3 0.0015552 0 0.00155512 0 0.00155522 3.3 0.00155514 3.3 0.00155524 0 0.0015551599999999999 0 0.00155526 3.3 0.00155518 3.3 0.00155528 0 0.0015551999999999999 0 0.0015553 3.3 0.00155522 3.3 0.00155532 0 0.0015552399999999998 0 0.0015553399999999999 3.3 0.00155526 3.3 0.00155536 0 0.0015552799999999998 0 0.0015553799999999999 3.3 0.0015553 3.3 0.0015554 0 0.00155532 0 0.00155542 3.3 0.0015553399999999999 3.3 0.00155544 0 0.00155536 0 0.00155546 3.3 0.0015553799999999999 3.3 0.00155548 0 0.0015554 0 0.0015555 3.3 0.0015554199999999998 3.3 0.00155552 0 0.00155544 0 0.00155554 3.3 0.0015554599999999998 3.3 0.0015555599999999999 0 0.00155548 0 0.00155558 3.3 0.0015554999999999998 3.3 0.0015555999999999999 0 0.00155552 0 0.00155562 3.3 0.00155554 3.3 0.00155564 0 0.0015555599999999999 0 0.00155566 3.3 0.00155558 3.3 0.00155568 0 0.0015555999999999999 0 0.0015557 3.3 0.00155562 3.3 0.00155572 0 0.0015556399999999998 0 0.00155574 3.3 0.00155566 3.3 0.00155576 0 0.0015556799999999998 0 0.0015557799999999999 3.3 0.0015557 3.3 0.0015558 0 0.00155572 0 0.00155582 3.3 0.00155574 3.3 0.00155584 0 0.00155576 0 0.00155586 3.3 0.0015557799999999999 3.3 0.00155588 0 0.0015558 0 0.0015559 3.3 0.0015558199999999999 3.3 0.00155592 0 0.00155584 0 0.00155594 3.3 0.0015558599999999998 3.3 0.00155596 0 0.00155588 0 0.00155598 3.3 0.0015558999999999998 3.3 0.0015559999999999999 0 0.00155592 0 0.00155602 3.3 0.00155594 3.3 0.00155604 0 0.00155596 0 0.00155606 3.3 0.00155598 3.3 0.00155608 0 0.0015559999999999999 0 0.0015561 3.3 0.00155602 3.3 0.00155612 0 0.0015560399999999999 0 0.00155614 3.3 0.00155606 3.3 0.00155616 0 0.0015560799999999998 0 0.0015561799999999999 3.3 0.0015561 3.3 0.0015562 0 0.0015561199999999998 0 0.0015562199999999999 3.3 0.00155614 3.3 0.00155624 0 0.00155616 0 0.00155626 3.3 0.0015561799999999999 3.3 0.00155628 0 0.0015562 0 0.0015563 3.3 0.0015562199999999999 3.3 0.00155632 0 0.00155624 0 0.00155634 3.3 0.0015562599999999998 3.3 0.00155636 0 0.00155628 0 0.00155638 3.3 0.0015562999999999998 3.3 0.0015563999999999999 0 0.00155632 0 0.00155642 3.3 0.0015563399999999998 3.3 0.0015564399999999999 0 0.00155636 0 0.00155646 3.3 0.00155638 3.3 0.00155648 0 0.0015563999999999999 0 0.0015565 3.3 0.00155642 3.3 0.00155652 0 0.0015564399999999999 0 0.00155654 3.3 0.00155646 3.3 0.00155656 0 0.0015564799999999998 0 0.00155658 3.3 0.0015565 3.3 0.0015566 0 0.0015565199999999998 0 0.0015566199999999999 3.3 0.00155654 3.3 0.00155664 0 0.00155656 0 0.00155666 3.3 0.00155658 3.3 0.00155668 0 0.0015566 0 0.0015567 3.3 0.0015566199999999999 3.3 0.00155672 0 0.00155664 0 0.00155674 3.3 0.0015566599999999999 3.3 0.00155676 0 0.00155668 0 0.00155678 3.3 0.0015566999999999998 3.3 0.0015568 0 0.00155672 0 0.00155682 3.3 0.0015567399999999998 3.3 0.0015568399999999999 0 0.00155676 0 0.00155686 3.3 0.00155678 3.3 0.00155688 0 0.0015568 0 0.0015569 3.3 0.00155682 3.3 0.00155692 0 0.0015568399999999999 0 0.00155694 3.3 0.00155686 3.3 0.00155696 0 0.0015568799999999999 0 0.00155698 3.3 0.0015569 3.3 0.001557 0 0.0015569199999999998 0 0.0015570199999999999 3.3 0.00155694 3.3 0.00155704 0 0.0015569599999999998 0 0.0015570599999999999 3.3 0.00155698 3.3 0.00155708 0 0.001557 0 0.0015571 3.3 0.0015570199999999999 3.3 0.00155712 0 0.00155704 0 0.00155714 3.3 0.0015570599999999999 3.3 0.00155716 0 0.00155708 0 0.00155718 3.3 0.0015570999999999998 3.3 0.0015572 0 0.00155712 0 0.00155722 3.3 0.0015571399999999998 3.3 0.0015572399999999999 0 0.00155716 0 0.00155726 3.3 0.0015571799999999998 3.3 0.0015572799999999999 0 0.0015572 0 0.0015573 3.3 0.00155722 3.3 0.00155732 0 0.0015572399999999999 0 0.00155734 3.3 0.00155726 3.3 0.00155736 0 0.0015572799999999999 0 0.00155738 3.3 0.0015573 3.3 0.0015574 0 0.0015573199999999998 0 0.00155742 3.3 0.00155734 3.3 0.00155744 0 0.0015573599999999998 0 0.0015574599999999999 3.3 0.00155738 3.3 0.00155748 0 0.0015574 0 0.0015575 3.3 0.00155742 3.3 0.00155752 0 0.00155744 0 0.00155754 3.3 0.0015574599999999999 3.3 0.00155756 0 0.00155748 0 0.00155758 3.3 0.0015574999999999999 3.3 0.0015576 0 0.00155752 0 0.00155762 3.3 0.0015575399999999998 3.3 0.00155764 0 0.00155756 0 0.00155766 3.3 0.0015575799999999998 3.3 0.0015576799999999999 0 0.0015576 0 0.0015577 3.3 0.00155762 3.3 0.00155772 0 0.00155764 0 0.00155774 3.3 0.00155766 3.3 0.00155776 0 0.0015576799999999999 0 0.00155778 3.3 0.0015577 3.3 0.0015578 0 0.0015577199999999999 0 0.00155782 3.3 0.00155774 3.3 0.00155784 0 0.0015577599999999998 0 0.0015578599999999999 3.3 0.00155778 3.3 0.00155788 0 0.0015577999999999998 0 0.0015578999999999999 3.3 0.00155782 3.3 0.00155792 0 0.00155784 0 0.00155794 3.3 0.0015578599999999999 3.3 0.00155796 0 0.00155788 0 0.00155798 3.3 0.0015578999999999999 3.3 0.001558 0 0.00155792 0 0.00155802 3.3 0.0015579399999999998 3.3 0.00155804 0 0.00155796 0 0.00155806 3.3 0.0015579799999999998 3.3 0.0015580799999999999 0 0.001558 0 0.0015581 3.3 0.0015580199999999998 3.3 0.0015581199999999999 0 0.00155804 0 0.00155814 3.3 0.00155806 3.3 0.00155816 0 0.0015580799999999999 0 0.00155818 3.3 0.0015581 3.3 0.0015582 0 0.0015581199999999999 0 0.00155822 3.3 0.00155814 3.3 0.00155824 0 0.0015581599999999998 0 0.00155826 3.3 0.00155818 3.3 0.00155828 0 0.0015581999999999998 0 0.0015582999999999999 3.3 0.00155822 3.3 0.00155832 0 0.00155824 0 0.00155834 3.3 0.00155826 3.3 0.00155836 0 0.00155828 0 0.00155838 3.3 0.0015582999999999999 3.3 0.0015584 0 0.00155832 0 0.00155842 3.3 0.0015583399999999999 3.3 0.00155844 0 0.00155836 0 0.00155846 3.3 0.0015583799999999998 3.3 0.0015584799999999999 0 0.0015584 0 0.0015585 3.3 0.0015584199999999998 3.3 0.0015585199999999999 0 0.00155844 0 0.00155854 3.3 0.00155846 3.3 0.00155856 0 0.0015584799999999999 0 0.00155858 3.3 0.0015585 3.3 0.0015586 0 0.0015585199999999999 0 0.00155862 3.3 0.00155854 3.3 0.00155864 0 0.0015585599999999999 0 0.00155866 3.3 0.00155858 3.3 0.00155868 0 0.0015585999999999998 0 0.0015586999999999999 3.3 0.00155862 3.3 0.00155872 0 0.0015586399999999998 0 0.0015587399999999999 3.3 0.00155866 3.3 0.00155876 0 0.00155868 0 0.00155878 3.3 0.0015586999999999999 3.3 0.0015588 0 0.00155872 0 0.00155882 3.3 0.0015587399999999999 3.3 0.00155884 0 0.00155876 0 0.00155886 3.3 0.0015587799999999998 3.3 0.00155888 0 0.0015588 0 0.0015589 3.3 0.0015588199999999998 3.3 0.0015589199999999999 0 0.00155884 0 0.00155894 3.3 0.00155886 3.3 0.00155896 0 0.00155888 0 0.00155898 3.3 0.0015589 3.3 0.001559 0 0.0015589199999999999 0 0.00155902 3.3 0.00155894 3.3 0.00155904 0 0.0015589599999999999 0 0.00155906 3.3 0.00155898 3.3 0.00155908 0 0.0015589999999999998 0 0.0015591 3.3 0.00155902 3.3 0.00155912 0 0.0015590399999999998 0 0.0015591399999999999 3.3 0.00155906 3.3 0.00155916 0 0.00155908 0 0.00155918 3.3 0.0015591 3.3 0.0015592 0 0.00155912 0 0.00155922 3.3 0.0015591399999999999 3.3 0.00155924 0 0.00155916 0 0.00155926 3.3 0.0015591799999999999 3.3 0.00155928 0 0.0015592 0 0.0015593 3.3 0.0015592199999999998 3.3 0.0015593199999999999 0 0.00155924 0 0.00155934 3.3 0.0015592599999999998 3.3 0.0015593599999999999 0 0.00155928 0 0.00155938 3.3 0.0015593 3.3 0.0015594 0 0.0015593199999999999 0 0.00155942 3.3 0.00155934 3.3 0.00155944 0 0.0015593599999999999 0 0.00155946 3.3 0.00155938 3.3 0.00155948 0 0.0015593999999999998 0 0.0015595 3.3 0.00155942 3.3 0.00155952 0 0.0015594399999999998 0 0.0015595399999999999 3.3 0.00155946 3.3 0.00155956 0 0.0015594799999999998 0 0.0015595799999999999 3.3 0.0015595 3.3 0.0015596 0 0.00155952 0 0.00155962 3.3 0.0015595399999999999 3.3 0.00155964 0 0.00155956 0 0.00155966 3.3 0.0015595799999999999 3.3 0.00155968 0 0.0015596 0 0.0015597 3.3 0.0015596199999999998 3.3 0.00155972 0 0.00155964 0 0.00155974 3.3 0.0015596599999999998 3.3 0.0015597599999999999 0 0.00155968 0 0.00155978 3.3 0.0015597 3.3 0.0015598 0 0.00155972 0 0.00155982 3.3 0.00155974 3.3 0.00155984 0 0.0015597599999999999 0 0.00155986 3.3 0.00155978 3.3 0.00155988 0 0.0015597999999999999 0 0.0015599 3.3 0.00155982 3.3 0.00155992 0 0.0015598399999999998 0 0.00155994 3.3 0.00155986 3.3 0.00155996 0 0.0015598799999999998 0 0.0015599799999999999 3.3 0.0015599 3.3 0.00156 0 0.00155992 0 0.00156002 3.3 0.00155994 3.3 0.00156004 0 0.00155996 0 0.00156006 3.3 0.0015599799999999999 3.3 0.00156008 0 0.00156 0 0.0015601 3.3 0.0015600199999999999 3.3 0.00156012 0 0.00156004 0 0.00156014 3.3 0.0015600599999999998 3.3 0.0015601599999999999 0 0.00156008 0 0.00156018 3.3 0.0015600999999999998 3.3 0.0015601999999999999 0 0.00156012 0 0.00156022 3.3 0.00156014 3.3 0.00156024 0 0.0015601599999999999 0 0.00156026 3.3 0.00156018 3.3 0.00156028 0 0.0015601999999999999 0 0.0015603 3.3 0.00156022 3.3 0.00156032 0 0.0015602399999999998 0 0.00156034 3.3 0.00156026 3.3 0.00156036 0 0.0015602799999999998 0 0.0015603799999999999 3.3 0.0015603 3.3 0.0015604 0 0.0015603199999999998 0 0.0015604199999999999 3.3 0.00156034 3.3 0.00156044 0 0.00156036 0 0.00156046 3.3 0.0015603799999999999 3.3 0.00156048 0 0.0015604 0 0.0015605 3.3 0.0015604199999999999 3.3 0.00156052 0 0.00156044 0 0.00156054 3.3 0.0015604599999999998 3.3 0.00156056 0 0.00156048 0 0.00156058 3.3 0.0015604999999999998 3.3 0.0015605999999999999 0 0.00156052 0 0.00156062 3.3 0.00156054 3.3 0.00156064 0 0.00156056 0 0.00156066 3.3 0.00156058 3.3 0.00156068 0 0.0015605999999999999 0 0.0015607 3.3 0.00156062 3.3 0.00156072 0 0.0015606399999999999 0 0.00156074 3.3 0.00156066 3.3 0.00156076 0 0.0015606799999999998 0 0.00156078 3.3 0.0015607 3.3 0.0015608 0 0.0015607199999999998 0 0.0015608199999999999 3.3 0.00156074 3.3 0.00156084 0 0.00156076 0 0.00156086 3.3 0.00156078 3.3 0.00156088 0 0.0015608 0 0.0015609 3.3 0.0015608199999999999 3.3 0.00156092 0 0.00156084 0 0.00156094 3.3 0.0015608599999999999 3.3 0.00156096 0 0.00156088 0 0.00156098 3.3 0.0015608999999999998 3.3 0.0015609999999999999 0 0.00156092 0 0.00156102 3.3 0.0015609399999999998 3.3 0.0015610399999999999 0 0.00156096 0 0.00156106 3.3 0.00156098 3.3 0.00156108 0 0.0015609999999999999 0 0.0015611 3.3 0.00156102 3.3 0.00156112 0 0.0015610399999999999 0 0.00156114 3.3 0.00156106 3.3 0.00156116 0 0.0015610799999999998 0 0.00156118 3.3 0.0015611 3.3 0.0015612 0 0.0015611199999999998 0 0.0015612199999999999 3.3 0.00156114 3.3 0.00156124 0 0.0015611599999999998 0 0.0015612599999999999 3.3 0.00156118 3.3 0.00156128 0 0.0015612 0 0.0015613 3.3 0.0015612199999999999 3.3 0.00156132 0 0.00156124 0 0.00156134 3.3 0.0015612599999999999 3.3 0.00156136 0 0.00156128 0 0.00156138 3.3 0.0015612999999999998 3.3 0.0015614 0 0.00156132 0 0.00156142 3.3 0.0015613399999999998 3.3 0.0015614399999999999 0 0.00156136 0 0.00156146 3.3 0.00156138 3.3 0.00156148 0 0.0015614 0 0.0015615 3.3 0.00156142 3.3 0.00156152 0 0.0015614399999999999 0 0.00156154 3.3 0.00156146 3.3 0.00156156 0 0.0015614799999999999 0 0.00156158 3.3 0.0015615 3.3 0.0015616 0 0.0015615199999999998 0 0.00156162 3.3 0.00156154 3.3 0.00156164 0 0.0015615599999999998 0 0.0015616599999999999 3.3 0.00156158 3.3 0.00156168 0 0.0015616 0 0.0015617 3.3 0.00156162 3.3 0.00156172 0 0.00156164 0 0.00156174 3.3 0.0015616599999999999 3.3 0.00156176 0 0.00156168 0 0.00156178 3.3 0.0015616999999999999 3.3 0.0015618 0 0.00156172 0 0.00156182 3.3 0.0015617399999999998 3.3 0.0015618399999999999 0 0.00156176 0 0.00156186 3.3 0.0015617799999999998 3.3 0.0015618799999999999 0 0.0015618 0 0.0015619 3.3 0.00156182 3.3 0.00156192 0 0.0015618399999999999 0 0.00156194 3.3 0.00156186 3.3 0.00156196 0 0.0015618799999999999 0 0.00156198 3.3 0.0015619 3.3 0.001562 0 0.0015619199999999998 0 0.00156202 3.3 0.00156194 3.3 0.00156204 0 0.0015619599999999998 0 0.0015620599999999999 3.3 0.00156198 3.3 0.00156208 0 0.0015619999999999998 0 0.0015620999999999999 3.3 0.00156202 3.3 0.00156212 0 0.00156204 0 0.00156214 3.3 0.0015620599999999999 3.3 0.00156216 0 0.00156208 0 0.00156218 3.3 0.0015620999999999999 3.3 0.0015622 0 0.00156212 0 0.00156222 3.3 0.0015621399999999998 3.3 0.00156224 0 0.00156216 0 0.00156226 3.3 0.0015621799999999998 3.3 0.0015622799999999999 0 0.0015622 0 0.0015623 3.3 0.00156222 3.3 0.00156232 0 0.00156224 0 0.00156234 3.3 0.00156226 3.3 0.00156236 0 0.0015622799999999999 0 0.00156238 3.3 0.0015623 3.3 0.0015624 0 0.0015623199999999999 0 0.00156242 3.3 0.00156234 3.3 0.00156244 0 0.0015623599999999998 0 0.0015624599999999999 3.3 0.00156238 3.3 0.00156248 0 0.0015623999999999998 0 0.0015624999999999999 3.3 0.00156242 3.3 0.00156252 0 0.00156244 0 0.00156254 3.3 0.0015624599999999999 3.3 0.00156256 0 0.00156248 0 0.00156258 3.3 0.0015624999999999999 3.3 0.0015626 0 0.00156252 0 0.00156262 3.3 0.0015625399999999998 3.3 0.00156264 0 0.00156256 0 0.00156266 3.3 0.0015625799999999998 3.3 0.0015626799999999999 0 0.0015626 0 0.0015627 3.3 0.0015626199999999998 3.3 0.0015627199999999999 0 0.00156264 0 0.00156274 3.3 0.00156266 3.3 0.00156276 0 0.0015626799999999999 0 0.00156278 3.3 0.0015627 3.3 0.0015628 0 0.0015627199999999999 0 0.00156282 3.3 0.00156274 3.3 0.00156284 0 0.0015627599999999998 0 0.00156286 3.3 0.00156278 3.3 0.00156288 0 0.0015627999999999998 0 0.0015628999999999999 3.3 0.00156282 3.3 0.00156292 0 0.00156284 0 0.00156294 3.3 0.00156286 3.3 0.00156296 0 0.00156288 0 0.00156298 3.3 0.0015628999999999999 3.3 0.001563 0 0.00156292 0 0.00156302 3.3 0.0015629399999999999 3.3 0.00156304 0 0.00156296 0 0.00156306 3.3 0.0015629799999999998 3.3 0.00156308 0 0.001563 0 0.0015631 3.3 0.0015630199999999998 3.3 0.0015631199999999999 0 0.00156304 0 0.00156314 3.3 0.00156306 3.3 0.00156316 0 0.00156308 0 0.00156318 3.3 0.0015631 3.3 0.0015632 0 0.0015631199999999999 0 0.00156322 3.3 0.00156314 3.3 0.00156324 0 0.0015631599999999999 0 0.00156326 3.3 0.00156318 3.3 0.00156328 0 0.0015631999999999998 0 0.0015632999999999999 3.3 0.00156322 3.3 0.00156332 0 0.0015632399999999998 0 0.0015633399999999999 3.3 0.00156326 3.3 0.00156336 0 0.00156328 0 0.00156338 3.3 0.0015632999999999999 3.3 0.0015634 0 0.00156332 0 0.00156342 3.3 0.0015633399999999999 3.3 0.00156344 0 0.00156336 0 0.00156346 3.3 0.0015633799999999998 3.3 0.00156348 0 0.0015634 0 0.0015635 3.3 0.0015634199999999998 3.3 0.0015635199999999999 0 0.00156344 0 0.00156354 3.3 0.0015634599999999998 3.3 0.0015635599999999999 0 0.00156348 0 0.00156358 3.3 0.0015635 3.3 0.0015636 0 0.0015635199999999999 0 0.00156362 3.3 0.00156354 3.3 0.00156364 0 0.0015635599999999999 0 0.00156366 3.3 0.00156358 3.3 0.00156368 0 0.0015635999999999998 0 0.0015637 3.3 0.00156362 3.3 0.00156372 0 0.0015636399999999998 0 0.0015637399999999999 3.3 0.00156366 3.3 0.00156376 0 0.00156368 0 0.00156378 3.3 0.0015637 3.3 0.0015638 0 0.00156372 0 0.00156382 3.3 0.0015637399999999999 3.3 0.00156384 0 0.00156376 0 0.00156386 3.3 0.0015637799999999999 3.3 0.00156388 0 0.0015638 0 0.0015639 3.3 0.0015638199999999998 3.3 0.00156392 0 0.00156384 0 0.00156394 3.3 0.0015638599999999998 3.3 0.0015639599999999999 0 0.00156388 0 0.00156398 3.3 0.0015639 3.3 0.001564 0 0.00156392 0 0.00156402 3.3 0.00156394 3.3 0.00156404 0 0.0015639599999999999 0 0.00156406 3.3 0.00156398 3.3 0.00156408 0 0.0015639999999999999 0 0.0015641 3.3 0.00156402 3.3 0.00156412 0 0.0015640399999999998 0 0.0015641399999999999 3.3 0.00156406 3.3 0.00156416 0 0.0015640799999999998 0 0.0015641799999999999 3.3 0.0015641 3.3 0.0015642 0 0.00156412 0 0.00156422 3.3 0.0015641399999999999 3.3 0.00156424 0 0.00156416 0 0.00156426 3.3 0.0015641799999999999 3.3 0.00156428 0 0.0015642 0 0.0015643 3.3 0.0015642199999999998 3.3 0.00156432 0 0.00156424 0 0.00156434 3.3 0.0015642599999999998 3.3 0.0015643599999999999 0 0.00156428 0 0.00156438 3.3 0.0015642999999999998 3.3 0.0015643999999999999 0 0.00156432 0 0.00156442 3.3 0.00156434 3.3 0.00156444 0 0.0015643599999999999 0 0.00156446 3.3 0.00156438 3.3 0.00156448 0 0.0015643999999999999 0 0.0015645 3.3 0.00156442 3.3 0.00156452 0 0.0015644399999999998 0 0.00156454 3.3 0.00156446 3.3 0.00156456 0 0.0015644799999999998 0 0.0015645799999999999 3.3 0.0015645 3.3 0.0015646 0 0.00156452 0 0.00156462 3.3 0.00156454 3.3 0.00156464 0 0.00156456 0 0.00156466 3.3 0.0015645799999999999 3.3 0.00156468 0 0.0015646 0 0.0015647 3.3 0.0015646199999999999 3.3 0.00156472 0 0.00156464 0 0.00156474 3.3 0.0015646599999999998 3.3 0.00156476 0 0.00156468 0 0.00156478 3.3 0.0015646999999999998 3.3 0.0015647999999999999 0 0.00156472 0 0.00156482 3.3 0.00156474 3.3 0.00156484 0 0.00156476 0 0.00156486 3.3 0.00156478 3.3 0.00156488 0 0.0015647999999999999 0 0.0015649 3.3 0.00156482 3.3 0.00156492 0 0.0015648399999999999 0 0.00156494 3.3 0.00156486 3.3 0.00156496 0 0.0015648799999999998 0 0.0015649799999999999 3.3 0.0015649 3.3 0.001565 0 0.0015649199999999998 0 0.0015650199999999999 3.3 0.00156494 3.3 0.00156504 0 0.00156496 0 0.00156506 3.3 0.0015649799999999999 3.3 0.00156508 0 0.001565 0 0.0015651 3.3 0.0015650199999999999 3.3 0.00156512 0 0.00156504 0 0.00156514 3.3 0.0015650599999999998 3.3 0.00156516 0 0.00156508 0 0.00156518 3.3 0.0015650999999999998 3.3 0.0015651999999999999 0 0.00156512 0 0.00156522 3.3 0.0015651399999999998 3.3 0.0015652399999999999 0 0.00156516 0 0.00156526 3.3 0.00156518 3.3 0.00156528 0 0.0015651999999999999 0 0.0015653 3.3 0.00156522 3.3 0.00156532 0 0.0015652399999999999 0 0.00156534 3.3 0.00156526 3.3 0.00156536 0 0.0015652799999999998 0 0.00156538 3.3 0.0015653 3.3 0.0015654 0 0.0015653199999999998 0 0.0015654199999999999 3.3 0.00156534 3.3 0.00156544 0 0.00156536 0 0.00156546 3.3 0.00156538 3.3 0.00156548 0 0.0015654 0 0.0015655 3.3 0.0015654199999999999 3.3 0.00156552 0 0.00156544 0 0.00156554 3.3 0.0015654599999999999 3.3 0.00156556 0 0.00156548 0 0.00156558 3.3 0.0015654999999999998 3.3 0.0015655999999999999 0 0.00156552 0 0.00156562 3.3 0.0015655399999999998 3.3 0.0015656399999999999 0 0.00156556 0 0.00156566 3.3 0.00156558 3.3 0.00156568 0 0.0015655999999999999 0 0.0015657 3.3 0.00156562 3.3 0.00156572 0 0.0015656399999999999 0 0.00156574 3.3 0.00156566 3.3 0.00156576 0 0.0015656799999999998 0 0.00156578 3.3 0.0015657 3.3 0.0015658 0 0.0015657199999999998 0 0.0015658199999999999 3.3 0.00156574 3.3 0.00156584 0 0.0015657599999999998 0 0.0015658599999999999 3.3 0.00156578 3.3 0.00156588 0 0.0015658 0 0.0015659 3.3 0.0015658199999999999 3.3 0.00156592 0 0.00156584 0 0.00156594 3.3 0.0015658599999999999 3.3 0.00156596 0 0.00156588 0 0.00156598 3.3 0.0015658999999999998 3.3 0.001566 0 0.00156592 0 0.00156602 3.3 0.0015659399999999998 3.3 0.0015660399999999999 0 0.00156596 0 0.00156606 3.3 0.00156598 3.3 0.00156608 0 0.001566 0 0.0015661 3.3 0.00156602 3.3 0.00156612 0 0.0015660399999999999 0 0.00156614 3.3 0.00156606 3.3 0.00156616 0 0.0015660799999999999 0 0.00156618 3.3 0.0015661 3.3 0.0015662 0 0.0015661199999999998 0 0.00156622 3.3 0.00156614 3.3 0.00156624 0 0.0015661599999999998 0 0.0015662599999999999 3.3 0.00156618 3.3 0.00156628 0 0.0015662 0 0.0015663 3.3 0.00156622 3.3 0.00156632 0 0.00156624 0 0.00156634 3.3 0.0015662599999999999 3.3 0.00156636 0 0.00156628 0 0.00156638 3.3 0.0015662999999999999 3.3 0.0015664 0 0.00156632 0 0.00156642 3.3 0.0015663399999999998 3.3 0.0015664399999999999 0 0.00156636 0 0.00156646 3.3 0.0015663799999999998 3.3 0.0015664799999999999 0 0.0015664 0 0.0015665 3.3 0.00156642 3.3 0.00156652 0 0.0015664399999999999 0 0.00156654 3.3 0.00156646 3.3 0.00156656 0 0.0015664799999999999 0 0.00156658 3.3 0.0015665 3.3 0.0015666 0 0.0015665199999999998 0 0.00156662 3.3 0.00156654 3.3 0.00156664 0 0.0015665599999999998 0 0.0015666599999999999 3.3 0.00156658 3.3 0.00156668 0 0.0015665999999999998 0 0.0015666999999999999 3.3 0.00156662 3.3 0.00156672 0 0.00156664 0 0.00156674 3.3 0.0015666599999999999 3.3 0.00156676 0 0.00156668 0 0.00156678 3.3 0.0015666999999999999 3.3 0.0015668 0 0.00156672 0 0.00156682 3.3 0.0015667399999999998 3.3 0.00156684 0 0.00156676 0 0.00156686 3.3 0.0015667799999999998 3.3 0.0015668799999999999 0 0.0015668 0 0.0015669 3.3 0.00156682 3.3 0.00156692 0 0.00156684 0 0.00156694 3.3 0.00156686 3.3 0.00156696 0 0.0015668799999999999 0 0.00156698 3.3 0.0015669 3.3 0.001567 0 0.0015669199999999999 0 0.00156702 3.3 0.00156694 3.3 0.00156704 0 0.0015669599999999998 0 0.00156706 3.3 0.00156698 3.3 0.00156708 0 0.0015669999999999998 0 0.0015670999999999999 3.3 0.00156702 3.3 0.00156712 0 0.00156704 0 0.00156714 3.3 0.00156706 3.3 0.00156716 0 0.00156708 0 0.00156718 3.3 0.0015670999999999999 3.3 0.0015672 0 0.00156712 0 0.00156722 3.3 0.0015671399999999999 3.3 0.00156724 0 0.00156716 0 0.00156726 3.3 0.0015671799999999998 3.3 0.0015672799999999999 0 0.0015672 0 0.0015673 3.3 0.0015672199999999998 3.3 0.0015673199999999999 0 0.00156724 0 0.00156734 3.3 0.00156726 3.3 0.00156736 0 0.0015672799999999999 0 0.00156738 3.3 0.0015673 3.3 0.0015674 0 0.0015673199999999999 0 0.00156742 3.3 0.00156734 3.3 0.00156744 0 0.0015673599999999998 0 0.00156746 3.3 0.00156738 3.3 0.00156748 0 0.0015673999999999998 0 0.0015674999999999999 3.3 0.00156742 3.3 0.00156752 0 0.0015674399999999998 0 0.0015675399999999999 3.3 0.00156746 3.3 0.00156756 0 0.00156748 0 0.00156758 3.3 0.0015674999999999999 3.3 0.0015676 0 0.00156752 0 0.00156762 3.3 0.0015675399999999999 3.3 0.00156764 0 0.00156756 0 0.00156766 3.3 0.0015675799999999998 3.3 0.00156768 0 0.0015676 0 0.0015677 3.3 0.0015676199999999998 3.3 0.0015677199999999999 0 0.00156764 0 0.00156774 3.3 0.00156766 3.3 0.00156776 0 0.00156768 0 0.00156778 3.3 0.0015677 3.3 0.0015678 0 0.0015677199999999999 0 0.00156782 3.3 0.00156774 3.3 0.00156784 0 0.0015677599999999999 0 0.00156786 3.3 0.00156778 3.3 0.00156788 0 0.0015677999999999998 0 0.0015679 3.3 0.00156782 3.3 0.00156792 0 0.0015678399999999998 0 0.0015679399999999999 3.3 0.00156786 3.3 0.00156796 0 0.00156788 0 0.00156798 3.3 0.0015679 3.3 0.001568 0 0.00156792 0 0.00156802 3.3 0.0015679399999999999 3.3 0.00156804 0 0.00156796 0 0.00156806 3.3 0.0015679799999999999 3.3 0.00156808 0 0.001568 0 0.0015681 3.3 0.0015680199999999998 3.3 0.0015681199999999999 0 0.00156804 0 0.00156814 3.3 0.0015680599999999998 3.3 0.0015681599999999999 0 0.00156808 0 0.00156818 3.3 0.0015681 3.3 0.0015682 0 0.0015681199999999999 0 0.00156822 3.3 0.00156814 3.3 0.00156824 0 0.0015681599999999999 0 0.00156826 3.3 0.00156818 3.3 0.00156828 0 0.0015681999999999998 0 0.0015683 3.3 0.00156822 3.3 0.00156832 0 0.0015682399999999998 0 0.0015683399999999999 3.3 0.00156826 3.3 0.00156836 0 0.0015682799999999998 0 0.0015683799999999999 3.3 0.0015683 3.3 0.0015684 0 0.00156832 0 0.00156842 3.3 0.0015683399999999999 3.3 0.00156844 0 0.00156836 0 0.00156846 3.3 0.0015683799999999999 3.3 0.00156848 0 0.0015684 0 0.0015685 3.3 0.0015684199999999998 3.3 0.00156852 0 0.00156844 0 0.00156854 3.3 0.0015684599999999998 3.3 0.0015685599999999999 0 0.00156848 0 0.00156858 3.3 0.0015685 3.3 0.0015686 0 0.00156852 0 0.00156862 3.3 0.00156854 3.3 0.00156864 0 0.0015685599999999999 0 0.00156866 3.3 0.00156858 3.3 0.00156868 0 0.0015685999999999999 0 0.0015687 3.3 0.00156862 3.3 0.00156872 0 0.0015686399999999998 0 0.0015687399999999999 3.3 0.00156866 3.3 0.00156876 0 0.0015686799999999998 0 0.0015687799999999999 3.3 0.0015687 3.3 0.0015688 0 0.00156872 0 0.00156882 3.3 0.0015687399999999999 3.3 0.00156884 0 0.00156876 0 0.00156886 3.3 0.0015687799999999999 3.3 0.00156888 0 0.0015688 0 0.0015689 3.3 0.0015688199999999999 3.3 0.00156892 0 0.00156884 0 0.00156894 3.3 0.0015688599999999998 3.3 0.0015689599999999999 0 0.00156888 0 0.00156898 3.3 0.0015688999999999998 3.3 0.0015689999999999999 0 0.00156892 0 0.00156902 3.3 0.00156894 3.3 0.00156904 0 0.0015689599999999999 0 0.00156906 3.3 0.00156898 3.3 0.00156908 0 0.0015689999999999999 0 0.0015691 3.3 0.00156902 3.3 0.00156912 0 0.0015690399999999998 0 0.00156914 3.3 0.00156906 3.3 0.00156916 0 0.0015690799999999998 0 0.0015691799999999999 3.3 0.0015691 3.3 0.0015692 0 0.00156912 0 0.00156922 3.3 0.00156914 3.3 0.00156924 0 0.00156916 0 0.00156926 3.3 0.0015691799999999999 3.3 0.00156928 0 0.0015692 0 0.0015693 3.3 0.0015692199999999999 3.3 0.00156932 0 0.00156924 0 0.00156934 3.3 0.0015692599999999998 3.3 0.00156936 0 0.00156928 0 0.00156938 3.3 0.0015692999999999998 3.3 0.0015693999999999999 0 0.00156932 0 0.00156942 3.3 0.00156934 3.3 0.00156944 0 0.00156936 0 0.00156946 3.3 0.00156938 3.3 0.00156948 0 0.0015693999999999999 0 0.0015695 3.3 0.00156942 3.3 0.00156952 0 0.0015694399999999999 0 0.00156954 3.3 0.00156946 3.3 0.00156956 0 0.0015694799999999998 0 0.0015695799999999999 3.3 0.0015695 3.3 0.0015696 0 0.0015695199999999998 0 0.0015696199999999999 3.3 0.00156954 3.3 0.00156964 0 0.00156956 0 0.00156966 3.3 0.0015695799999999999 3.3 0.00156968 0 0.0015696 0 0.0015697 3.3 0.0015696199999999999 3.3 0.00156972 0 0.00156964 0 0.00156974 3.3 0.0015696599999999998 3.3 0.00156976 0 0.00156968 0 0.00156978 3.3 0.0015696999999999998 3.3 0.0015697999999999999 0 0.00156972 0 0.00156982 3.3 0.0015697399999999998 3.3 0.0015698399999999999 0 0.00156976 0 0.00156986 3.3 0.00156978 3.3 0.00156988 0 0.0015697999999999999 0 0.0015699 3.3 0.00156982 3.3 0.00156992 0 0.0015698399999999999 0 0.00156994 3.3 0.00156986 3.3 0.00156996 0 0.0015698799999999998 0 0.00156998 3.3 0.0015699 3.3 0.00157 0 0.0015699199999999998 0 0.0015700199999999999 3.3 0.00156994 3.3 0.00157004 0 0.00156996 0 0.00157006 3.3 0.00156998 3.3 0.00157008 0 0.00157 0 0.0015701 3.3 0.0015700199999999999 3.3 0.00157012 0 0.00157004 0 0.00157014 3.3 0.0015700599999999999 3.3 0.00157016 0 0.00157008 0 0.00157018 3.3 0.0015700999999999998 3.3 0.0015702 0 0.00157012 0 0.00157022 3.3 0.0015701399999999998 3.3 0.0015702399999999999 0 0.00157016 0 0.00157026 3.3 0.00157018 3.3 0.00157028 0 0.0015702 0 0.0015703 3.3 0.00157022 3.3 0.00157032 0 0.0015702399999999999 0 0.00157034 3.3 0.00157026 3.3 0.00157036 0 0.0015702799999999999 0 0.00157038 3.3 0.0015703 3.3 0.0015704 0 0.0015703199999999998 0 0.0015704199999999999 3.3 0.00157034 3.3 0.00157044 0 0.0015703599999999998 0 0.0015704599999999999 3.3 0.00157038 3.3 0.00157048 0 0.0015704 0 0.0015705 3.3 0.0015704199999999999 3.3 0.00157052 0 0.00157044 0 0.00157054 3.3 0.0015704599999999999 3.3 0.00157056 0 0.00157048 0 0.00157058 3.3 0.0015704999999999998 3.3 0.0015706 0 0.00157052 0 0.00157062 3.3 0.0015705399999999998 3.3 0.0015706399999999999 0 0.00157056 0 0.00157066 3.3 0.0015705799999999998 3.3 0.0015706799999999999 0 0.0015706 0 0.0015707 3.3 0.00157062 3.3 0.00157072 0 0.0015706399999999999 0 0.00157074 3.3 0.00157066 3.3 0.00157076 0 0.0015706799999999999 0 0.00157078 3.3 0.0015707 3.3 0.0015708 0 0.0015707199999999998 0 0.00157082 3.3 0.00157074 3.3 0.00157084 0 0.0015707599999999998 0 0.0015708599999999999 3.3 0.00157078 3.3 0.00157088 0 0.0015708 0 0.0015709 3.3 0.00157082 3.3 0.00157092 0 0.00157084 0 0.00157094 3.3 0.0015708599999999999 3.3 0.00157096 0 0.00157088 0 0.00157098 3.3 0.0015708999999999999 3.3 0.001571 0 0.00157092 0 0.00157102 3.3 0.0015709399999999998 3.3 0.00157104 0 0.00157096 0 0.00157106 3.3 0.0015709799999999998 3.3 0.0015710799999999999 0 0.001571 0 0.0015711 3.3 0.00157102 3.3 0.00157112 0 0.00157104 0 0.00157114 3.3 0.00157106 3.3 0.00157116 0 0.0015710799999999999 0 0.00157118 3.3 0.0015711 3.3 0.0015712 0 0.0015711199999999999 0 0.00157122 3.3 0.00157114 3.3 0.00157124 0 0.0015711599999999998 0 0.0015712599999999999 3.3 0.00157118 3.3 0.00157128 0 0.0015711999999999998 0 0.0015712999999999999 3.3 0.00157122 3.3 0.00157132 0 0.00157124 0 0.00157134 3.3 0.0015712599999999999 3.3 0.00157136 0 0.00157128 0 0.00157138 3.3 0.0015712999999999999 3.3 0.0015714 0 0.00157132 0 0.00157142 3.3 0.0015713399999999998 3.3 0.00157144 0 0.00157136 0 0.00157146 3.3 0.0015713799999999998 3.3 0.0015714799999999999 0 0.0015714 0 0.0015715 3.3 0.0015714199999999998 3.3 0.0015715199999999999 0 0.00157144 0 0.00157154 3.3 0.00157146 3.3 0.00157156 0 0.0015714799999999999 0 0.00157158 3.3 0.0015715 3.3 0.0015716 0 0.0015715199999999999 0 0.00157162 3.3 0.00157154 3.3 0.00157164 0 0.0015715599999999998 0 0.00157166 3.3 0.00157158 3.3 0.00157168 0 0.0015715999999999998 0 0.0015716999999999999 3.3 0.00157162 3.3 0.00157172 0 0.00157164 0 0.00157174 3.3 0.00157166 3.3 0.00157176 0 0.00157168 0 0.00157178 3.3 0.0015716999999999999 3.3 0.0015718 0 0.00157172 0 0.00157182 3.3 0.0015717399999999999 3.3 0.00157184 0 0.00157176 0 0.00157186 3.3 0.0015717799999999998 3.3 0.00157188 0 0.0015718 0 0.0015719 3.3 0.0015718199999999998 3.3 0.0015719199999999999 0 0.00157184 0 0.00157194 3.3 0.00157186 3.3 0.00157196 0 0.00157188 0 0.00157198 3.3 0.0015719 3.3 0.001572 0 0.0015719199999999999 0 0.00157202 3.3 0.00157194 3.3 0.00157204 0 0.0015719599999999999 0 0.00157206 3.3 0.00157198 3.3 0.00157208 0 0.0015719999999999998 0 0.0015720999999999999 3.3 0.00157202 3.3 0.00157212 0 0.0015720399999999998 0 0.0015721399999999999 3.3 0.00157206 3.3 0.00157216 0 0.00157208 0 0.00157218 3.3 0.0015720999999999999 3.3 0.0015722 0 0.00157212 0 0.00157222 3.3 0.0015721399999999999 3.3 0.00157224 0 0.00157216 0 0.00157226 3.3 0.0015721799999999998 3.3 0.00157228 0 0.0015722 0 0.0015723 3.3 0.0015722199999999998 3.3 0.0015723199999999999 0 0.00157224 0 0.00157234 3.3 0.0015722599999999998 3.3 0.0015723599999999999 0 0.00157228 0 0.00157238 3.3 0.0015723 3.3 0.0015724 0 0.0015723199999999999 0 0.00157242 3.3 0.00157234 3.3 0.00157244 0 0.0015723599999999999 0 0.00157246 3.3 0.00157238 3.3 0.00157248 0 0.0015723999999999998 0 0.0015725 3.3 0.00157242 3.3 0.00157252 0 0.0015724399999999998 0 0.0015725399999999999 3.3 0.00157246 3.3 0.00157256 0 0.00157248 0 0.00157258 3.3 0.0015725 3.3 0.0015726 0 0.00157252 0 0.00157262 3.3 0.0015725399999999999 3.3 0.00157264 0 0.00157256 0 0.00157266 3.3 0.0015725799999999999 3.3 0.00157268 0 0.0015726 0 0.0015727 3.3 0.0015726199999999998 3.3 0.0015727199999999999 0 0.00157264 0 0.00157274 3.3 0.0015726599999999998 3.3 0.0015727599999999999 0 0.00157268 0 0.00157278 3.3 0.0015727 3.3 0.0015728 0 0.0015727199999999999 0 0.00157282 3.3 0.00157274 3.3 0.00157284 0 0.0015727599999999999 0 0.00157286 3.3 0.00157278 3.3 0.00157288 0 0.0015727999999999998 0 0.0015729 3.3 0.00157282 3.3 0.00157292 0 0.0015728399999999998 0 0.0015729399999999999 3.3 0.00157286 3.3 0.00157296 0 0.0015728799999999998 0 0.0015729799999999999 3.3 0.0015729 3.3 0.001573 0 0.00157292 0 0.00157302 3.3 0.0015729399999999999 3.3 0.00157304 0 0.00157296 0 0.00157306 3.3 0.0015729799999999999 3.3 0.00157308 0 0.001573 0 0.0015731 3.3 0.0015730199999999998 3.3 0.00157312 0 0.00157304 0 0.00157314 3.3 0.0015730599999999998 3.3 0.0015731599999999999 0 0.00157308 0 0.00157318 3.3 0.0015731 3.3 0.0015732 0 0.00157312 0 0.00157322 3.3 0.00157314 3.3 0.00157324 0 0.0015731599999999999 0 0.00157326 3.3 0.00157318 3.3 0.00157328 0 0.0015731999999999999 0 0.0015733 3.3 0.00157322 3.3 0.00157332 0 0.0015732399999999998 0 0.00157334 3.3 0.00157326 3.3 0.00157336 0 0.0015732799999999998 0 0.0015733799999999999 3.3 0.0015733 3.3 0.0015734 0 0.00157332 0 0.00157342 3.3 0.00157334 3.3 0.00157344 0 0.00157336 0 0.00157346 3.3 0.0015733799999999999 3.3 0.00157348 0 0.0015734 0 0.0015735 3.3 0.0015734199999999999 3.3 0.00157352 0 0.00157344 0 0.00157354 3.3 0.0015734599999999998 3.3 0.0015735599999999999 0 0.00157348 0 0.00157358 3.3 0.0015734999999999998 3.3 0.0015735999999999999 0 0.00157352 0 0.00157362 3.3 0.00157354 3.3 0.00157364 0 0.0015735599999999999 0 0.00157366 3.3 0.00157358 3.3 0.00157368 0 0.0015735999999999999 0 0.0015737 3.3 0.00157362 3.3 0.00157372 0 0.0015736399999999998 0 0.00157374 3.3 0.00157366 3.3 0.00157376 0 0.0015736799999999998 0 0.0015737799999999999 3.3 0.0015737 3.3 0.0015738 0 0.0015737199999999998 0 0.0015738199999999999 3.3 0.00157374 3.3 0.00157384 0 0.00157376 0 0.00157386 3.3 0.0015737799999999999 3.3 0.00157388 0 0.0015738 0 0.0015739 3.3 0.0015738199999999999 3.3 0.00157392 0 0.00157384 0 0.00157394 3.3 0.0015738599999999998 3.3 0.00157396 0 0.00157388 0 0.00157398 3.3 0.0015738999999999998 3.3 0.0015739999999999999 0 0.00157392 0 0.00157402 3.3 0.00157394 3.3 0.00157404 0 0.00157396 0 0.00157406 3.3 0.00157398 3.3 0.00157408 0 0.0015739999999999999 0 0.0015741 3.3 0.00157402 3.3 0.00157412 0 0.0015740399999999999 0 0.00157414 3.3 0.00157406 3.3 0.00157416 0 0.0015740799999999998 0 0.00157418 3.3 0.0015741 3.3 0.0015742 0 0.0015741199999999998 0 0.0015742199999999999 3.3 0.00157414 3.3 0.00157424 0 0.00157416 0 0.00157426 3.3 0.00157418 3.3 0.00157428 0 0.0015742 0 0.0015743 3.3 0.0015742199999999999 3.3 0.00157432 0 0.00157424 0 0.00157434 3.3 0.0015742599999999999 3.3 0.00157436 0 0.00157428 0 0.00157438 3.3 0.0015742999999999998 3.3 0.0015743999999999999 0 0.00157432 0 0.00157442 3.3 0.0015743399999999998 3.3 0.0015744399999999999 0 0.00157436 0 0.00157446 3.3 0.00157438 3.3 0.00157448 0 0.0015743999999999999 0 0.0015745 3.3 0.00157442 3.3 0.00157452 0 0.0015744399999999999 0 0.00157454 3.3 0.00157446 3.3 0.00157456 0 0.0015744799999999998 0 0.00157458 3.3 0.0015745 3.3 0.0015746 0 0.0015745199999999998 0 0.0015746199999999999 3.3 0.00157454 3.3 0.00157464 0 0.0015745599999999998 0 0.0015746599999999999 3.3 0.00157458 3.3 0.00157468 0 0.0015746 0 0.0015747 3.3 0.0015746199999999999 3.3 0.00157472 0 0.00157464 0 0.00157474 3.3 0.0015746599999999999 3.3 0.00157476 0 0.00157468 0 0.00157478 3.3 0.0015746999999999998 3.3 0.0015748 0 0.00157472 0 0.00157482 3.3 0.0015747399999999998 3.3 0.0015748399999999999 0 0.00157476 0 0.00157486 3.3 0.00157478 3.3 0.00157488 0 0.0015748 0 0.0015749 3.3 0.00157482 3.3 0.00157492 0 0.0015748399999999999 0 0.00157494 3.3 0.00157486 3.3 0.00157496 0 0.0015748799999999999 0 0.00157498 3.3 0.0015749 3.3 0.001575 0 0.0015749199999999998 0 0.00157502 3.3 0.00157494 3.3 0.00157504 0 0.0015749599999999998 0 0.0015750599999999999 3.3 0.00157498 3.3 0.00157508 0 0.001575 0 0.0015751 3.3 0.00157502 3.3 0.00157512 0 0.00157504 0 0.00157514 3.3 0.0015750599999999999 3.3 0.00157516 0 0.00157508 0 0.00157518 3.3 0.0015750999999999999 3.3 0.0015752 0 0.00157512 0 0.00157522 3.3 0.0015751399999999998 3.3 0.0015752399999999999 0 0.00157516 0 0.00157526 3.3 0.0015751799999999998 3.3 0.0015752799999999999 0 0.0015752 0 0.0015753 3.3 0.00157522 3.3 0.00157532 0 0.0015752399999999999 0 0.00157534 3.3 0.00157526 3.3 0.00157536 0 0.0015752799999999999 0 0.00157538 3.3 0.0015753 3.3 0.0015754 0 0.0015753199999999998 0 0.00157542 3.3 0.00157534 3.3 0.00157544 0 0.0015753599999999998 0 0.0015754599999999999 3.3 0.00157538 3.3 0.00157548 0 0.0015753999999999998 0 0.0015754999999999999 3.3 0.00157542 3.3 0.00157552 0 0.00157544 0 0.00157554 3.3 0.0015754599999999999 3.3 0.00157556 0 0.00157548 0 0.00157558 3.3 0.0015754999999999999 3.3 0.0015756 0 0.00157552 0 0.00157562 3.3 0.0015755399999999998 3.3 0.00157564 0 0.00157556 0 0.00157566 3.3 0.0015755799999999998 3.3 0.0015756799999999999 0 0.0015756 0 0.0015757 3.3 0.00157562 3.3 0.00157572 0 0.00157564 0 0.00157574 3.3 0.00157566 3.3 0.00157576 0 0.0015756799999999999 0 0.00157578 3.3 0.0015757 3.3 0.0015758 0 0.0015757199999999999 0 0.00157582 3.3 0.00157574 3.3 0.00157584 0 0.0015757599999999998 0 0.0015758599999999999 3.3 0.00157578 3.3 0.00157588 0 0.0015757999999999998 0 0.0015758999999999999 3.3 0.00157582 3.3 0.00157592 0 0.00157584 0 0.00157594 3.3 0.0015758599999999999 3.3 0.00157596 0 0.00157588 0 0.00157598 3.3 0.0015758999999999999 3.3 0.001576 0 0.00157592 0 0.00157602 3.3 0.0015759399999999998 3.3 0.00157604 0 0.00157596 0 0.00157606 3.3 0.0015759799999999998 3.3 0.0015760799999999999 0 0.001576 0 0.0015761 3.3 0.0015760199999999998 3.3 0.0015761199999999999 0 0.00157604 0 0.00157614 3.3 0.00157606 3.3 0.00157616 0 0.0015760799999999999 0 0.00157618 3.3 0.0015761 3.3 0.0015762 0 0.0015761199999999999 0 0.00157622 3.3 0.00157614 3.3 0.00157624 0 0.0015761599999999998 0 0.00157626 3.3 0.00157618 3.3 0.00157628 0 0.0015761999999999998 0 0.0015762999999999999 3.3 0.00157622 3.3 0.00157632 0 0.00157624 0 0.00157634 3.3 0.00157626 3.3 0.00157636 0 0.00157628 0 0.00157638 3.3 0.0015762999999999999 3.3 0.0015764 0 0.00157632 0 0.00157642 3.3 0.0015763399999999999 3.3 0.00157644 0 0.00157636 0 0.00157646 3.3 0.0015763799999999998 3.3 0.00157648 0 0.0015764 0 0.0015765 3.3 0.0015764199999999998 3.3 0.0015765199999999999 0 0.00157644 0 0.00157654 3.3 0.00157646 3.3 0.00157656 0 0.00157648 0 0.00157658 3.3 0.0015765 3.3 0.0015766 0 0.0015765199999999999 0 0.00157662 3.3 0.00157654 3.3 0.00157664 0 0.0015765599999999999 0 0.00157666 3.3 0.00157658 3.3 0.00157668 0 0.0015765999999999998 0 0.0015766999999999999 3.3 0.00157662 3.3 0.00157672 0 0.0015766399999999998 0 0.0015767399999999999 3.3 0.00157666 3.3 0.00157676 0 0.00157668 0 0.00157678 3.3 0.0015766999999999999 3.3 0.0015768 0 0.00157672 0 0.00157682 3.3 0.0015767399999999999 3.3 0.00157684 0 0.00157676 0 0.00157686 3.3 0.0015767799999999998 3.3 0.00157688 0 0.0015768 0 0.0015769 3.3 0.0015768199999999998 3.3 0.0015769199999999999 0 0.00157684 0 0.00157694 3.3 0.0015768599999999998 3.3 0.0015769599999999999 0 0.00157688 0 0.00157698 3.3 0.0015769 3.3 0.001577 0 0.0015769199999999999 0 0.00157702 3.3 0.00157694 3.3 0.00157704 0 0.0015769599999999999 0 0.00157706 3.3 0.00157698 3.3 0.00157708 0 0.0015769999999999998 0 0.0015771 3.3 0.00157702 3.3 0.00157712 0 0.0015770399999999998 0 0.0015771399999999999 3.3 0.00157706 3.3 0.00157716 0 0.00157708 0 0.00157718 3.3 0.0015771 3.3 0.0015772 0 0.00157712 0 0.00157722 3.3 0.0015771399999999999 3.3 0.00157724 0 0.00157716 0 0.00157726 3.3 0.0015771799999999999 3.3 0.00157728 0 0.0015772 0 0.0015773 3.3 0.0015772199999999998 3.3 0.00157732 0 0.00157724 0 0.00157734 3.3 0.0015772599999999998 3.3 0.0015773599999999999 0 0.00157728 0 0.00157738 3.3 0.0015773 3.3 0.0015774 0 0.00157732 0 0.00157742 3.3 0.00157734 3.3 0.00157744 0 0.0015773599999999999 0 0.00157746 3.3 0.00157738 3.3 0.00157748 0 0.0015773999999999999 0 0.0015775 3.3 0.00157742 3.3 0.00157752 0 0.0015774399999999998 0 0.0015775399999999999 3.3 0.00157746 3.3 0.00157756 0 0.0015774799999999998 0 0.0015775799999999999 3.3 0.0015775 3.3 0.0015776 0 0.00157752 0 0.00157762 3.3 0.0015775399999999999 3.3 0.00157764 0 0.00157756 0 0.00157766 3.3 0.0015775799999999999 3.3 0.00157768 0 0.0015776 0 0.0015777 3.3 0.0015776199999999998 3.3 0.00157772 0 0.00157764 0 0.00157774 3.3 0.0015776599999999998 3.3 0.0015777599999999999 0 0.00157768 0 0.00157778 3.3 0.0015776999999999998 3.3 0.0015777999999999999 0 0.00157772 0 0.00157782 3.3 0.00157774 3.3 0.00157784 0 0.0015777599999999999 0 0.00157786 3.3 0.00157778 3.3 0.00157788 0 0.0015777999999999999 0 0.0015779 3.3 0.00157782 3.3 0.00157792 0 0.0015778399999999998 0 0.00157794 3.3 0.00157786 3.3 0.00157796 0 0.0015778799999999998 0 0.0015779799999999999 3.3 0.0015779 3.3 0.001578 0 0.00157792 0 0.00157802 3.3 0.00157794 3.3 0.00157804 0 0.00157796 0 0.00157806 3.3 0.0015779799999999999 3.3 0.00157808 0 0.001578 0 0.0015781 3.3 0.0015780199999999999 3.3 0.00157812 0 0.00157804 0 0.00157814 3.3 0.0015780599999999998 3.3 0.00157816 0 0.00157808 0 0.00157818 3.3 0.0015780999999999998 3.3 0.0015781999999999999 0 0.00157812 0 0.00157822 3.3 0.00157814 3.3 0.00157824 0 0.00157816 0 0.00157826 3.3 0.00157818 3.3 0.00157828 0 0.0015781999999999999 0 0.0015783 3.3 0.00157822 3.3 0.00157832 0 0.0015782399999999999 0 0.00157834 3.3 0.00157826 3.3 0.00157836 0 0.0015782799999999998 0 0.0015783799999999999 3.3 0.0015783 3.3 0.0015784 0 0.0015783199999999998 0 0.0015784199999999999 3.3 0.00157834 3.3 0.00157844 0 0.00157836 0 0.00157846 3.3 0.0015783799999999999 3.3 0.00157848 0 0.0015784 0 0.0015785 3.3 0.0015784199999999999 3.3 0.00157852 0 0.00157844 0 0.00157854 3.3 0.0015784599999999998 3.3 0.00157856 0 0.00157848 0 0.00157858 3.3 0.0015784999999999998 3.3 0.0015785999999999999 0 0.00157852 0 0.00157862 3.3 0.0015785399999999998 3.3 0.0015786399999999999 0 0.00157856 0 0.00157866 3.3 0.00157858 3.3 0.00157868 0 0.0015785999999999999 0 0.0015787 3.3 0.00157862 3.3 0.00157872 0 0.0015786399999999999 0 0.00157874 3.3 0.00157866 3.3 0.00157876 0 0.0015786799999999998 0 0.00157878 3.3 0.0015787 3.3 0.0015788 0 0.0015787199999999998 0 0.0015788199999999999 3.3 0.00157874 3.3 0.00157884 0 0.00157876 0 0.00157886 3.3 0.00157878 3.3 0.00157888 0 0.0015788 0 0.0015789 3.3 0.0015788199999999999 3.3 0.00157892 0 0.00157884 0 0.00157894 3.3 0.0015788599999999999 3.3 0.00157896 0 0.00157888 0 0.00157898 3.3 0.0015788999999999998 3.3 0.0015789999999999999 0 0.00157892 0 0.00157902 3.3 0.0015789399999999998 3.3 0.0015790399999999999 0 0.00157896 0 0.00157906 3.3 0.00157898 3.3 0.00157908 0 0.0015789999999999999 0 0.0015791 3.3 0.00157902 3.3 0.00157912 0 0.0015790399999999999 0 0.00157914 3.3 0.00157906 3.3 0.00157916 0 0.0015790799999999999 0 0.00157918 3.3 0.0015791 3.3 0.0015792 0 0.0015791199999999998 0 0.0015792199999999999 3.3 0.00157914 3.3 0.00157924 0 0.0015791599999999998 0 0.0015792599999999999 3.3 0.00157918 3.3 0.00157928 0 0.0015792 0 0.0015793 3.3 0.0015792199999999999 3.3 0.00157932 0 0.00157924 0 0.00157934 3.3 0.0015792599999999999 3.3 0.00157936 0 0.00157928 0 0.00157938 3.3 0.0015792999999999998 3.3 0.0015794 0 0.00157932 0 0.00157942 3.3 0.0015793399999999998 3.3 0.0015794399999999999 0 0.00157936 0 0.00157946 3.3 0.00157938 3.3 0.00157948 0 0.0015794 0 0.0015795 3.3 0.00157942 3.3 0.00157952 0 0.0015794399999999999 0 0.00157954 3.3 0.00157946 3.3 0.00157956 0 0.0015794799999999999 0 0.00157958 3.3 0.0015795 3.3 0.0015796 0 0.0015795199999999998 0 0.00157962 3.3 0.00157954 3.3 0.00157964 0 0.0015795599999999998 0 0.0015796599999999999 3.3 0.00157958 3.3 0.00157968 0 0.0015796 0 0.0015797 3.3 0.00157962 3.3 0.00157972 0 0.00157964 0 0.00157974 3.3 0.0015796599999999999 3.3 0.00157976 0 0.00157968 0 0.00157978 3.3 0.0015796999999999999 3.3 0.0015798 0 0.00157972 0 0.00157982 3.3 0.0015797399999999998 3.3 0.0015798399999999999 0 0.00157976 0 0.00157986 3.3 0.0015797799999999998 3.3 0.0015798799999999999 0 0.0015798 0 0.0015799 3.3 0.00157982 3.3 0.00157992 0 0.0015798399999999999 0 0.00157994 3.3 0.00157986 3.3 0.00157996 0 0.0015798799999999999 0 0.00157998 3.3 0.0015799 3.3 0.00158 0 0.0015799199999999998 0 0.00158002 3.3 0.00157994 3.3 0.00158004 0 0.0015799599999999998 0 0.0015800599999999999 3.3 0.00157998 3.3 0.00158008 0 0.0015799999999999998 0 0.0015800999999999999 3.3 0.00158002 3.3 0.00158012 0 0.00158004 0 0.00158014 3.3 0.0015800599999999999 3.3 0.00158016 0 0.00158008 0 0.00158018 3.3 0.0015800999999999999 3.3 0.0015802 0 0.00158012 0 0.00158022 3.3 0.0015801399999999998 3.3 0.00158024 0 0.00158016 0 0.00158026 3.3 0.0015801799999999998 3.3 0.0015802799999999999 0 0.0015802 0 0.0015803 3.3 0.00158022 3.3 0.00158032 0 0.00158024 0 0.00158034 3.3 0.00158026 3.3 0.00158036 0 0.0015802799999999999 0 0.00158038 3.3 0.0015803 3.3 0.0015804 0 0.0015803199999999999 0 0.00158042 3.3 0.00158034 3.3 0.00158044 0 0.0015803599999999998 0 0.00158046 3.3 0.00158038 3.3 0.00158048 0 0.0015803999999999998 0 0.0015804999999999999 3.3 0.00158042 3.3 0.00158052 0 0.00158044 0 0.00158054 3.3 0.00158046 3.3 0.00158056 0 0.00158048 0 0.00158058 3.3 0.0015804999999999999 3.3 0.0015806 0 0.00158052 0 0.00158062 3.3 0.0015805399999999999 3.3 0.00158064 0 0.00158056 0 0.00158066 3.3 0.0015805799999999998 3.3 0.0015806799999999999 0 0.0015806 0 0.0015807 3.3 0.0015806199999999998 3.3 0.0015807199999999999 0 0.00158064 0 0.00158074 3.3 0.00158066 3.3 0.00158076 0 0.0015806799999999999 0 0.00158078 3.3 0.0015807 3.3 0.0015808 0 0.0015807199999999999 0 0.00158082 3.3 0.00158074 3.3 0.00158084 0 0.0015807599999999998 0 0.00158086 3.3 0.00158078 3.3 0.00158088 0 0.0015807999999999998 0 0.0015808999999999999 3.3 0.00158082 3.3 0.00158092 0 0.0015808399999999998 0 0.0015809399999999999 3.3 0.00158086 3.3 0.00158096 0 0.00158088 0 0.00158098 3.3 0.0015808999999999999 3.3 0.001581 0 0.00158092 0 0.00158102 3.3 0.0015809399999999999 3.3 0.00158104 0 0.00158096 0 0.00158106 3.3 0.0015809799999999998 3.3 0.00158108 0 0.001581 0 0.0015811 3.3 0.0015810199999999998 3.3 0.0015811199999999999 0 0.00158104 0 0.00158114 3.3 0.00158106 3.3 0.00158116 0 0.00158108 0 0.00158118 3.3 0.0015811 3.3 0.0015812 0 0.0015811199999999999 0 0.00158122 3.3 0.00158114 3.3 0.00158124 0 0.0015811599999999999 0 0.00158126 3.3 0.00158118 3.3 0.00158128 0 0.0015811999999999998 0 0.0015813 3.3 0.00158122 3.3 0.00158132 0 0.0015812399999999998 0 0.0015813399999999999 3.3 0.00158126 3.3 0.00158136 0 0.00158128 0 0.00158138 3.3 0.0015813 3.3 0.0015814 0 0.00158132 0 0.00158142 3.3 0.0015813399999999999 3.3 0.00158144 0 0.00158136 0 0.00158146 3.3 0.0015813799999999999 3.3 0.00158148 0 0.0015814 0 0.0015815 3.3 0.0015814199999999998 3.3 0.0015815199999999999 0 0.00158144 0 0.00158154 3.3 0.0015814599999999998 3.3 0.0015815599999999999 0 0.00158148 0 0.00158158 3.3 0.0015815 3.3 0.0015816 0 0.0015815199999999999 0 0.00158162 3.3 0.00158154 3.3 0.00158164 0 0.0015815599999999999 0 0.00158166 3.3 0.00158158 3.3 0.00158168 0 0.0015815999999999998 0 0.0015817 3.3 0.00158162 3.3 0.00158172 0 0.0015816399999999998 0 0.0015817399999999999 3.3 0.00158166 3.3 0.00158176 0 0.0015816799999999998 0 0.0015817799999999999 3.3 0.0015817 3.3 0.0015818 0 0.00158172 0 0.00158182 3.3 0.0015817399999999999 3.3 0.00158184 0 0.00158176 0 0.00158186 3.3 0.0015817799999999999 3.3 0.00158188 0 0.0015818 0 0.0015819 3.3 0.0015818199999999998 3.3 0.00158192 0 0.00158184 0 0.00158194 3.3 0.0015818599999999998 3.3 0.0015819599999999999 0 0.00158188 0 0.00158198 3.3 0.0015819 3.3 0.001582 0 0.00158192 0 0.00158202 3.3 0.00158194 3.3 0.00158204 0 0.0015819599999999999 0 0.00158206 3.3 0.00158198 3.3 0.00158208 0 0.0015819999999999999 0 0.0015821 3.3 0.00158202 3.3 0.00158212 0 0.0015820399999999998 0 0.00158214 3.3 0.00158206 3.3 0.00158216 0 0.0015820799999999998 0 0.0015821799999999999 3.3 0.0015821 3.3 0.0015822 0 0.00158212 0 0.00158222 3.3 0.00158214 3.3 0.00158224 0 0.00158216 0 0.00158226 3.3 0.0015821799999999999 3.3 0.00158228 0 0.0015822 0 0.0015823 3.3 0.0015822199999999999 3.3 0.00158232 0 0.00158224 0 0.00158234 3.3 0.0015822599999999998 3.3 0.0015823599999999999 0 0.00158228 0 0.00158238 3.3 0.0015822999999999998 3.3 0.0015823999999999999 0 0.00158232 0 0.00158242 3.3 0.00158234 3.3 0.00158244 0 0.0015823599999999999 0 0.00158246 3.3 0.00158238 3.3 0.00158248 0 0.0015823999999999999 0 0.0015825 3.3 0.00158242 3.3 0.00158252 0 0.0015824399999999998 0 0.00158254 3.3 0.00158246 3.3 0.00158256 0 0.0015824799999999998 0 0.0015825799999999999 3.3 0.0015825 3.3 0.0015826 0 0.0015825199999999998 0 0.0015826199999999999 3.3 0.00158254 3.3 0.00158264 0 0.00158256 0 0.00158266 3.3 0.0015825799999999999 3.3 0.00158268 0 0.0015826 0 0.0015827 3.3 0.0015826199999999999 3.3 0.00158272 0 0.00158264 0 0.00158274 3.3 0.0015826599999999998 3.3 0.00158276 0 0.00158268 0 0.00158278 3.3 0.0015826999999999998 3.3 0.0015827999999999999 0 0.00158272 0 0.00158282 3.3 0.00158274 3.3 0.00158284 0 0.00158276 0 0.00158286 3.3 0.00158278 3.3 0.00158288 0 0.0015827999999999999 0 0.0015829 3.3 0.00158282 3.3 0.00158292 0 0.0015828399999999999 0 0.00158294 3.3 0.00158286 3.3 0.00158296 0 0.0015828799999999998 0 0.0015829799999999999 3.3 0.0015829 3.3 0.001583 0 0.0015829199999999998 0 0.0015830199999999999 3.3 0.00158294 3.3 0.00158304 0 0.00158296 0 0.00158306 3.3 0.0015829799999999999 3.3 0.00158308 0 0.001583 0 0.0015831 3.3 0.0015830199999999999 3.3 0.00158312 0 0.00158304 0 0.00158314 3.3 0.0015830599999999998 3.3 0.00158316 0 0.00158308 0 0.00158318 3.3 0.0015830999999999998 3.3 0.0015831999999999999 0 0.00158312 0 0.00158322 3.3 0.0015831399999999998 3.3 0.0015832399999999999 0 0.00158316 0 0.00158326 3.3 0.00158318 3.3 0.00158328 0 0.0015831999999999999 0 0.0015833 3.3 0.00158322 3.3 0.00158332 0 0.0015832399999999999 0 0.00158334 3.3 0.00158326 3.3 0.00158336 0 0.0015832799999999998 0 0.00158338 3.3 0.0015833 3.3 0.0015834 0 0.0015833199999999998 0 0.0015834199999999999 3.3 0.00158334 3.3 0.00158344 0 0.00158336 0 0.00158346 3.3 0.00158338 3.3 0.00158348 0 0.0015834 0 0.0015835 3.3 0.0015834199999999999 3.3 0.00158352 0 0.00158344 0 0.00158354 3.3 0.0015834599999999999 3.3 0.00158356 0 0.00158348 0 0.00158358 3.3 0.0015834999999999998 3.3 0.0015836 0 0.00158352 0 0.00158362 3.3 0.0015835399999999998 3.3 0.0015836399999999999 0 0.00158356 0 0.00158366 3.3 0.00158358 3.3 0.00158368 0 0.0015836 0 0.0015837 3.3 0.00158362 3.3 0.00158372 0 0.0015836399999999999 0 0.00158374 3.3 0.00158366 3.3 0.00158376 0 0.0015836799999999999 0 0.00158378 3.3 0.0015837 3.3 0.0015838 0 0.0015837199999999998 0 0.0015838199999999999 3.3 0.00158374 3.3 0.00158384 0 0.0015837599999999998 0 0.0015838599999999999 3.3 0.00158378 3.3 0.00158388 0 0.0015838 0 0.0015839 3.3 0.0015838199999999999 3.3 0.00158392 0 0.00158384 0 0.00158394 3.3 0.0015838599999999999 3.3 0.00158396 0 0.00158388 0 0.00158398 3.3 0.0015838999999999998 3.3 0.001584 0 0.00158392 0 0.00158402 3.3 0.0015839399999999998 3.3 0.0015840399999999999 0 0.00158396 0 0.00158406 3.3 0.0015839799999999998 3.3 0.0015840799999999999 0 0.001584 0 0.0015841 3.3 0.00158402 3.3 0.00158412 0 0.0015840399999999999 0 0.00158414 3.3 0.00158406 3.3 0.00158416 0 0.0015840799999999999 0 0.00158418 3.3 0.0015841 3.3 0.0015842 0 0.0015841199999999998 0 0.00158422 3.3 0.00158414 3.3 0.00158424 0 0.0015841599999999998 0 0.0015842599999999999 3.3 0.00158418 3.3 0.00158428 0 0.0015842 0 0.0015843 3.3 0.00158422 3.3 0.00158432 0 0.00158424 0 0.00158434 3.3 0.0015842599999999999 3.3 0.00158436 0 0.00158428 0 0.00158438 3.3 0.0015842999999999999 3.3 0.0015844 0 0.00158432 0 0.00158442 3.3 0.0015843399999999998 3.3 0.00158444 0 0.00158436 0 0.00158446 3.3 0.0015843799999999998 3.3 0.0015844799999999999 0 0.0015844 0 0.0015845 3.3 0.00158442 3.3 0.00158452 0 0.00158444 0 0.00158454 3.3 0.00158446 3.3 0.00158456 0 0.0015844799999999999 0 0.00158458 3.3 0.0015845 3.3 0.0015846 0 0.0015845199999999999 0 0.00158462 3.3 0.00158454 3.3 0.00158464 0 0.0015845599999999998 0 0.0015846599999999999 3.3 0.00158458 3.3 0.00158468 0 0.0015845999999999998 0 0.0015846999999999999 3.3 0.00158462 3.3 0.00158472 0 0.00158464 0 0.00158474 3.3 0.0015846599999999999 3.3 0.00158476 0 0.00158468 0 0.00158478 3.3 0.0015846999999999999 3.3 0.0015848 0 0.00158472 0 0.00158482 3.3 0.0015847399999999998 3.3 0.00158484 0 0.00158476 0 0.00158486 3.3 0.0015847799999999998 3.3 0.0015848799999999999 0 0.0015848 0 0.0015849 3.3 0.0015848199999999998 3.3 0.0015849199999999999 0 0.00158484 0 0.00158494 3.3 0.00158486 3.3 0.00158496 0 0.0015848799999999999 0 0.00158498 3.3 0.0015849 3.3 0.001585 0 0.0015849199999999999 0 0.00158502 3.3 0.00158494 3.3 0.00158504 0 0.0015849599999999998 0 0.00158506 3.3 0.00158498 3.3 0.00158508 0 0.0015849999999999998 0 0.0015850999999999999 3.3 0.00158502 3.3 0.00158512 0 0.00158504 0 0.00158514 3.3 0.00158506 3.3 0.00158516 0 0.00158508 0 0.00158518 3.3 0.0015850999999999999 3.3 0.0015852 0 0.00158512 0 0.00158522 3.3 0.0015851399999999999 3.3 0.00158524 0 0.00158516 0 0.00158526 3.3 0.0015851799999999998 3.3 0.00158528 0 0.0015852 0 0.0015853 3.3 0.0015852199999999998 3.3 0.0015853199999999999 0 0.00158524 0 0.00158534 3.3 0.00158526 3.3 0.00158536 0 0.00158528 0 0.00158538 3.3 0.0015853 3.3 0.0015854 0 0.0015853199999999999 0 0.00158542 3.3 0.00158534 3.3 0.00158544 0 0.0015853599999999999 0 0.00158546 3.3 0.00158538 3.3 0.00158548 0 0.0015853999999999998 0 0.0015854999999999999 3.3 0.00158542 3.3 0.00158552 0 0.0015854399999999998 0 0.0015855399999999999 3.3 0.00158546 3.3 0.00158556 0 0.00158548 0 0.00158558 3.3 0.0015854999999999999 3.3 0.0015856 0 0.00158552 0 0.00158562 3.3 0.0015855399999999999 3.3 0.00158564 0 0.00158556 0 0.00158566 3.3 0.0015855799999999998 3.3 0.00158568 0 0.0015856 0 0.0015857 3.3 0.0015856199999999998 3.3 0.0015857199999999999 0 0.00158564 0 0.00158574 3.3 0.0015856599999999998 3.3 0.0015857599999999999 0 0.00158568 0 0.00158578 3.3 0.0015857 3.3 0.0015858 0 0.0015857199999999999 0 0.00158582 3.3 0.00158574 3.3 0.00158584 0 0.0015857599999999999 0 0.00158586 3.3 0.00158578 3.3 0.00158588 0 0.0015857999999999998 0 0.0015859 3.3 0.00158582 3.3 0.00158592 0 0.0015858399999999998 0 0.0015859399999999999 3.3 0.00158586 3.3 0.00158596 0 0.00158588 0 0.00158598 3.3 0.0015859 3.3 0.001586 0 0.00158592 0 0.00158602 3.3 0.0015859399999999999 3.3 0.00158604 0 0.00158596 0 0.00158606 3.3 0.0015859799999999999 3.3 0.00158608 0 0.001586 0 0.0015861 3.3 0.0015860199999999998 3.3 0.0015861199999999999 0 0.00158604 0 0.00158614 3.3 0.0015860599999999998 3.3 0.0015861599999999999 0 0.00158608 0 0.00158618 3.3 0.0015861 3.3 0.0015862 0 0.0015861199999999999 0 0.00158622 3.3 0.00158614 3.3 0.00158624 0 0.0015861599999999999 0 0.00158626 3.3 0.00158618 3.3 0.00158628 0 0.0015861999999999998 0 0.0015863 3.3 0.00158622 3.3 0.00158632 0 0.0015862399999999998 0 0.0015863399999999999 3.3 0.00158626 3.3 0.00158636 0 0.0015862799999999998 0 0.0015863799999999999 3.3 0.0015863 3.3 0.0015864 0 0.00158632 0 0.00158642 3.3 0.0015863399999999999 3.3 0.00158644 0 0.00158636 0 0.00158646 3.3 0.0015863799999999999 3.3 0.00158648 0 0.0015864 0 0.0015865 3.3 0.0015864199999999998 3.3 0.00158652 0 0.00158644 0 0.00158654 3.3 0.0015864599999999998 3.3 0.0015865599999999999 0 0.00158648 0 0.00158658 3.3 0.0015865 3.3 0.0015866 0 0.00158652 0 0.00158662 3.3 0.00158654 3.3 0.00158664 0 0.0015865599999999999 0 0.00158666 3.3 0.00158658 3.3 0.00158668 0 0.0015865999999999999 0 0.0015867 3.3 0.00158662 3.3 0.00158672 0 0.0015866399999999998 0 0.00158674 3.3 0.00158666 3.3 0.00158676 0 0.0015866799999999998 0 0.0015867799999999999 3.3 0.0015867 3.3 0.0015868 0 0.00158672 0 0.00158682 3.3 0.00158674 3.3 0.00158684 0 0.00158676 0 0.00158686 3.3 0.0015867799999999999 3.3 0.00158688 0 0.0015868 0 0.0015869 3.3 0.0015868199999999999 3.3 0.00158692 0 0.00158684 0 0.00158694 3.3 0.0015868599999999998 3.3 0.0015869599999999999 0 0.00158688 0 0.00158698 3.3 0.0015868999999999998 3.3 0.0015869999999999999 0 0.00158692 0 0.00158702 3.3 0.00158694 3.3 0.00158704 0 0.0015869599999999999 0 0.00158706 3.3 0.00158698 3.3 0.00158708 0 0.0015869999999999999 0 0.0015871 3.3 0.00158702 3.3 0.00158712 0 0.0015870399999999998 0 0.00158714 3.3 0.00158706 3.3 0.00158716 0 0.0015870799999999998 0 0.0015871799999999999 3.3 0.0015871 3.3 0.0015872 0 0.0015871199999999998 0 0.0015872199999999999 3.3 0.00158714 3.3 0.00158724 0 0.00158716 0 0.00158726 3.3 0.0015871799999999999 3.3 0.00158728 0 0.0015872 0 0.0015873 3.3 0.0015872199999999999 3.3 0.00158732 0 0.00158724 0 0.00158734 3.3 0.0015872599999999998 3.3 0.00158736 0 0.00158728 0 0.00158738 3.3 0.0015872999999999998 3.3 0.0015873999999999999 0 0.00158732 0 0.00158742 3.3 0.00158734 3.3 0.00158744 0 0.00158736 0 0.00158746 3.3 0.00158738 3.3 0.00158748 0 0.0015873999999999999 0 0.0015875 3.3 0.00158742 3.3 0.00158752 0 0.0015874399999999999 0 0.00158754 3.3 0.00158746 3.3 0.00158756 0 0.0015874799999999998 0 0.00158758 3.3 0.0015875 3.3 0.0015876 0 0.0015875199999999998 0 0.0015876199999999999 3.3 0.00158754 3.3 0.00158764 0 0.00158756 0 0.00158766 3.3 0.00158758 3.3 0.00158768 0 0.0015876 0 0.0015877 3.3 0.0015876199999999999 3.3 0.00158772 0 0.00158764 0 0.00158774 3.3 0.0015876599999999999 3.3 0.00158776 0 0.00158768 0 0.00158778 3.3 0.0015876999999999998 3.3 0.0015877999999999999 0 0.00158772 0 0.00158782 3.3 0.0015877399999999998 3.3 0.0015878399999999999 0 0.00158776 0 0.00158786 3.3 0.00158778 3.3 0.00158788 0 0.0015877999999999999 0 0.0015879 3.3 0.00158782 3.3 0.00158792 0 0.0015878399999999999 0 0.00158794 3.3 0.00158786 3.3 0.00158796 0 0.0015878799999999998 0 0.00158798 3.3 0.0015879 3.3 0.001588 0 0.0015879199999999998 0 0.0015880199999999999 3.3 0.00158794 3.3 0.00158804 0 0.0015879599999999998 0 0.0015880599999999999 3.3 0.00158798 3.3 0.00158808 0 0.001588 0 0.0015881 3.3 0.0015880199999999999 3.3 0.00158812 0 0.00158804 0 0.00158814 3.3 0.0015880599999999999 3.3 0.00158816 0 0.00158808 0 0.00158818 3.3 0.0015880999999999998 3.3 0.0015882 0 0.00158812 0 0.00158822 3.3 0.0015881399999999998 3.3 0.0015882399999999999 0 0.00158816 0 0.00158826 3.3 0.00158818 3.3 0.00158828 0 0.0015882 0 0.0015883 3.3 0.00158822 3.3 0.00158832 0 0.0015882399999999999 0 0.00158834 3.3 0.00158826 3.3 0.00158836 0 0.0015882799999999999 0 0.00158838 3.3 0.0015883 3.3 0.0015884 0 0.0015883199999999998 0 0.00158842 3.3 0.00158834 3.3 0.00158844 0 0.0015883599999999998 0 0.0015884599999999999 3.3 0.00158838 3.3 0.00158848 0 0.0015884 0 0.0015885 3.3 0.00158842 3.3 0.00158852 0 0.00158844 0 0.00158854 3.3 0.0015884599999999999 3.3 0.00158856 0 0.00158848 0 0.00158858 3.3 0.0015884999999999999 3.3 0.0015886 0 0.00158852 0 0.00158862 3.3 0.0015885399999999998 3.3 0.0015886399999999999 0 0.00158856 0 0.00158866 3.3 0.0015885799999999998 3.3 0.0015886799999999999 0 0.0015886 0 0.0015887 3.3 0.00158862 3.3 0.00158872 0 0.0015886399999999999 0 0.00158874 3.3 0.00158866 3.3 0.00158876 0 0.0015886799999999999 0 0.00158878 3.3 0.0015887 3.3 0.0015888 0 0.0015887199999999998 0 0.00158882 3.3 0.00158874 3.3 0.00158884 0 0.0015887599999999998 0 0.0015888599999999999 3.3 0.00158878 3.3 0.00158888 0 0.0015887999999999998 0 0.0015888999999999999 3.3 0.00158882 3.3 0.00158892 0 0.00158884 0 0.00158894 3.3 0.0015888599999999999 3.3 0.00158896 0 0.00158888 0 0.00158898 3.3 0.0015888999999999999 3.3 0.001589 0 0.00158892 0 0.00158902 3.3 0.0015889399999999998 3.3 0.00158904 0 0.00158896 0 0.00158906 3.3 0.0015889799999999998 3.3 0.0015890799999999999 0 0.001589 0 0.0015891 3.3 0.00158902 3.3 0.00158912 0 0.00158904 0 0.00158914 3.3 0.00158906 3.3 0.00158916 0 0.0015890799999999999 0 0.00158918 3.3 0.0015891 3.3 0.0015892 0 0.0015891199999999999 0 0.00158922 3.3 0.00158914 3.3 0.00158924 0 0.0015891599999999998 0 0.0015892599999999999 3.3 0.00158918 3.3 0.00158928 0 0.0015891999999999998 0 0.0015892999999999999 3.3 0.00158922 3.3 0.00158932 0 0.00158924 0 0.00158934 3.3 0.0015892599999999999 3.3 0.00158936 0 0.00158928 0 0.00158938 3.3 0.0015892999999999999 3.3 0.0015894 0 0.00158932 0 0.00158942 3.3 0.0015893399999999999 3.3 0.00158944 0 0.00158936 0 0.00158946 3.3 0.0015893799999999998 3.3 0.0015894799999999999 0 0.0015894 0 0.0015895 3.3 0.0015894199999999998 3.3 0.0015895199999999999 0 0.00158944 0 0.00158954 3.3 0.00158946 3.3 0.00158956 0 0.0015894799999999999 0 0.00158958 3.3 0.0015895 3.3 0.0015896 0 0.0015895199999999999 0 0.00158962 3.3 0.00158954 3.3 0.00158964 0 0.0015895599999999998 0 0.00158966 3.3 0.00158958 3.3 0.00158968 0 0.0015895999999999998 0 0.0015896999999999999 3.3 0.00158962 3.3 0.00158972 0 0.0015896399999999998 0 0.0015897399999999999 3.3 0.00158966 3.3 0.00158976 0 0.00158968 0 0.00158978 3.3 0.0015896999999999999 3.3 0.0015898 0 0.00158972 0 0.00158982 3.3 0.0015897399999999999 3.3 0.00158984 0 0.00158976 0 0.00158986 3.3 0.0015897799999999998 3.3 0.00158988 0 0.0015898 0 0.0015899 3.3 0.0015898199999999998 3.3 0.0015899199999999999 0 0.00158984 0 0.00158994 3.3 0.00158986 3.3 0.00158996 0 0.00158988 0 0.00158998 3.3 0.0015899 3.3 0.00159 0 0.0015899199999999999 0 0.00159002 3.3 0.00158994 3.3 0.00159004 0 0.0015899599999999999 0 0.00159006 3.3 0.00158998 3.3 0.00159008 0 0.0015899999999999998 0 0.0015900999999999999 3.3 0.00159002 3.3 0.00159012 0 0.0015900399999999998 0 0.0015901399999999999 3.3 0.00159006 3.3 0.00159016 0 0.00159008 0 0.00159018 3.3 0.0015900999999999999 3.3 0.0015902 0 0.00159012 0 0.00159022 3.3 0.0015901399999999999 3.3 0.00159024 0 0.00159016 0 0.00159026 3.3 0.0015901799999999998 3.3 0.00159028 0 0.0015902 0 0.0015903 3.3 0.0015902199999999998 3.3 0.0015903199999999999 0 0.00159024 0 0.00159034 3.3 0.0015902599999999998 3.3 0.0015903599999999999 0 0.00159028 0 0.00159038 3.3 0.0015903 3.3 0.0015904 0 0.0015903199999999999 0 0.00159042 3.3 0.00159034 3.3 0.00159044 0 0.0015903599999999999 0 0.00159046 3.3 0.00159038 3.3 0.00159048 0 0.0015903999999999998 0 0.0015905 3.3 0.00159042 3.3 0.00159052 0 0.0015904399999999998 0 0.0015905399999999999 3.3 0.00159046 3.3 0.00159056 0 0.00159048 0 0.00159058 3.3 0.0015905 3.3 0.0015906 0 0.00159052 0 0.00159062 3.3 0.0015905399999999999 3.3 0.00159064 0 0.00159056 0 0.00159066 3.3 0.0015905799999999999 3.3 0.00159068 0 0.0015906 0 0.0015907 3.3 0.0015906199999999998 3.3 0.00159072 0 0.00159064 0 0.00159074 3.3 0.0015906599999999998 3.3 0.0015907599999999999 0 0.00159068 0 0.00159078 3.3 0.0015907 3.3 0.0015908 0 0.00159072 0 0.00159082 3.3 0.00159074 3.3 0.00159084 0 0.0015907599999999999 0 0.00159086 3.3 0.00159078 3.3 0.00159088 0 0.0015907999999999999 0 0.0015909 3.3 0.00159082 3.3 0.00159092 0 0.0015908399999999998 0 0.0015909399999999999 3.3 0.00159086 3.3 0.00159096 0 0.0015908799999999998 0 0.0015909799999999999 3.3 0.0015909 3.3 0.001591 0 0.00159092 0 0.00159102 3.3 0.0015909399999999999 3.3 0.00159104 0 0.00159096 0 0.00159106 3.3 0.0015909799999999999 3.3 0.00159108 0 0.001591 0 0.0015911 3.3 0.0015910199999999998 3.3 0.00159112 0 0.00159104 0 0.00159114 3.3 0.0015910599999999998 3.3 0.0015911599999999999 0 0.00159108 0 0.00159118 3.3 0.0015910999999999998 3.3 0.0015911999999999999 0 0.00159112 0 0.00159122 3.3 0.00159114 3.3 0.00159124 0 0.0015911599999999999 0 0.00159126 3.3 0.00159118 3.3 0.00159128 0 0.0015911999999999999 0 0.0015913 3.3 0.00159122 3.3 0.00159132 0 0.0015912399999999998 0 0.00159134 3.3 0.00159126 3.3 0.00159136 0 0.0015912799999999998 0 0.0015913799999999999 3.3 0.0015913 3.3 0.0015914 0 0.00159132 0 0.00159142 3.3 0.00159134 3.3 0.00159144 0 0.00159136 0 0.00159146 3.3 0.0015913799999999999 3.3 0.00159148 0 0.0015914 0 0.0015915 3.3 0.0015914199999999999 3.3 0.00159152 0 0.00159144 0 0.00159154 3.3 0.0015914599999999998 3.3 0.00159156 0 0.00159148 0 0.00159158 3.3 0.0015914999999999998 3.3 0.0015915999999999999 0 0.00159152 0 0.00159162 3.3 0.00159154 3.3 0.00159164 0 0.00159156 0 0.00159166 3.3 0.00159158 3.3 0.00159168 0 0.0015915999999999999 0 0.0015917 3.3 0.00159162 3.3 0.00159172 0 0.0015916399999999999 0 0.00159174 3.3 0.00159166 3.3 0.00159176 0 0.0015916799999999998 0 0.0015917799999999999 3.3 0.0015917 3.3 0.0015918 0 0.0015917199999999998 0 0.0015918199999999999 3.3 0.00159174 3.3 0.00159184 0 0.00159176 0 0.00159186 3.3 0.0015917799999999999 3.3 0.00159188 0 0.0015918 0 0.0015919 3.3 0.0015918199999999999 3.3 0.00159192 0 0.00159184 0 0.00159194 3.3 0.0015918599999999998 3.3 0.00159196 0 0.00159188 0 0.00159198 3.3 0.0015918999999999998 3.3 0.0015919999999999999 0 0.00159192 0 0.00159202 3.3 0.0015919399999999998 3.3 0.0015920399999999999 0 0.00159196 0 0.00159206 3.3 0.00159198 3.3 0.00159208 0 0.0015919999999999999 0 0.0015921 3.3 0.00159202 3.3 0.00159212 0 0.0015920399999999999 0 0.00159214 3.3 0.00159206 3.3 0.00159216 0 0.0015920799999999998 0 0.00159218 3.3 0.0015921 3.3 0.0015922 0 0.0015921199999999998 0 0.0015922199999999999 3.3 0.00159214 3.3 0.00159224 0 0.00159216 0 0.00159226 3.3 0.00159218 3.3 0.00159228 0 0.0015922 0 0.0015923 3.3 0.0015922199999999999 3.3 0.00159232 0 0.00159224 0 0.00159234 3.3 0.0015922599999999999 3.3 0.00159236 0 0.00159228 0 0.00159238 3.3 0.0015922999999999998 3.3 0.0015924 0 0.00159232 0 0.00159242 3.3 0.0015923399999999998 3.3 0.0015924399999999999 0 0.00159236 0 0.00159246 3.3 0.00159238 3.3 0.00159248 0 0.0015924 0 0.0015925 3.3 0.00159242 3.3 0.00159252 0 0.0015924399999999999 0 0.00159254 3.3 0.00159246 3.3 0.00159256 0 0.0015924799999999999 0 0.00159258 3.3 0.0015925 3.3 0.0015926 0 0.0015925199999999998 0 0.0015926199999999999 3.3 0.00159254 3.3 0.00159264 0 0.0015925599999999998 0 0.0015926599999999999 3.3 0.00159258 3.3 0.00159268 0 0.0015926 0 0.0015927 3.3 0.0015926199999999999 3.3 0.00159272 0 0.00159264 0 0.00159274 3.3 0.0015926599999999999 3.3 0.00159276 0 0.00159268 0 0.00159278 3.3 0.0015926999999999998 3.3 0.0015928 0 0.00159272 0 0.00159282 3.3 0.0015927399999999998 3.3 0.0015928399999999999 0 0.00159276 0 0.00159286 3.3 0.0015927799999999998 3.3 0.0015928799999999999 0 0.0015928 0 0.0015929 3.3 0.00159282 3.3 0.00159292 0 0.0015928399999999999 0 0.00159294 3.3 0.00159286 3.3 0.00159296 0 0.0015928799999999999 0 0.00159298 3.3 0.0015929 3.3 0.001593 0 0.0015929199999999998 0 0.00159302 3.3 0.00159294 3.3 0.00159304 0 0.0015929599999999998 0 0.0015930599999999999 3.3 0.00159298 3.3 0.00159308 0 0.001593 0 0.0015931 3.3 0.00159302 3.3 0.00159312 0 0.00159304 0 0.00159314 3.3 0.0015930599999999999 3.3 0.00159316 0 0.00159308 0 0.00159318 3.3 0.0015930999999999999 3.3 0.0015932 0 0.00159312 0 0.00159322 3.3 0.0015931399999999998 3.3 0.0015932399999999999 0 0.00159316 0 0.00159326 3.3 0.0015931799999999998 3.3 0.0015932799999999999 0 0.0015932 0 0.0015933 3.3 0.00159322 3.3 0.00159332 0 0.0015932399999999999 0 0.00159334 3.3 0.00159326 3.3 0.00159336 0 0.0015932799999999999 0 0.00159338 3.3 0.0015933 3.3 0.0015934 0 0.0015933199999999998 0 0.00159342 3.3 0.00159334 3.3 0.00159344 0 0.0015933599999999998 0 0.0015934599999999999 3.3 0.00159338 3.3 0.00159348 0 0.0015933999999999998 0 0.0015934999999999999 3.3 0.00159342 3.3 0.00159352 0 0.00159344 0 0.00159354 3.3 0.0015934599999999999 3.3 0.00159356 0 0.00159348 0 0.00159358 3.3 0.0015934999999999999 3.3 0.0015936 0 0.00159352 0 0.00159362 3.3 0.0015935399999999998 3.3 0.00159364 0 0.00159356 0 0.00159366 3.3 0.0015935799999999998 3.3 0.0015936799999999999 0 0.0015936 0 0.0015937 3.3 0.00159362 3.3 0.00159372 0 0.00159364 0 0.00159374 3.3 0.00159366 3.3 0.00159376 0 0.0015936799999999999 0 0.00159378 3.3 0.0015937 3.3 0.0015938 0 0.0015937199999999999 0 0.00159382 3.3 0.00159374 3.3 0.00159384 0 0.0015937599999999998 0 0.00159386 3.3 0.00159378 3.3 0.00159388 0 0.0015937999999999998 0 0.0015938999999999999 3.3 0.00159382 3.3 0.00159392 0 0.00159384 0 0.00159394 3.3 0.00159386 3.3 0.00159396 0 0.00159388 0 0.00159398 3.3 0.0015938999999999999 3.3 0.001594 0 0.00159392 0 0.00159402 3.3 0.0015939399999999999 3.3 0.00159404 0 0.00159396 0 0.00159406 3.3 0.0015939799999999998 3.3 0.0015940799999999999 0 0.001594 0 0.0015941 3.3 0.0015940199999999998 3.3 0.0015941199999999999 0 0.00159404 0 0.00159414 3.3 0.00159406 3.3 0.00159416 0 0.0015940799999999999 0 0.00159418 3.3 0.0015941 3.3 0.0015942 0 0.0015941199999999999 0 0.00159422 3.3 0.00159414 3.3 0.00159424 0 0.0015941599999999998 0 0.00159426 3.3 0.00159418 3.3 0.00159428 0 0.0015941999999999998 0 0.0015942999999999999 3.3 0.00159422 3.3 0.00159432 0 0.0015942399999999998 0 0.0015943399999999999 3.3 0.00159426 3.3 0.00159436 0 0.00159428 0 0.00159438 3.3 0.0015942999999999999 3.3 0.0015944 0 0.00159432 0 0.00159442 3.3 0.0015943399999999999 3.3 0.00159444 0 0.00159436 0 0.00159446 3.3 0.0015943799999999998 3.3 0.00159448 0 0.0015944 0 0.0015945 3.3 0.0015944199999999998 3.3 0.0015945199999999999 0 0.00159444 0 0.00159454 3.3 0.00159446 3.3 0.00159456 0 0.00159448 0 0.00159458 3.3 0.0015945 3.3 0.0015946 0 0.0015945199999999999 0 0.00159462 3.3 0.00159454 3.3 0.00159464 0 0.0015945599999999999 0 0.00159466 3.3 0.00159458 3.3 0.00159468 0 0.0015945999999999998 0 0.0015947 3.3 0.00159462 3.3 0.00159472 0 0.0015946399999999998 0 0.0015947399999999999 3.3 0.00159466 3.3 0.00159476 0 0.00159468 0 0.00159478 3.3 0.0015947 3.3 0.0015948 0 0.00159472 0 0.00159482 3.3 0.0015947399999999999 3.3 0.00159484 0 0.00159476 0 0.00159486 3.3 0.0015947799999999999 3.3 0.00159488 0 0.0015948 0 0.0015949 3.3 0.0015948199999999998 3.3 0.0015949199999999999 0 0.00159484 0 0.00159494 3.3 0.0015948599999999998 3.3 0.0015949599999999999 0 0.00159488 0 0.00159498 3.3 0.0015949 3.3 0.001595 0 0.0015949199999999999 0 0.00159502 3.3 0.00159494 3.3 0.00159504 0 0.0015949599999999999 0 0.00159506 3.3 0.00159498 3.3 0.00159508 0 0.0015949999999999998 0 0.0015951 3.3 0.00159502 3.3 0.00159512 0 0.0015950399999999998 0 0.0015951399999999999 3.3 0.00159506 3.3 0.00159516 0 0.0015950799999999998 0 0.0015951799999999999 3.3 0.0015951 3.3 0.0015952 0 0.00159512 0 0.00159522 3.3 0.0015951399999999999 3.3 0.00159524 0 0.00159516 0 0.00159526 3.3 0.0015951799999999999 3.3 0.00159528 0 0.0015952 0 0.0015953 3.3 0.0015952199999999998 3.3 0.00159532 0 0.00159524 0 0.00159534 3.3 0.0015952599999999998 3.3 0.0015953599999999999 0 0.00159528 0 0.00159538 3.3 0.0015953 3.3 0.0015954 0 0.00159532 0 0.00159542 3.3 0.00159534 3.3 0.00159544 0 0.0015953599999999999 0 0.00159546 3.3 0.00159538 3.3 0.00159548 0 0.0015953999999999999 0 0.0015955 3.3 0.00159542 3.3 0.00159552 0 0.0015954399999999998 0 0.00159554 3.3 0.00159546 3.3 0.00159556 0 0.0015954799999999998 0 0.0015955799999999999 3.3 0.0015955 3.3 0.0015956 0 0.00159552 0 0.00159562 3.3 0.00159554 3.3 0.00159564 0 0.00159556 0 0.00159566 3.3 0.0015955799999999999 3.3 0.00159568 0 0.0015956 0 0.0015957 3.3 0.0015956199999999999 3.3 0.00159572 0 0.00159564 0 0.00159574 3.3 0.0015956599999999998 3.3 0.0015957599999999999 0 0.00159568 0 0.00159578 3.3 0.0015956999999999998 3.3 0.0015957999999999999 0 0.00159572 0 0.00159582 3.3 0.00159574 3.3 0.00159584 0 0.0015957599999999999 0 0.00159586 3.3 0.00159578 3.3 0.00159588 0 0.0015957999999999999 0 0.0015959 3.3 0.00159582 3.3 0.00159592 0 0.0015958399999999998 0 0.00159594 3.3 0.00159586 3.3 0.00159596 0 0.0015958799999999998 0 0.0015959799999999999 3.3 0.0015959 3.3 0.001596 0 0.0015959199999999998 0 0.0015960199999999999 3.3 0.00159594 3.3 0.00159604 0 0.00159596 0 0.00159606 3.3 0.0015959799999999999 3.3 0.00159608 0 0.001596 0 0.0015961 3.3 0.0015960199999999999 3.3 0.00159612 0 0.00159604 0 0.00159614 3.3 0.0015960599999999998 3.3 0.00159616 0 0.00159608 0 0.00159618 3.3 0.0015960999999999998 3.3 0.0015961999999999999 0 0.00159612 0 0.00159622 3.3 0.00159614 3.3 0.00159624 0 0.00159616 0 0.00159626 3.3 0.00159618 3.3 0.00159628 0 0.0015961999999999999 0 0.0015963 3.3 0.00159622 3.3 0.00159632 0 0.0015962399999999999 0 0.00159634 3.3 0.00159626 3.3 0.00159636 0 0.0015962799999999998 0 0.0015963799999999999 3.3 0.0015963 3.3 0.0015964 0 0.0015963199999999998 0 0.0015964199999999999 3.3 0.00159634 3.3 0.00159644 0 0.00159636 0 0.00159646 3.3 0.0015963799999999999 3.3 0.00159648 0 0.0015964 0 0.0015965 3.3 0.0015964199999999999 3.3 0.00159652 0 0.00159644 0 0.00159654 3.3 0.0015964599999999998 3.3 0.00159656 0 0.00159648 0 0.00159658 3.3 0.0015964999999999998 3.3 0.0015965999999999999 0 0.00159652 0 0.00159662 3.3 0.0015965399999999998 3.3 0.0015966399999999999 0 0.00159656 0 0.00159666 3.3 0.00159658 3.3 0.00159668 0 0.0015965999999999999 0 0.0015967 3.3 0.00159662 3.3 0.00159672 0 0.0015966399999999999 0 0.00159674 3.3 0.00159666 3.3 0.00159676 0 0.0015966799999999998 0 0.00159678 3.3 0.0015967 3.3 0.0015968 0 0.0015967199999999998 0 0.0015968199999999999 3.3 0.00159674 3.3 0.00159684 0 0.00159676 0 0.00159686 3.3 0.00159678 3.3 0.00159688 0 0.0015968 0 0.0015969 3.3 0.0015968199999999999 3.3 0.00159692 0 0.00159684 0 0.00159694 3.3 0.0015968599999999999 3.3 0.00159696 0 0.00159688 0 0.00159698 3.3 0.0015968999999999998 3.3 0.001597 0 0.00159692 0 0.00159702 3.3 0.0015969399999999998 3.3 0.0015970399999999999 0 0.00159696 0 0.00159706 3.3 0.00159698 3.3 0.00159708 0 0.001597 0 0.0015971 3.3 0.00159702 3.3 0.00159712 0 0.0015970399999999999 0 0.00159714 3.3 0.00159706 3.3 0.00159716 0 0.0015970799999999999 0 0.00159718 3.3 0.0015971 3.3 0.0015972 0 0.0015971199999999998 0 0.0015972199999999999 3.3 0.00159714 3.3 0.00159724 0 0.0015971599999999998 0 0.0015972599999999999 3.3 0.00159718 3.3 0.00159728 0 0.0015972 0 0.0015973 3.3 0.0015972199999999999 3.3 0.00159732 0 0.00159724 0 0.00159734 3.3 0.0015972599999999999 3.3 0.00159736 0 0.00159728 0 0.00159738 3.3 0.0015972999999999998 3.3 0.0015974 0 0.00159732 0 0.00159742 3.3 0.0015973399999999998 3.3 0.0015974399999999999 0 0.00159736 0 0.00159746 3.3 0.0015973799999999998 3.3 0.0015974799999999999 0 0.0015974 0 0.0015975 3.3 0.00159742 3.3 0.00159752 0 0.0015974399999999999 0 0.00159754 3.3 0.00159746 3.3 0.00159756 0 0.0015974799999999999 0 0.00159758 3.3 0.0015975 3.3 0.0015976 0 0.0015975199999999998 0 0.00159762 3.3 0.00159754 3.3 0.00159764 0 0.0015975599999999998 0 0.0015976599999999999 3.3 0.00159758 3.3 0.00159768 0 0.0015976 0 0.0015977 3.3 0.00159762 3.3 0.00159772 0 0.00159764 0 0.00159774 3.3 0.0015976599999999999 3.3 0.00159776 0 0.00159768 0 0.00159778 3.3 0.0015976999999999999 3.3 0.0015978 0 0.00159772 0 0.00159782 3.3 0.0015977399999999998 3.3 0.00159784 0 0.00159776 0 0.00159786 3.3 0.0015977799999999998 3.3 0.0015978799999999999 0 0.0015978 0 0.0015979 3.3 0.00159782 3.3 0.00159792 0 0.00159784 0 0.00159794 3.3 0.00159786 3.3 0.00159796 0 0.0015978799999999999 0 0.00159798 3.3 0.0015979 3.3 0.001598 0 0.0015979199999999999 0 0.00159802 3.3 0.00159794 3.3 0.00159804 0 0.0015979599999999998 0 0.0015980599999999999 3.3 0.00159798 3.3 0.00159808 0 0.0015979999999999998 0 0.0015980999999999999 3.3 0.00159802 3.3 0.00159812 0 0.00159804 0 0.00159814 3.3 0.0015980599999999999 3.3 0.00159816 0 0.00159808 0 0.00159818 3.3 0.0015980999999999999 3.3 0.0015982 0 0.00159812 0 0.00159822 3.3 0.0015981399999999998 3.3 0.00159824 0 0.00159816 0 0.00159826 3.3 0.0015981799999999998 3.3 0.0015982799999999999 0 0.0015982 0 0.0015983 3.3 0.0015982199999999998 3.3 0.0015983199999999999 0 0.00159824 0 0.00159834 3.3 0.00159826 3.3 0.00159836 0 0.0015982799999999999 0 0.00159838 3.3 0.0015983 3.3 0.0015984 0 0.0015983199999999999 0 0.00159842 3.3 0.00159834 3.3 0.00159844 0 0.0015983599999999998 0 0.00159846 3.3 0.00159838 3.3 0.00159848 0 0.0015983999999999998 0 0.0015984999999999999 3.3 0.00159842 3.3 0.00159852 0 0.00159844 0 0.00159854 3.3 0.00159846 3.3 0.00159856 0 0.00159848 0 0.00159858 3.3 0.0015984999999999999 3.3 0.0015986 0 0.00159852 0 0.00159862 3.3 0.0015985399999999999 3.3 0.00159864 0 0.00159856 0 0.00159866 3.3 0.0015985799999999998 3.3 0.00159868 0 0.0015986 0 0.0015987 3.3 0.0015986199999999998 3.3 0.0015987199999999999 0 0.00159864 0 0.00159874 3.3 0.00159866 3.3 0.00159876 0 0.00159868 0 0.00159878 3.3 0.0015987 3.3 0.0015988 0 0.0015987199999999999 0 0.00159882 3.3 0.00159874 3.3 0.00159884 0 0.0015987599999999999 0 0.00159886 3.3 0.00159878 3.3 0.00159888 0 0.0015987999999999998 0 0.0015988999999999999 3.3 0.00159882 3.3 0.00159892 0 0.0015988399999999998 0 0.0015989399999999999 3.3 0.00159886 3.3 0.00159896 0 0.00159888 0 0.00159898 3.3 0.0015988999999999999 3.3 0.001599 0 0.00159892 0 0.00159902 3.3 0.0015989399999999999 3.3 0.00159904 0 0.00159896 0 0.00159906 3.3 0.0015989799999999998 3.3 0.00159908 0 0.001599 0 0.0015991 3.3 0.0015990199999999998 3.3 0.0015991199999999999 0 0.00159904 0 0.00159914 3.3 0.0015990599999999998 3.3 0.0015991599999999999 0 0.00159908 0 0.00159918 3.3 0.0015991 3.3 0.0015992 0 0.0015991199999999999 0 0.00159922 3.3 0.00159914 3.3 0.00159924 0 0.0015991599999999999 0 0.00159926 3.3 0.00159918 3.3 0.00159928 0 0.0015991999999999998 0 0.0015993 3.3 0.00159922 3.3 0.00159932 0 0.0015992399999999998 0 0.0015993399999999999 3.3 0.00159926 3.3 0.00159936 0 0.00159928 0 0.00159938 3.3 0.0015993 3.3 0.0015994 0 0.00159932 0 0.00159942 3.3 0.0015993399999999999 3.3 0.00159944 0 0.00159936 0 0.00159946 3.3 0.0015993799999999999 3.3 0.00159948 0 0.0015994 0 0.0015995 3.3 0.0015994199999999998 3.3 0.0015995199999999999 0 0.00159944 0 0.00159954 3.3 0.0015994599999999998 3.3 0.0015995599999999999 0 0.00159948 0 0.00159958 3.3 0.0015995 3.3 0.0015996 0 0.0015995199999999999 0 0.00159962 3.3 0.00159954 3.3 0.00159964 0 0.0015995599999999999 0 0.00159966 3.3 0.00159958 3.3 0.00159968 0 0.0015995999999999999 0 0.0015997 3.3 0.00159962 3.3 0.00159972 0 0.0015996399999999998 0 0.0015997399999999999 3.3 0.00159966 3.3 0.00159976 0 0.0015996799999999998 0 0.0015997799999999999 3.3 0.0015997 3.3 0.0015998 0 0.00159972 0 0.00159982 3.3 0.0015997399999999999 3.3 0.00159984 0 0.00159976 0 0.00159986 3.3 0.0015997799999999999 3.3 0.00159988 0 0.0015998 0 0.0015999 3.3 0.0015998199999999998 3.3 0.00159992 0 0.00159984 0 0.00159994 3.3 0.0015998599999999998 3.3 0.0015999599999999999 0 0.00159988 0 0.00159998 3.3 0.0015998999999999998 3.3 0.0015999999999999999 0 0.00159992 0 0.00160002 3.3 0.00159994 3.3 0.00160004 0 0.0015999599999999999 0 0.00160006 3.3 0.00159998 3.3 0.00160008 0 0.0015999999999999999 0 0.0016001 3.3 0.00160002 3.3 0.00160012 0 0.0016000399999999998 0 0.00160014 3.3 0.00160006 3.3 0.00160016 0 0.0016000799999999998 0 0.0016001799999999999 3.3 0.0016001 3.3 0.0016002 0 0.00160012 0 0.00160022 3.3 0.00160014 3.3 0.00160024 0 0.00160016 0 0.00160026 3.3 0.0016001799999999999 3.3 0.00160028 0 0.0016002 0 0.0016003 3.3 0.0016002199999999999 3.3 0.00160032 0 0.00160024 0 0.00160034 3.3 0.0016002599999999998 3.3 0.0016003599999999999 0 0.00160028 0 0.00160038 3.3 0.0016002999999999998 3.3 0.0016003999999999999 0 0.00160032 0 0.00160042 3.3 0.00160034 3.3 0.00160044 0 0.0016003599999999999 0 0.00160046 3.3 0.00160038 3.3 0.00160048 0 0.0016003999999999999 0 0.0016005 3.3 0.00160042 3.3 0.00160052 0 0.0016004399999999998 0 0.00160054 3.3 0.00160046 3.3 0.00160056 0 0.0016004799999999998 0 0.0016005799999999999 3.3 0.0016005 3.3 0.0016006 0 0.0016005199999999998 0 0.0016006199999999999 3.3 0.00160054 3.3 0.00160064 0 0.00160056 0 0.00160066 3.3 0.0016005799999999999 3.3 0.00160068 0 0.0016006 0 0.0016007 3.3 0.0016006199999999999 3.3 0.00160072 0 0.00160064 0 0.00160074 3.3 0.0016006599999999998 3.3 0.00160076 0 0.00160068 0 0.00160078 3.3 0.0016006999999999998 3.3 0.0016007999999999999 0 0.00160072 0 0.00160082 3.3 0.00160074 3.3 0.00160084 0 0.00160076 0 0.00160086 3.3 0.00160078 3.3 0.00160088 0 0.0016007999999999999 0 0.0016009 3.3 0.00160082 3.3 0.00160092 0 0.0016008399999999999 0 0.00160094 3.3 0.00160086 3.3 0.00160096 0 0.0016008799999999998 0 0.00160098 3.3 0.0016009 3.3 0.001601 0 0.0016009199999999998 0 0.0016010199999999999 3.3 0.00160094 3.3 0.00160104 0 0.00160096 0 0.00160106 3.3 0.00160098 3.3 0.00160108 0 0.001601 0 0.0016011 3.3 0.0016010199999999999 3.3 0.00160112 0 0.00160104 0 0.00160114 3.3 0.0016010599999999999 3.3 0.00160116 0 0.00160108 0 0.00160118 3.3 0.0016010999999999998 3.3 0.0016011999999999999 0 0.00160112 0 0.00160122 3.3 0.0016011399999999998 3.3 0.0016012399999999999 0 0.00160116 0 0.00160126 3.3 0.00160118 3.3 0.00160128 0 0.0016011999999999999 0 0.0016013 3.3 0.00160122 3.3 0.00160132 0 0.0016012399999999999 0 0.00160134 3.3 0.00160126 3.3 0.00160136 0 0.0016012799999999998 0 0.00160138 3.3 0.0016013 3.3 0.0016014 0 0.0016013199999999998 0 0.0016014199999999999 3.3 0.00160134 3.3 0.00160144 0 0.0016013599999999998 0 0.0016014599999999999 3.3 0.00160138 3.3 0.00160148 0 0.0016014 0 0.0016015 3.3 0.0016014199999999999 3.3 0.00160152 0 0.00160144 0 0.00160154 3.3 0.0016014599999999999 3.3 0.00160156 0 0.00160148 0 0.00160158 3.3 0.0016014999999999998 3.3 0.0016016 0 0.00160152 0 0.00160162 3.3 0.0016015399999999998 3.3 0.0016016399999999999 0 0.00160156 0 0.00160166 3.3 0.00160158 3.3 0.00160168 0 0.0016016 0 0.0016017 3.3 0.00160162 3.3 0.00160172 0 0.0016016399999999999 0 0.00160174 3.3 0.00160166 3.3 0.00160176 0 0.0016016799999999999 0 0.00160178 3.3 0.0016017 3.3 0.0016018 0 0.0016017199999999998 0 0.00160182 3.3 0.00160174 3.3 0.00160184 0 0.0016017599999999998 0 0.0016018599999999999 3.3 0.00160178 3.3 0.00160188 0 0.0016018 0 0.0016019 3.3 0.00160182 3.3 0.00160192 0 0.00160184 0 0.00160194 3.3 0.0016018599999999999 3.3 0.00160196 0 0.00160188 0 0.00160198 3.3 0.0016018999999999999 3.3 0.001602 0 0.00160192 0 0.00160202 3.3 0.0016019399999999998 3.3 0.0016020399999999999 0 0.00160196 0 0.00160206 3.3 0.0016019799999999998 3.3 0.0016020799999999999 0 0.001602 0 0.0016021 3.3 0.00160202 3.3 0.00160212 0 0.0016020399999999999 0 0.00160214 3.3 0.00160206 3.3 0.00160216 0 0.0016020799999999999 0 0.00160218 3.3 0.0016021 3.3 0.0016022 0 0.0016021199999999998 0 0.00160222 3.3 0.00160214 3.3 0.00160224 0 0.0016021599999999998 0 0.0016022599999999999 3.3 0.00160218 3.3 0.00160228 0 0.0016021999999999998 0 0.0016022999999999999 3.3 0.00160222 3.3 0.00160232 0 0.00160224 0 0.00160234 3.3 0.0016022599999999999 3.3 0.00160236 0 0.00160228 0 0.00160238 3.3 0.0016022999999999999 3.3 0.0016024 0 0.00160232 0 0.00160242 3.3 0.0016023399999999998 3.3 0.00160244 0 0.00160236 0 0.00160246 3.3 0.0016023799999999998 3.3 0.0016024799999999999 0 0.0016024 0 0.0016025 3.3 0.00160242 3.3 0.00160252 0 0.00160244 0 0.00160254 3.3 0.00160246 3.3 0.00160256 0 0.0016024799999999999 0 0.00160258 3.3 0.0016025 3.3 0.0016026 0 0.0016025199999999999 0 0.00160262 3.3 0.00160254 3.3 0.00160264 0 0.0016025599999999998 0 0.00160266 3.3 0.00160258 3.3 0.00160268 0 0.0016025999999999998 0 0.0016026999999999999 3.3 0.00160262 3.3 0.00160272 0 0.00160264 0 0.00160274 3.3 0.00160266 3.3 0.00160276 0 0.00160268 0 0.00160278 3.3 0.0016026999999999999 3.3 0.0016028 0 0.00160272 0 0.00160282 3.3 0.0016027399999999999 3.3 0.00160284 0 0.00160276 0 0.00160286 3.3 0.0016027799999999998 3.3 0.0016028799999999999 0 0.0016028 0 0.0016029 3.3 0.0016028199999999998 3.3 0.0016029199999999999 0 0.00160284 0 0.00160294 3.3 0.00160286 3.3 0.00160296 0 0.0016028799999999999 0 0.00160298 3.3 0.0016029 3.3 0.001603 0 0.0016029199999999999 0 0.00160302 3.3 0.00160294 3.3 0.00160304 0 0.0016029599999999998 0 0.00160306 3.3 0.00160298 3.3 0.00160308 0 0.0016029999999999998 0 0.0016030999999999999 3.3 0.00160302 3.3 0.00160312 0 0.0016030399999999998 0 0.0016031399999999999 3.3 0.00160306 3.3 0.00160316 0 0.00160308 0 0.00160318 3.3 0.0016030999999999999 3.3 0.0016032 0 0.00160312 0 0.00160322 3.3 0.0016031399999999999 3.3 0.00160324 0 0.00160316 0 0.00160326 3.3 0.0016031799999999998 3.3 0.00160328 0 0.0016032 0 0.0016033 3.3 0.0016032199999999998 3.3 0.0016033199999999999 0 0.00160324 0 0.00160334 3.3 0.00160326 3.3 0.00160336 0 0.00160328 0 0.00160338 3.3 0.0016033 3.3 0.0016034 0 0.0016033199999999999 0 0.00160342 3.3 0.00160334 3.3 0.00160344 0 0.0016033599999999999 0 0.00160346 3.3 0.00160338 3.3 0.00160348 0 0.0016033999999999998 0 0.0016034999999999999 3.3 0.00160342 3.3 0.00160352 0 0.0016034399999999998 0 0.0016035399999999999 3.3 0.00160346 3.3 0.00160356 0 0.00160348 0 0.00160358 3.3 0.0016034999999999999 3.3 0.0016036 0 0.00160352 0 0.00160362 3.3 0.0016035399999999999 3.3 0.00160364 0 0.00160356 0 0.00160366 3.3 0.0016035799999999998 3.3 0.00160368 0 0.0016036 0 0.0016037 3.3 0.0016036199999999998 3.3 0.0016037199999999999 0 0.00160364 0 0.00160374 3.3 0.0016036599999999998 3.3 0.0016037599999999999 0 0.00160368 0 0.00160378 3.3 0.0016037 3.3 0.0016038 0 0.0016037199999999999 0 0.00160382 3.3 0.00160374 3.3 0.00160384 0 0.0016037599999999999 0 0.00160386 3.3 0.00160378 3.3 0.00160388 0 0.0016037999999999998 0 0.0016039 3.3 0.00160382 3.3 0.00160392 0 0.0016038399999999998 0 0.0016039399999999999 3.3 0.00160386 3.3 0.00160396 0 0.00160388 0 0.00160398 3.3 0.0016039 3.3 0.001604 0 0.00160392 0 0.00160402 3.3 0.0016039399999999999 3.3 0.00160404 0 0.00160396 0 0.00160406 3.3 0.0016039799999999999 3.3 0.00160408 0 0.001604 0 0.0016041 3.3 0.0016040199999999998 3.3 0.00160412 0 0.00160404 0 0.00160414 3.3 0.0016040599999999998 3.3 0.0016041599999999999 0 0.00160408 0 0.00160418 3.3 0.0016041 3.3 0.0016042 0 0.00160412 0 0.00160422 3.3 0.00160414 3.3 0.00160424 0 0.0016041599999999999 0 0.00160426 3.3 0.00160418 3.3 0.00160428 0 0.0016041999999999999 0 0.0016043 3.3 0.00160422 3.3 0.00160432 0 0.0016042399999999998 0 0.0016043399999999999 3.3 0.00160426 3.3 0.00160436 0 0.0016042799999999998 0 0.0016043799999999999 3.3 0.0016043 3.3 0.0016044 0 0.00160432 0 0.00160442 3.3 0.0016043399999999999 3.3 0.00160444 0 0.00160436 0 0.00160446 3.3 0.0016043799999999999 3.3 0.00160448 0 0.0016044 0 0.0016045 3.3 0.0016044199999999998 3.3 0.00160452 0 0.00160444 0 0.00160454 3.3 0.0016044599999999998 3.3 0.0016045599999999999 0 0.00160448 0 0.00160458 3.3 0.0016044999999999998 3.3 0.0016045999999999999 0 0.00160452 0 0.00160462 3.3 0.00160454 3.3 0.00160464 0 0.0016045599999999999 0 0.00160466 3.3 0.00160458 3.3 0.00160468 0 0.0016045999999999999 0 0.0016047 3.3 0.00160462 3.3 0.00160472 0 0.0016046399999999998 0 0.00160474 3.3 0.00160466 3.3 0.00160476 0 0.0016046799999999998 0 0.0016047799999999999 3.3 0.0016047 3.3 0.0016048 0 0.00160472 0 0.00160482 3.3 0.00160474 3.3 0.00160484 0 0.00160476 0 0.00160486 3.3 0.0016047799999999999 3.3 0.00160488 0 0.0016048 0 0.0016049 3.3 0.0016048199999999999 3.3 0.00160492 0 0.00160484 0 0.00160494 3.3 0.0016048599999999998 3.3 0.00160496 0 0.00160488 0 0.00160498 3.3 0.0016048999999999998 3.3 0.0016049999999999999 0 0.00160492 0 0.00160502 3.3 0.00160494 3.3 0.00160504 0 0.00160496 0 0.00160506 3.3 0.00160498 3.3 0.00160508 0 0.0016049999999999999 0 0.0016051 3.3 0.00160502 3.3 0.00160512 0 0.0016050399999999999 0 0.00160514 3.3 0.00160506 3.3 0.00160516 0 0.0016050799999999998 0 0.0016051799999999999 3.3 0.0016051 3.3 0.0016052 0 0.0016051199999999998 0 0.0016052199999999999 3.3 0.00160514 3.3 0.00160524 0 0.00160516 0 0.00160526 3.3 0.0016051799999999999 3.3 0.00160528 0 0.0016052 0 0.0016053 3.3 0.0016052199999999999 3.3 0.00160532 0 0.00160524 0 0.00160534 3.3 0.0016052599999999998 3.3 0.00160536 0 0.00160528 0 0.00160538 3.3 0.0016052999999999998 3.3 0.0016053999999999999 0 0.00160532 0 0.00160542 3.3 0.0016053399999999998 3.3 0.0016054399999999999 0 0.00160536 0 0.00160546 3.3 0.00160538 3.3 0.00160548 0 0.0016053999999999999 0 0.0016055 3.3 0.00160542 3.3 0.00160552 0 0.0016054399999999999 0 0.00160554 3.3 0.00160546 3.3 0.00160556 0 0.0016054799999999998 0 0.00160558 3.3 0.0016055 3.3 0.0016056 0 0.0016055199999999998 0 0.0016056199999999999 3.3 0.00160554 3.3 0.00160564 0 0.00160556 0 0.00160566 3.3 0.00160558 3.3 0.00160568 0 0.0016056 0 0.0016057 3.3 0.0016056199999999999 3.3 0.00160572 0 0.00160564 0 0.00160574 3.3 0.0016056599999999999 3.3 0.00160576 0 0.00160568 0 0.00160578 3.3 0.0016056999999999998 3.3 0.0016058 0 0.00160572 0 0.00160582 3.3 0.0016057399999999998 3.3 0.0016058399999999999 0 0.00160576 0 0.00160586 3.3 0.00160578 3.3 0.00160588 0 0.0016058 0 0.0016059 3.3 0.00160582 3.3 0.00160592 0 0.0016058399999999999 0 0.00160594 3.3 0.00160586 3.3 0.00160596 0 0.0016058799999999999 0 0.00160598 3.3 0.0016059 3.3 0.001606 0 0.0016059199999999998 0 0.0016060199999999999 3.3 0.00160594 3.3 0.00160604 0 0.0016059599999999998 0 0.0016060599999999999 3.3 0.00160598 3.3 0.00160608 0 0.001606 0 0.0016061 3.3 0.0016060199999999999 3.3 0.00160612 0 0.00160604 0 0.00160614 3.3 0.0016060599999999999 3.3 0.00160616 0 0.00160608 0 0.00160618 3.3 0.0016060999999999998 3.3 0.0016062 0 0.00160612 0 0.00160622 3.3 0.0016061399999999998 3.3 0.0016062399999999999 0 0.00160616 0 0.00160626 3.3 0.0016061799999999998 3.3 0.0016062799999999999 0 0.0016062 0 0.0016063 3.3 0.00160622 3.3 0.00160632 0 0.0016062399999999999 0 0.00160634 3.3 0.00160626 3.3 0.00160636 0 0.0016062799999999999 0 0.00160638 3.3 0.0016063 3.3 0.0016064 0 0.0016063199999999998 0 0.00160642 3.3 0.00160634 3.3 0.00160644 0 0.0016063599999999998 0 0.0016064599999999999 3.3 0.00160638 3.3 0.00160648 0 0.0016064 0 0.0016065 3.3 0.00160642 3.3 0.00160652 0 0.00160644 0 0.00160654 3.3 0.0016064599999999999 3.3 0.00160656 0 0.00160648 0 0.00160658 3.3 0.0016064999999999999 3.3 0.0016066 0 0.00160652 0 0.00160662 3.3 0.0016065399999999998 3.3 0.0016066399999999999 0 0.00160656 0 0.00160666 3.3 0.0016065799999999998 3.3 0.0016066799999999999 0 0.0016066 0 0.0016067 3.3 0.00160662 3.3 0.00160672 0 0.0016066399999999999 0 0.00160674 3.3 0.00160666 3.3 0.00160676 0 0.0016066799999999999 0 0.00160678 3.3 0.0016067 3.3 0.0016068 0 0.0016067199999999998 0 0.00160682 3.3 0.00160674 3.3 0.00160684 0 0.0016067599999999998 0 0.0016068599999999999 3.3 0.00160678 3.3 0.00160688 0 0.0016067999999999998 0 0.0016068999999999999 3.3 0.00160682 3.3 0.00160692 0 0.00160684 0 0.00160694 3.3 0.0016068599999999999 3.3 0.00160696 0 0.00160688 0 0.00160698 3.3 0.0016068999999999999 3.3 0.001607 0 0.00160692 0 0.00160702 3.3 0.0016069399999999998 3.3 0.00160704 0 0.00160696 0 0.00160706 3.3 0.0016069799999999998 3.3 0.0016070799999999999 0 0.001607 0 0.0016071 3.3 0.0016070199999999998 3.3 0.0016071199999999999 0 0.00160704 0 0.00160714 3.3 0.00160706 3.3 0.00160716 0 0.0016070799999999999 0 0.00160718 3.3 0.0016071 3.3 0.0016072 0 0.0016071199999999999 0 0.00160722 3.3 0.00160714 3.3 0.00160724 0 0.0016071599999999998 0 0.00160726 3.3 0.00160718 3.3 0.00160728 0 0.0016071999999999998 0 0.0016072999999999999 3.3 0.00160722 3.3 0.00160732 0 0.00160724 0 0.00160734 3.3 0.00160726 3.3 0.00160736 0 0.00160728 0 0.00160738 3.3 0.0016072999999999999 3.3 0.0016074 0 0.00160732 0 0.00160742 3.3 0.0016073399999999999 3.3 0.00160744 0 0.00160736 0 0.00160746 3.3 0.0016073799999999998 3.3 0.0016074799999999999 0 0.0016074 0 0.0016075 3.3 0.0016074199999999998 3.3 0.0016075199999999999 0 0.00160744 0 0.00160754 3.3 0.00160746 3.3 0.00160756 0 0.0016074799999999999 0 0.00160758 3.3 0.0016075 3.3 0.0016076 0 0.0016075199999999999 0 0.00160762 3.3 0.00160754 3.3 0.00160764 0 0.0016075599999999998 0 0.00160766 3.3 0.00160758 3.3 0.00160768 0 0.0016075999999999998 0 0.0016076999999999999 3.3 0.00160762 3.3 0.00160772 0 0.0016076399999999998 0 0.0016077399999999999 3.3 0.00160766 3.3 0.00160776 0 0.00160768 0 0.00160778 3.3 0.0016076999999999999 3.3 0.0016078 0 0.00160772 0 0.00160782 3.3 0.0016077399999999999 3.3 0.00160784 0 0.00160776 0 0.00160786 3.3 0.0016077799999999998 3.3 0.00160788 0 0.0016078 0 0.0016079 3.3 0.0016078199999999998 3.3 0.0016079199999999999 0 0.00160784 0 0.00160794 3.3 0.00160786 3.3 0.00160796 0 0.00160788 0 0.00160798 3.3 0.0016079 3.3 0.001608 0 0.0016079199999999999 0 0.00160802 3.3 0.00160794 3.3 0.00160804 0 0.0016079599999999999 0 0.00160806 3.3 0.00160798 3.3 0.00160808 0 0.0016079999999999998 0 0.0016081 3.3 0.00160802 3.3 0.00160812 0 0.0016080399999999998 0 0.0016081399999999999 3.3 0.00160806 3.3 0.00160816 0 0.00160808 0 0.00160818 3.3 0.0016081 3.3 0.0016082 0 0.00160812 0 0.00160822 3.3 0.0016081399999999999 3.3 0.00160824 0 0.00160816 0 0.00160826 3.3 0.0016081799999999999 3.3 0.00160828 0 0.0016082 0 0.0016083 3.3 0.0016082199999999998 3.3 0.0016083199999999999 0 0.00160824 0 0.00160834 3.3 0.0016082599999999998 3.3 0.0016083599999999999 0 0.00160828 0 0.00160838 3.3 0.0016083 3.3 0.0016084 0 0.0016083199999999999 0 0.00160842 3.3 0.00160834 3.3 0.00160844 0 0.0016083599999999999 0 0.00160846 3.3 0.00160838 3.3 0.00160848 0 0.0016083999999999998 0 0.0016085 3.3 0.00160842 3.3 0.00160852 0 0.0016084399999999998 0 0.0016085399999999999 3.3 0.00160846 3.3 0.00160856 0 0.0016084799999999998 0 0.0016085799999999999 3.3 0.0016085 3.3 0.0016086 0 0.00160852 0 0.00160862 3.3 0.0016085399999999999 3.3 0.00160864 0 0.00160856 0 0.00160866 3.3 0.0016085799999999999 3.3 0.00160868 0 0.0016086 0 0.0016087 3.3 0.0016086199999999998 3.3 0.00160872 0 0.00160864 0 0.00160874 3.3 0.0016086599999999998 3.3 0.0016087599999999999 0 0.00160868 0 0.00160878 3.3 0.0016087 3.3 0.0016088 0 0.00160872 0 0.00160882 3.3 0.00160874 3.3 0.00160884 0 0.0016087599999999999 0 0.00160886 3.3 0.00160878 3.3 0.00160888 0 0.0016087999999999999 0 0.0016089 3.3 0.00160882 3.3 0.00160892 0 0.0016088399999999998 0 0.00160894 3.3 0.00160886 3.3 0.00160896 0 0.0016088799999999998 0 0.0016089799999999999 3.3 0.0016089 3.3 0.001609 0 0.00160892 0 0.00160902 3.3 0.00160894 3.3 0.00160904 0 0.00160896 0 0.00160906 3.3 0.0016089799999999999 3.3 0.00160908 0 0.001609 0 0.0016091 3.3 0.0016090199999999999 3.3 0.00160912 0 0.00160904 0 0.00160914 3.3 0.0016090599999999998 3.3 0.0016091599999999999 0 0.00160908 0 0.00160918 3.3 0.0016090999999999998 3.3 0.0016091999999999999 0 0.00160912 0 0.00160922 3.3 0.00160914 3.3 0.00160924 0 0.0016091599999999999 0 0.00160926 3.3 0.00160918 3.3 0.00160928 0 0.0016091999999999999 0 0.0016093 3.3 0.00160922 3.3 0.00160932 0 0.0016092399999999998 0 0.00160934 3.3 0.00160926 3.3 0.00160936 0 0.0016092799999999998 0 0.0016093799999999999 3.3 0.0016093 3.3 0.0016094 0 0.0016093199999999998 0 0.0016094199999999999 3.3 0.00160934 3.3 0.00160944 0 0.00160936 0 0.00160946 3.3 0.0016093799999999999 3.3 0.00160948 0 0.0016094 0 0.0016095 3.3 0.0016094199999999999 3.3 0.00160952 0 0.00160944 0 0.00160954 3.3 0.0016094599999999998 3.3 0.00160956 0 0.00160948 0 0.00160958 3.3 0.0016094999999999998 3.3 0.0016095999999999999 0 0.00160952 0 0.00160962 3.3 0.00160954 3.3 0.00160964 0 0.00160956 0 0.00160966 3.3 0.00160958 3.3 0.00160968 0 0.0016095999999999999 0 0.0016097 3.3 0.00160962 3.3 0.00160972 0 0.0016096399999999999 0 0.00160974 3.3 0.00160966 3.3 0.00160976 0 0.0016096799999999998 0 0.0016097799999999999 3.3 0.0016097 3.3 0.0016098 0 0.0016097199999999998 0 0.0016098199999999999 3.3 0.00160974 3.3 0.00160984 0 0.00160976 0 0.00160986 3.3 0.0016097799999999999 3.3 0.00160988 0 0.0016098 0 0.0016099 3.3 0.0016098199999999999 3.3 0.00160992 0 0.00160984 0 0.00160994 3.3 0.0016098599999999999 3.3 0.00160996 0 0.00160988 0 0.00160998 3.3 0.0016098999999999998 3.3 0.0016099999999999999 0 0.00160992 0 0.00161002 3.3 0.0016099399999999998 3.3 0.0016100399999999999 0 0.00160996 0 0.00161006 3.3 0.00160998 3.3 0.00161008 0 0.0016099999999999999 0 0.0016101 3.3 0.00161002 3.3 0.00161012 0 0.0016100399999999999 0 0.00161014 3.3 0.00161006 3.3 0.00161016 0 0.0016100799999999998 0 0.00161018 3.3 0.0016101 3.3 0.0016102 0 0.0016101199999999998 0 0.0016102199999999999 3.3 0.00161014 3.3 0.00161024 0 0.0016101599999999998 0 0.0016102599999999999 3.3 0.00161018 3.3 0.00161028 0 0.0016102 0 0.0016103 3.3 0.0016102199999999999 3.3 0.00161032 0 0.00161024 0 0.00161034 3.3 0.0016102599999999999 3.3 0.00161036 0 0.00161028 0 0.00161038 3.3 0.0016102999999999998 3.3 0.0016104 0 0.00161032 0 0.00161042 3.3 0.0016103399999999998 3.3 0.0016104399999999999 0 0.00161036 0 0.00161046 3.3 0.00161038 3.3 0.00161048 0 0.0016104 0 0.0016105 3.3 0.00161042 3.3 0.00161052 0 0.0016104399999999999 0 0.00161054 3.3 0.00161046 3.3 0.00161056 0 0.0016104799999999999 0 0.00161058 3.3 0.0016105 3.3 0.0016106 0 0.0016105199999999998 0 0.0016106199999999999 3.3 0.00161054 3.3 0.00161064 0 0.0016105599999999998 0 0.0016106599999999999 3.3 0.00161058 3.3 0.00161068 0 0.0016106 0 0.0016107 3.3 0.0016106199999999999 3.3 0.00161072 0 0.00161064 0 0.00161074 3.3 0.0016106599999999999 3.3 0.00161076 0 0.00161068 0 0.00161078 3.3 0.0016106999999999998 3.3 0.0016108 0 0.00161072 0 0.00161082 3.3 0.0016107399999999998 3.3 0.0016108399999999999 0 0.00161076 0 0.00161086 3.3 0.0016107799999999998 3.3 0.0016108799999999999 0 0.0016108 0 0.0016109 3.3 0.00161082 3.3 0.00161092 0 0.0016108399999999999 0 0.00161094 3.3 0.00161086 3.3 0.00161096 0 0.0016108799999999999 0 0.00161098 3.3 0.0016109 3.3 0.001611 0 0.0016109199999999998 0 0.00161102 3.3 0.00161094 3.3 0.00161104 0 0.0016109599999999998 0 0.0016110599999999999 3.3 0.00161098 3.3 0.00161108 0 0.001611 0 0.0016111 3.3 0.00161102 3.3 0.00161112 0 0.00161104 0 0.00161114 3.3 0.0016110599999999999 3.3 0.00161116 0 0.00161108 0 0.00161118 3.3 0.0016110999999999999 3.3 0.0016112 0 0.00161112 0 0.00161122 3.3 0.0016111399999999998 3.3 0.00161124 0 0.00161116 0 0.00161126 3.3 0.0016111799999999998 3.3 0.0016112799999999999 0 0.0016112 0 0.0016113 3.3 0.00161122 3.3 0.00161132 0 0.00161124 0 0.00161134 3.3 0.00161126 3.3 0.00161136 0 0.0016112799999999999 0 0.00161138 3.3 0.0016113 3.3 0.0016114 0 0.0016113199999999999 0 0.00161142 3.3 0.00161134 3.3 0.00161144 0 0.0016113599999999998 0 0.0016114599999999999 3.3 0.00161138 3.3 0.00161148 0 0.0016113999999999998 0 0.0016114999999999999 3.3 0.00161142 3.3 0.00161152 0 0.00161144 0 0.00161154 3.3 0.0016114599999999999 3.3 0.00161156 0 0.00161148 0 0.00161158 3.3 0.0016114999999999999 3.3 0.0016116 0 0.00161152 0 0.00161162 3.3 0.0016115399999999998 3.3 0.00161164 0 0.00161156 0 0.00161166 3.3 0.0016115799999999998 3.3 0.0016116799999999999 0 0.0016116 0 0.0016117 3.3 0.0016116199999999998 3.3 0.0016117199999999999 0 0.00161164 0 0.00161174 3.3 0.00161166 3.3 0.00161176 0 0.0016116799999999999 0 0.00161178 3.3 0.0016117 3.3 0.0016118 0 0.0016117199999999999 0 0.00161182 3.3 0.00161174 3.3 0.00161184 0 0.0016117599999999998 0 0.00161186 3.3 0.00161178 3.3 0.00161188 0 0.0016117999999999998 0 0.0016118999999999999 3.3 0.00161182 3.3 0.00161192 0 0.00161184 0 0.00161194 3.3 0.00161186 3.3 0.00161196 0 0.00161188 0 0.00161198 3.3 0.0016118999999999999 3.3 0.001612 0 0.00161192 0 0.00161202 3.3 0.0016119399999999999 3.3 0.00161204 0 0.00161196 0 0.00161206 3.3 0.0016119799999999998 3.3 0.00161208 0 0.001612 0 0.0016121 3.3 0.0016120199999999998 3.3 0.0016121199999999999 0 0.00161204 0 0.00161214 3.3 0.00161206 3.3 0.00161216 0 0.00161208 0 0.00161218 3.3 0.0016121 3.3 0.0016122 0 0.0016121199999999999 0 0.00161222 3.3 0.00161214 3.3 0.00161224 0 0.0016121599999999999 0 0.00161226 3.3 0.00161218 3.3 0.00161228 0 0.0016121999999999998 0 0.0016122999999999999 3.3 0.00161222 3.3 0.00161232 0 0.0016122399999999998 0 0.0016123399999999999 3.3 0.00161226 3.3 0.00161236 0 0.00161228 0 0.00161238 3.3 0.0016122999999999999 3.3 0.0016124 0 0.00161232 0 0.00161242 3.3 0.0016123399999999999 3.3 0.00161244 0 0.00161236 0 0.00161246 3.3 0.0016123799999999998 3.3 0.00161248 0 0.0016124 0 0.0016125 3.3 0.0016124199999999998 3.3 0.0016125199999999999 0 0.00161244 0 0.00161254 3.3 0.0016124599999999998 3.3 0.0016125599999999999 0 0.00161248 0 0.00161258 3.3 0.0016125 3.3 0.0016126 0 0.0016125199999999999 0 0.00161262 3.3 0.00161254 3.3 0.00161264 0 0.0016125599999999999 0 0.00161266 3.3 0.00161258 3.3 0.00161268 0 0.0016125999999999998 0 0.0016127 3.3 0.00161262 3.3 0.00161272 0 0.0016126399999999998 0 0.0016127399999999999 3.3 0.00161266 3.3 0.00161276 0 0.00161268 0 0.00161278 3.3 0.0016127 3.3 0.0016128 0 0.00161272 0 0.00161282 3.3 0.0016127399999999999 3.3 0.00161284 0 0.00161276 0 0.00161286 3.3 0.0016127799999999999 3.3 0.00161288 0 0.0016128 0 0.0016129 3.3 0.0016128199999999998 3.3 0.00161292 0 0.00161284 0 0.00161294 3.3 0.0016128599999999998 3.3 0.0016129599999999999 0 0.00161288 0 0.00161298 3.3 0.0016129 3.3 0.001613 0 0.00161292 0 0.00161302 3.3 0.00161294 3.3 0.00161304 0 0.0016129599999999999 0 0.00161306 3.3 0.00161298 3.3 0.00161308 0 0.0016129999999999999 0 0.0016131 3.3 0.00161302 3.3 0.00161312 0 0.0016130399999999998 0 0.0016131399999999999 3.3 0.00161306 3.3 0.00161316 0 0.0016130799999999998 0 0.0016131799999999999 3.3 0.0016131 3.3 0.0016132 0 0.00161312 0 0.00161322 3.3 0.0016131399999999999 3.3 0.00161324 0 0.00161316 0 0.00161326 3.3 0.0016131799999999999 3.3 0.00161328 0 0.0016132 0 0.0016133 3.3 0.0016132199999999998 3.3 0.00161332 0 0.00161324 0 0.00161334 3.3 0.0016132599999999998 3.3 0.0016133599999999999 0 0.00161328 0 0.00161338 3.3 0.0016132999999999998 3.3 0.0016133999999999999 0 0.00161332 0 0.00161342 3.3 0.00161334 3.3 0.00161344 0 0.0016133599999999999 0 0.00161346 3.3 0.00161338 3.3 0.00161348 0 0.0016133999999999999 0 0.0016135 3.3 0.00161342 3.3 0.00161352 0 0.0016134399999999998 0 0.00161354 3.3 0.00161346 3.3 0.00161356 0 0.0016134799999999998 0 0.0016135799999999999 3.3 0.0016135 3.3 0.0016136 0 0.00161352 0 0.00161362 3.3 0.00161354 3.3 0.00161364 0 0.00161356 0 0.00161366 3.3 0.0016135799999999999 3.3 0.00161368 0 0.0016136 0 0.0016137 3.3 0.0016136199999999999 3.3 0.00161372 0 0.00161364 0 0.00161374 3.3 0.0016136599999999998 3.3 0.0016137599999999999 0 0.00161368 0 0.00161378 3.3 0.0016136999999999998 3.3 0.0016137999999999999 0 0.00161372 0 0.00161382 3.3 0.00161374 3.3 0.00161384 0 0.0016137599999999999 0 0.00161386 3.3 0.00161378 3.3 0.00161388 0 0.0016137999999999999 0 0.0016139 3.3 0.00161382 3.3 0.00161392 0 0.0016138399999999998 0 0.00161394 3.3 0.00161386 3.3 0.00161396 0 0.0016138799999999998 0 0.0016139799999999999 3.3 0.0016139 3.3 0.001614 0 0.0016139199999999998 0 0.0016140199999999999 3.3 0.00161394 3.3 0.00161404 0 0.00161396 0 0.00161406 3.3 0.0016139799999999999 3.3 0.00161408 0 0.001614 0 0.0016141 3.3 0.0016140199999999999 3.3 0.00161412 0 0.00161404 0 0.00161414 3.3 0.0016140599999999998 3.3 0.00161416 0 0.00161408 0 0.00161418 3.3 0.0016140999999999998 3.3 0.0016141999999999999 0 0.00161412 0 0.00161422 3.3 0.00161414 3.3 0.00161424 0 0.00161416 0 0.00161426 3.3 0.00161418 3.3 0.00161428 0 0.0016141999999999999 0 0.0016143 3.3 0.00161422 3.3 0.00161432 0 0.0016142399999999999 0 0.00161434 3.3 0.00161426 3.3 0.00161436 0 0.0016142799999999998 0 0.00161438 3.3 0.0016143 3.3 0.0016144 0 0.0016143199999999998 0 0.0016144199999999999 3.3 0.00161434 3.3 0.00161444 0 0.00161436 0 0.00161446 3.3 0.00161438 3.3 0.00161448 0 0.0016144 0 0.0016145 3.3 0.0016144199999999999 3.3 0.00161452 0 0.00161444 0 0.00161454 3.3 0.0016144599999999999 3.3 0.00161456 0 0.00161448 0 0.00161458 3.3 0.0016144999999999998 3.3 0.0016145999999999999 0 0.00161452 0 0.00161462 3.3 0.0016145399999999998 3.3 0.0016146399999999999 0 0.00161456 0 0.00161466 3.3 0.00161458 3.3 0.00161468 0 0.0016145999999999999 0 0.0016147 3.3 0.00161462 3.3 0.00161472 0 0.0016146399999999999 0 0.00161474 3.3 0.00161466 3.3 0.00161476 0 0.0016146799999999998 0 0.00161478 3.3 0.0016147 3.3 0.0016148 0 0.0016147199999999998 0 0.0016148199999999999 3.3 0.00161474 3.3 0.00161484 0 0.0016147599999999998 0 0.0016148599999999999 3.3 0.00161478 3.3 0.00161488 0 0.0016148 0 0.0016149 3.3 0.0016148199999999999 3.3 0.00161492 0 0.00161484 0 0.00161494 3.3 0.0016148599999999999 3.3 0.00161496 0 0.00161488 0 0.00161498 3.3 0.0016148999999999998 3.3 0.001615 0 0.00161492 0 0.00161502 3.3 0.0016149399999999998 3.3 0.0016150399999999999 0 0.00161496 0 0.00161506 3.3 0.00161498 3.3 0.00161508 0 0.001615 0 0.0016151 3.3 0.00161502 3.3 0.00161512 0 0.0016150399999999999 0 0.00161514 3.3 0.00161506 3.3 0.00161516 0 0.0016150799999999999 0 0.00161518 3.3 0.0016151 3.3 0.0016152 0 0.0016151199999999998 0 0.00161522 3.3 0.00161514 3.3 0.00161524 0 0.0016151599999999998 0 0.0016152599999999999 3.3 0.00161518 3.3 0.00161528 0 0.0016152 0 0.0016153 3.3 0.00161522 3.3 0.00161532 0 0.00161524 0 0.00161534 3.3 0.0016152599999999999 3.3 0.00161536 0 0.00161528 0 0.00161538 3.3 0.0016152999999999999 3.3 0.0016154 0 0.00161532 0 0.00161542 3.3 0.0016153399999999998 3.3 0.0016154399999999999 0 0.00161536 0 0.00161546 3.3 0.0016153799999999998 3.3 0.0016154799999999999 0 0.0016154 0 0.0016155 3.3 0.00161542 3.3 0.00161552 0 0.0016154399999999999 0 0.00161554 3.3 0.00161546 3.3 0.00161556 0 0.0016154799999999999 0 0.00161558 3.3 0.0016155 3.3 0.0016156 0 0.0016155199999999998 0 0.00161562 3.3 0.00161554 3.3 0.00161564 0 0.0016155599999999998 0 0.0016156599999999999 3.3 0.00161558 3.3 0.00161568 0 0.0016155999999999998 0 0.0016156999999999999 3.3 0.00161562 3.3 0.00161572 0 0.00161564 0 0.00161574 3.3 0.0016156599999999999 3.3 0.00161576 0 0.00161568 0 0.00161578 3.3 0.0016156999999999999 3.3 0.0016158 0 0.00161572 0 0.00161582 3.3 0.0016157399999999998 3.3 0.00161584 0 0.00161576 0 0.00161586 3.3 0.0016157799999999998 3.3 0.0016158799999999999 0 0.0016158 0 0.0016159 3.3 0.00161582 3.3 0.00161592 0 0.00161584 0 0.00161594 3.3 0.00161586 3.3 0.00161596 0 0.0016158799999999999 0 0.00161598 3.3 0.0016159 3.3 0.001616 0 0.0016159199999999999 0 0.00161602 3.3 0.00161594 3.3 0.00161604 0 0.0016159599999999998 0 0.00161606 3.3 0.00161598 3.3 0.00161608 0 0.0016159999999999998 0 0.0016160999999999999 3.3 0.00161602 3.3 0.00161612 0 0.00161604 0 0.00161614 3.3 0.00161606 3.3 0.00161616 0 0.00161608 0 0.00161618 3.3 0.0016160999999999999 3.3 0.0016162 0 0.00161612 0 0.00161622 3.3 0.0016161399999999999 3.3 0.00161624 0 0.00161616 0 0.00161626 3.3 0.0016161799999999998 3.3 0.0016162799999999999 0 0.0016162 0 0.0016163 3.3 0.0016162199999999998 3.3 0.0016163199999999999 0 0.00161624 0 0.00161634 3.3 0.00161626 3.3 0.00161636 0 0.0016162799999999999 0 0.00161638 3.3 0.0016163 3.3 0.0016164 0 0.0016163199999999999 0 0.00161642 3.3 0.00161634 3.3 0.00161644 0 0.0016163599999999998 0 0.00161646 3.3 0.00161638 3.3 0.00161648 0 0.0016163999999999998 0 0.0016164999999999999 3.3 0.00161642 3.3 0.00161652 0 0.0016164399999999998 0 0.0016165399999999999 3.3 0.00161646 3.3 0.00161656 0 0.00161648 0 0.00161658 3.3 0.0016164999999999999 3.3 0.0016166 0 0.00161652 0 0.00161662 3.3 0.0016165399999999999 3.3 0.00161664 0 0.00161656 0 0.00161666 3.3 0.0016165799999999998 3.3 0.00161668 0 0.0016166 0 0.0016167 3.3 0.0016166199999999998 3.3 0.0016167199999999999 0 0.00161664 0 0.00161674 3.3 0.00161666 3.3 0.00161676 0 0.00161668 0 0.00161678 3.3 0.0016167 3.3 0.0016168 0 0.0016167199999999999 0 0.00161682 3.3 0.00161674 3.3 0.00161684 0 0.0016167599999999999 0 0.00161686 3.3 0.00161678 3.3 0.00161688 0 0.0016167999999999998 0 0.0016168999999999999 3.3 0.00161682 3.3 0.00161692 0 0.0016168399999999998 0 0.0016169399999999999 3.3 0.00161686 3.3 0.00161696 0 0.00161688 0 0.00161698 3.3 0.0016168999999999999 3.3 0.001617 0 0.00161692 0 0.00161702 3.3 0.0016169399999999999 3.3 0.00161704 0 0.00161696 0 0.00161706 3.3 0.0016169799999999998 3.3 0.00161708 0 0.001617 0 0.0016171 3.3 0.0016170199999999998 3.3 0.0016171199999999999 0 0.00161704 0 0.00161714 3.3 0.0016170599999999998 3.3 0.0016171599999999999 0 0.00161708 0 0.00161718 3.3 0.0016171 3.3 0.0016172 0 0.0016171199999999999 0 0.00161722 3.3 0.00161714 3.3 0.00161724 0 0.0016171599999999999 0 0.00161726 3.3 0.00161718 3.3 0.00161728 0 0.0016171999999999998 0 0.0016173 3.3 0.00161722 3.3 0.00161732 0 0.0016172399999999998 0 0.0016173399999999999 3.3 0.00161726 3.3 0.00161736 0 0.0016172799999999998 0 0.0016173799999999999 3.3 0.0016173 3.3 0.0016174 0 0.00161732 0 0.00161742 3.3 0.0016173399999999999 3.3 0.00161744 0 0.00161736 0 0.00161746 3.3 0.0016173799999999999 3.3 0.00161748 0 0.0016174 0 0.0016175 3.3 0.0016174199999999998 3.3 0.00161752 0 0.00161744 0 0.00161754 3.3 0.0016174599999999998 3.3 0.0016175599999999999 0 0.00161748 0 0.00161758 3.3 0.0016175 3.3 0.0016176 0 0.00161752 0 0.00161762 3.3 0.00161754 3.3 0.00161764 0 0.0016175599999999999 0 0.00161766 3.3 0.00161758 3.3 0.00161768 0 0.0016175999999999999 0 0.0016177 3.3 0.00161762 3.3 0.00161772 0 0.0016176399999999998 0 0.0016177399999999999 3.3 0.00161766 3.3 0.00161776 0 0.0016176799999999998 0 0.0016177799999999999 3.3 0.0016177 3.3 0.0016178 0 0.00161772 0 0.00161782 3.3 0.0016177399999999999 3.3 0.00161784 0 0.00161776 0 0.00161786 3.3 0.0016177799999999999 3.3 0.00161788 0 0.0016178 0 0.0016179 3.3 0.0016178199999999998 3.3 0.00161792 0 0.00161784 0 0.00161794 3.3 0.0016178599999999998 3.3 0.0016179599999999999 0 0.00161788 0 0.00161798 3.3 0.0016178999999999998 3.3 0.0016179999999999999 0 0.00161792 0 0.00161802 3.3 0.00161794 3.3 0.00161804 0 0.0016179599999999999 0 0.00161806 3.3 0.00161798 3.3 0.00161808 0 0.0016179999999999999 0 0.0016181 3.3 0.00161802 3.3 0.00161812 0 0.0016180399999999998 0 0.00161814 3.3 0.00161806 3.3 0.00161816 0 0.0016180799999999998 0 0.0016181799999999999 3.3 0.0016181 3.3 0.0016182 0 0.00161812 0 0.00161822 3.3 0.00161814 3.3 0.00161824 0 0.00161816 0 0.00161826 3.3 0.0016181799999999999 3.3 0.00161828 0 0.0016182 0 0.0016183 3.3 0.0016182199999999999 3.3 0.00161832 0 0.00161824 0 0.00161834 3.3 0.0016182599999999998 3.3 0.00161836 0 0.00161828 0 0.00161838 3.3 0.0016182999999999998 3.3 0.0016183999999999999 0 0.00161832 0 0.00161842 3.3 0.00161834 3.3 0.00161844 0 0.00161836 0 0.00161846 3.3 0.00161838 3.3 0.00161848 0 0.0016183999999999999 0 0.0016185 3.3 0.00161842 3.3 0.00161852 0 0.0016184399999999999 0 0.00161854 3.3 0.00161846 3.3 0.00161856 0 0.0016184799999999998 0 0.0016185799999999999 3.3 0.0016185 3.3 0.0016186 0 0.0016185199999999998 0 0.0016186199999999999 3.3 0.00161854 3.3 0.00161864 0 0.00161856 0 0.00161866 3.3 0.0016185799999999999 3.3 0.00161868 0 0.0016186 0 0.0016187 3.3 0.0016186199999999999 3.3 0.00161872 0 0.00161864 0 0.00161874 3.3 0.0016186599999999998 3.3 0.00161876 0 0.00161868 0 0.00161878 3.3 0.0016186999999999998 3.3 0.0016187999999999999 0 0.00161872 0 0.00161882 3.3 0.0016187399999999998 3.3 0.0016188399999999999 0 0.00161876 0 0.00161886 3.3 0.00161878 3.3 0.00161888 0 0.0016187999999999999 0 0.0016189 3.3 0.00161882 3.3 0.00161892 0 0.0016188399999999999 0 0.00161894 3.3 0.00161886 3.3 0.00161896 0 0.0016188799999999998 0 0.00161898 3.3 0.0016189 3.3 0.001619 0 0.0016189199999999998 0 0.0016190199999999999 3.3 0.00161894 3.3 0.00161904 0 0.00161896 0 0.00161906 3.3 0.00161898 3.3 0.00161908 0 0.001619 0 0.0016191 3.3 0.0016190199999999999 3.3 0.00161912 0 0.00161904 0 0.00161914 3.3 0.0016190599999999999 3.3 0.00161916 0 0.00161908 0 0.00161918 3.3 0.0016190999999999998 3.3 0.0016192 0 0.00161912 0 0.00161922 3.3 0.0016191399999999998 3.3 0.0016192399999999999 0 0.00161916 0 0.00161926 3.3 0.00161918 3.3 0.00161928 0 0.0016192 0 0.0016193 3.3 0.00161922 3.3 0.00161932 0 0.0016192399999999999 0 0.00161934 3.3 0.00161926 3.3 0.00161936 0 0.0016192799999999999 0 0.00161938 3.3 0.0016193 3.3 0.0016194 0 0.0016193199999999998 0 0.0016194199999999999 3.3 0.00161934 3.3 0.00161944 0 0.0016193599999999998 0 0.0016194599999999999 3.3 0.00161938 3.3 0.00161948 0 0.0016194 0 0.0016195 3.3 0.0016194199999999999 3.3 0.00161952 0 0.00161944 0 0.00161954 3.3 0.0016194599999999999 3.3 0.00161956 0 0.00161948 0 0.00161958 3.3 0.0016194999999999998 3.3 0.0016196 0 0.00161952 0 0.00161962 3.3 0.0016195399999999998 3.3 0.0016196399999999999 0 0.00161956 0 0.00161966 3.3 0.0016195799999999998 3.3 0.0016196799999999999 0 0.0016196 0 0.0016197 3.3 0.00161962 3.3 0.00161972 0 0.0016196399999999999 0 0.00161974 3.3 0.00161966 3.3 0.00161976 0 0.0016196799999999999 0 0.00161978 3.3 0.0016197 3.3 0.0016198 0 0.0016197199999999998 0 0.00161982 3.3 0.00161974 3.3 0.00161984 0 0.0016197599999999998 0 0.0016198599999999999 3.3 0.00161978 3.3 0.00161988 0 0.0016198 0 0.0016199 3.3 0.00161982 3.3 0.00161992 0 0.00161984 0 0.00161994 3.3 0.0016198599999999999 3.3 0.00161996 0 0.00161988 0 0.00161998 3.3 0.0016198999999999999 3.3 0.00162 0 0.00161992 0 0.00162002 3.3 0.0016199399999999998 3.3 0.00162004 0 0.00161996 0 0.00162006 3.3 0.0016199799999999998 3.3 0.0016200799999999999 0 0.00162 0 0.0016201 3.3 0.00162002 3.3 0.00162012 0 0.00162004 0 0.00162014 3.3 0.00162006 3.3 0.00162016 0 0.0016200799999999999 0 0.00162018 3.3 0.0016201 3.3 0.0016202 0 0.0016201199999999999 0 0.00162022 3.3 0.00162014 3.3 0.00162024 0 0.0016201599999999998 0 0.0016202599999999999 3.3 0.00162018 3.3 0.00162028 0 0.0016201999999999998 0 0.0016202999999999999 3.3 0.00162022 3.3 0.00162032 0 0.00162024 0 0.00162034 3.3 0.0016202599999999999 3.3 0.00162036 0 0.00162028 0 0.00162038 3.3 0.0016202999999999999 3.3 0.0016204 0 0.00162032 0 0.00162042 3.3 0.0016203399999999998 3.3 0.00162044 0 0.00162036 0 0.00162046 3.3 0.0016203799999999998 3.3 0.0016204799999999999 0 0.0016204 0 0.0016205 3.3 0.0016204199999999998 3.3 0.0016205199999999999 0 0.00162044 0 0.00162054 3.3 0.00162046 3.3 0.00162056 0 0.0016204799999999999 0 0.00162058 3.3 0.0016205 3.3 0.0016206 0 0.0016205199999999999 0 0.00162062 3.3 0.00162054 3.3 0.00162064 0 0.0016205599999999998 0 0.00162066 3.3 0.00162058 3.3 0.00162068 0 0.0016205999999999998 0 0.0016206999999999999 3.3 0.00162062 3.3 0.00162072 0 0.00162064 0 0.00162074 3.3 0.00162066 3.3 0.00162076 0 0.00162068 0 0.00162078 3.3 0.0016206999999999999 3.3 0.0016208 0 0.00162072 0 0.00162082 3.3 0.0016207399999999999 3.3 0.00162084 0 0.00162076 0 0.00162086 3.3 0.0016207799999999998 3.3 0.0016208799999999999 0 0.0016208 0 0.0016209 3.3 0.0016208199999999998 3.3 0.0016209199999999999 0 0.00162084 0 0.00162094 3.3 0.00162086 3.3 0.00162096 0 0.0016208799999999999 0 0.00162098 3.3 0.0016209 3.3 0.001621 0 0.0016209199999999999 0 0.00162102 3.3 0.00162094 3.3 0.00162104 0 0.0016209599999999998 0 0.00162106 3.3 0.00162098 3.3 0.00162108 0 0.0016209999999999998 0 0.0016210999999999999 3.3 0.00162102 3.3 0.00162112 0 0.0016210399999999998 0 0.0016211399999999999 3.3 0.00162106 3.3 0.00162116 0 0.00162108 0 0.00162118 3.3 0.0016210999999999999 3.3 0.0016212 0 0.00162112 0 0.00162122 3.3 0.0016211399999999999 3.3 0.00162124 0 0.00162116 0 0.00162126 3.3 0.0016211799999999998 3.3 0.00162128 0 0.0016212 0 0.0016213 3.3 0.0016212199999999998 3.3 0.0016213199999999999 0 0.00162124 0 0.00162134 3.3 0.00162126 3.3 0.00162136 0 0.00162128 0 0.00162138 3.3 0.0016213 3.3 0.0016214 0 0.0016213199999999999 0 0.00162142 3.3 0.00162134 3.3 0.00162144 0 0.0016213599999999999 0 0.00162146 3.3 0.00162138 3.3 0.00162148 0 0.0016213999999999998 0 0.0016215 3.3 0.00162142 3.3 0.00162152 0 0.0016214399999999998 0 0.0016215399999999999 3.3 0.00162146 3.3 0.00162156 0 0.00162148 0 0.00162158 3.3 0.0016215 3.3 0.0016216 0 0.00162152 0 0.00162162 3.3 0.0016215399999999999 3.3 0.00162164 0 0.00162156 0 0.00162166 3.3 0.0016215799999999999 3.3 0.00162168 0 0.0016216 0 0.0016217 3.3 0.0016216199999999998 3.3 0.0016217199999999999 0 0.00162164 0 0.00162174 3.3 0.0016216599999999998 3.3 0.0016217599999999999 0 0.00162168 0 0.00162178 3.3 0.0016217 3.3 0.0016218 0 0.0016217199999999999 0 0.00162182 3.3 0.00162174 3.3 0.00162184 0 0.0016217599999999999 0 0.00162186 3.3 0.00162178 3.3 0.00162188 0 0.0016217999999999998 0 0.0016219 3.3 0.00162182 3.3 0.00162192 0 0.0016218399999999998 0 0.0016219399999999999 3.3 0.00162186 3.3 0.00162196 0 0.0016218799999999998 0 0.0016219799999999999 3.3 0.0016219 3.3 0.001622 0 0.00162192 0 0.00162202 3.3 0.0016219399999999999 3.3 0.00162204 0 0.00162196 0 0.00162206 3.3 0.0016219799999999999 3.3 0.00162208 0 0.001622 0 0.0016221 3.3 0.0016220199999999998 3.3 0.00162212 0 0.00162204 0 0.00162214 3.3 0.0016220599999999998 3.3 0.0016221599999999999 0 0.00162208 0 0.00162218 3.3 0.0016221 3.3 0.0016222 0 0.00162212 0 0.00162222 3.3 0.00162214 3.3 0.00162224 0 0.0016221599999999999 0 0.00162226 3.3 0.00162218 3.3 0.00162228 0 0.0016221999999999999 0 0.0016223 3.3 0.00162222 3.3 0.00162232 0 0.0016222399999999998 0 0.00162234 3.3 0.00162226 3.3 0.00162236 0 0.0016222799999999998 0 0.0016223799999999999 3.3 0.0016223 3.3 0.0016224 0 0.00162232 0 0.00162242 3.3 0.00162234 3.3 0.00162244 0 0.00162236 0 0.00162246 3.3 0.0016223799999999999 3.3 0.00162248 0 0.0016224 0 0.0016225 3.3 0.0016224199999999999 3.3 0.00162252 0 0.00162244 0 0.00162254 3.3 0.0016224599999999998 3.3 0.0016225599999999999 0 0.00162248 0 0.00162258 3.3 0.0016224999999999998 3.3 0.0016225999999999999 0 0.00162252 0 0.00162262 3.3 0.00162254 3.3 0.00162264 0 0.0016225599999999999 0 0.00162266 3.3 0.00162258 3.3 0.00162268 0 0.0016225999999999999 0 0.0016227 3.3 0.00162262 3.3 0.00162272 0 0.0016226399999999998 0 0.00162274 3.3 0.00162266 3.3 0.00162276 0 0.0016226799999999998 0 0.0016227799999999999 3.3 0.0016227 3.3 0.0016228 0 0.0016227199999999998 0 0.0016228199999999999 3.3 0.00162274 3.3 0.00162284 0 0.00162276 0 0.00162286 3.3 0.0016227799999999999 3.3 0.00162288 0 0.0016228 0 0.0016229 3.3 0.0016228199999999999 3.3 0.00162292 0 0.00162284 0 0.00162294 3.3 0.0016228599999999998 3.3 0.00162296 0 0.00162288 0 0.00162298 3.3 0.0016228999999999998 3.3 0.0016229999999999999 0 0.00162292 0 0.00162302 3.3 0.00162294 3.3 0.00162304 0 0.00162296 0 0.00162306 3.3 0.00162298 3.3 0.00162308 0 0.0016229999999999999 0 0.0016231 3.3 0.00162302 3.3 0.00162312 0 0.0016230399999999999 0 0.00162314 3.3 0.00162306 3.3 0.00162316 0 0.0016230799999999998 0 0.00162318 3.3 0.0016231 3.3 0.0016232 0 0.0016231199999999998 0 0.0016232199999999999 3.3 0.00162314 3.3 0.00162324 0 0.00162316 0 0.00162326 3.3 0.00162318 3.3 0.00162328 0 0.0016232 0 0.0016233 3.3 0.0016232199999999999 3.3 0.00162332 0 0.00162324 0 0.00162334 3.3 0.0016232599999999999 3.3 0.00162336 0 0.00162328 0 0.00162338 3.3 0.0016232999999999998 3.3 0.0016233999999999999 0 0.00162332 0 0.00162342 3.3 0.0016233399999999998 3.3 0.0016234399999999999 0 0.00162336 0 0.00162346 3.3 0.00162338 3.3 0.00162348 0 0.0016233999999999999 0 0.0016235 3.3 0.00162342 3.3 0.00162352 0 0.0016234399999999999 0 0.00162354 3.3 0.00162346 3.3 0.00162356 0 0.0016234799999999998 0 0.00162358 3.3 0.0016235 3.3 0.0016236 0 0.0016235199999999998 0 0.0016236199999999999 3.3 0.00162354 3.3 0.00162364 0 0.0016235599999999998 0 0.0016236599999999999 3.3 0.00162358 3.3 0.00162368 0 0.0016236 0 0.0016237 3.3 0.0016236199999999999 3.3 0.00162372 0 0.00162364 0 0.00162374 3.3 0.0016236599999999999 3.3 0.00162376 0 0.00162368 0 0.00162378 3.3 0.0016236999999999998 3.3 0.0016238 0 0.00162372 0 0.00162382 3.3 0.0016237399999999998 3.3 0.0016238399999999999 0 0.00162376 0 0.00162386 3.3 0.00162378 3.3 0.00162388 0 0.0016238 0 0.0016239 3.3 0.00162382 3.3 0.00162392 0 0.0016238399999999999 0 0.00162394 3.3 0.00162386 3.3 0.00162396 0 0.0016238799999999999 0 0.00162398 3.3 0.0016239 3.3 0.001624 0 0.0016239199999999998 0 0.0016240199999999999 3.3 0.00162394 3.3 0.00162404 0 0.0016239599999999998 0 0.0016240599999999999 3.3 0.00162398 3.3 0.00162408 0 0.001624 0 0.0016241 3.3 0.0016240199999999999 3.3 0.00162412 0 0.00162404 0 0.00162414 3.3 0.0016240599999999999 3.3 0.00162416 0 0.00162408 0 0.00162418 3.3 0.0016240999999999998 3.3 0.0016242 0 0.00162412 0 0.00162422 3.3 0.0016241399999999998 3.3 0.0016242399999999999 0 0.00162416 0 0.00162426 3.3 0.0016241799999999998 3.3 0.0016242799999999999 0 0.0016242 0 0.0016243 3.3 0.00162422 3.3 0.00162432 0 0.0016242399999999999 0 0.00162434 3.3 0.00162426 3.3 0.00162436 0 0.0016242799999999999 0 0.00162438 3.3 0.0016243 3.3 0.0016244 0 0.0016243199999999998 0 0.00162442 3.3 0.00162434 3.3 0.00162444 0 0.0016243599999999998 0 0.0016244599999999999 3.3 0.00162438 3.3 0.00162448 0 0.0016243999999999998 0 0.0016244999999999999 3.3 0.00162442 3.3 0.00162452 0 0.00162444 0 0.00162454 3.3 0.0016244599999999999 3.3 0.00162456 0 0.00162448 0 0.00162458 3.3 0.0016244999999999999 3.3 0.0016246 0 0.00162452 0 0.00162462 3.3 0.0016245399999999998 3.3 0.00162464 0 0.00162456 0 0.00162466 3.3 0.0016245799999999998 3.3 0.0016246799999999999 0 0.0016246 0 0.0016247 3.3 0.00162462 3.3 0.00162472 0 0.00162464 0 0.00162474 3.3 0.00162466 3.3 0.00162476 0 0.0016246799999999999 0 0.00162478 3.3 0.0016247 3.3 0.0016248 0 0.0016247199999999999 0 0.00162482 3.3 0.00162474 3.3 0.00162484 0 0.0016247599999999998 0 0.0016248599999999999 3.3 0.00162478 3.3 0.00162488 0 0.0016247999999999998 0 0.0016248999999999999 3.3 0.00162482 3.3 0.00162492 0 0.00162484 0 0.00162494 3.3 0.0016248599999999999 3.3 0.00162496 0 0.00162488 0 0.00162498 3.3 0.0016248999999999999 3.3 0.001625 0 0.00162492 0 0.00162502 3.3 0.0016249399999999998 3.3 0.00162504 0 0.00162496 0 0.00162506 3.3 0.0016249799999999998 3.3 0.0016250799999999999 0 0.001625 0 0.0016251 3.3 0.0016250199999999998 3.3 0.0016251199999999999 0 0.00162504 0 0.00162514 3.3 0.00162506 3.3 0.00162516 0 0.0016250799999999999 0 0.00162518 3.3 0.0016251 3.3 0.0016252 0 0.0016251199999999999 0 0.00162522 3.3 0.00162514 3.3 0.00162524 0 0.0016251599999999998 0 0.00162526 3.3 0.00162518 3.3 0.00162528 0 0.0016251999999999998 0 0.0016252999999999999 3.3 0.00162522 3.3 0.00162532 0 0.00162524 0 0.00162534 3.3 0.00162526 3.3 0.00162536 0 0.00162528 0 0.00162538 3.3 0.0016252999999999999 3.3 0.0016254 0 0.00162532 0 0.00162542 3.3 0.0016253399999999999 3.3 0.00162544 0 0.00162536 0 0.00162546 3.3 0.0016253799999999998 3.3 0.00162548 0 0.0016254 0 0.0016255 3.3 0.0016254199999999998 3.3 0.0016255199999999999 0 0.00162544 0 0.00162554 3.3 0.00162546 3.3 0.00162556 0 0.00162548 0 0.00162558 3.3 0.0016255 3.3 0.0016256 0 0.0016255199999999999 0 0.00162562 3.3 0.00162554 3.3 0.00162564 0 0.0016255599999999999 0 0.00162566 3.3 0.00162558 3.3 0.00162568 0 0.0016255999999999998 0 0.0016256999999999999 3.3 0.00162562 3.3 0.00162572 0 0.0016256399999999998 0 0.0016257399999999999 3.3 0.00162566 3.3 0.00162576 0 0.00162568 0 0.00162578 3.3 0.0016256999999999999 3.3 0.0016258 0 0.00162572 0 0.00162582 3.3 0.0016257399999999999 3.3 0.00162584 0 0.00162576 0 0.00162586 3.3 0.0016257799999999998 3.3 0.00162588 0 0.0016258 0 0.0016259 3.3 0.0016258199999999998 3.3 0.0016259199999999999 0 0.00162584 0 0.00162594 3.3 0.0016258599999999998 3.3 0.0016259599999999999 0 0.00162588 0 0.00162598 3.3 0.0016259 3.3 0.001626 0 0.0016259199999999999 0 0.00162602 3.3 0.00162594 3.3 0.00162604 0 0.0016259599999999999 0 0.00162606 3.3 0.00162598 3.3 0.00162608 0 0.0016259999999999998 0 0.0016261 3.3 0.00162602 3.3 0.00162612 0 0.0016260399999999998 0 0.0016261399999999999 3.3 0.00162606 3.3 0.00162616 0 0.00162608 0 0.00162618 3.3 0.0016261 3.3 0.0016262 0 0.00162612 0 0.00162622 3.3 0.0016261399999999999 3.3 0.00162624 0 0.00162616 0 0.00162626 3.3 0.0016261799999999999 3.3 0.00162628 0 0.0016262 0 0.0016263 3.3 0.0016262199999999998 3.3 0.00162632 0 0.00162624 0 0.00162634 3.3 0.0016262599999999998 3.3 0.0016263599999999999 0 0.00162628 0 0.00162638 3.3 0.0016263 3.3 0.0016264 0 0.00162632 0 0.00162642 3.3 0.00162634 3.3 0.00162644 0 0.0016263599999999999 0 0.00162646 3.3 0.00162638 3.3 0.00162648 0 0.0016263999999999999 0 0.0016265 3.3 0.00162642 3.3 0.00162652 0 0.0016264399999999998 0 0.0016265399999999999 3.3 0.00162646 3.3 0.00162656 0 0.0016264799999999998 0 0.0016265799999999999 3.3 0.0016265 3.3 0.0016266 0 0.00162652 0 0.00162662 3.3 0.0016265399999999999 3.3 0.00162664 0 0.00162656 0 0.00162666 3.3 0.0016265799999999999 3.3 0.00162668 0 0.0016266 0 0.0016267 3.3 0.0016266199999999998 3.3 0.00162672 0 0.00162664 0 0.00162674 3.3 0.0016266599999999998 3.3 0.0016267599999999999 0 0.00162668 0 0.00162678 3.3 0.0016266999999999998 3.3 0.0016267999999999999 0 0.00162672 0 0.00162682 3.3 0.00162674 3.3 0.00162684 0 0.0016267599999999999 0 0.00162686 3.3 0.00162678 3.3 0.00162688 0 0.0016267999999999999 0 0.0016269 3.3 0.00162682 3.3 0.00162692 0 0.0016268399999999998 0 0.00162694 3.3 0.00162686 3.3 0.00162696 0 0.0016268799999999998 0 0.0016269799999999999 3.3 0.0016269 3.3 0.001627 0 0.00162692 0 0.00162702 3.3 0.00162694 3.3 0.00162704 0 0.00162696 0 0.00162706 3.3 0.0016269799999999999 3.3 0.00162708 0 0.001627 0 0.0016271 3.3 0.0016270199999999999 3.3 0.00162712 0 0.00162704 0 0.00162714 3.3 0.0016270599999999998 3.3 0.0016271599999999999 0 0.00162708 0 0.00162718 3.3 0.0016270999999999998 3.3 0.0016271999999999999 0 0.00162712 0 0.00162722 3.3 0.00162714 3.3 0.00162724 0 0.0016271599999999999 0 0.00162726 3.3 0.00162718 3.3 0.00162728 0 0.0016271999999999999 0 0.0016273 3.3 0.00162722 3.3 0.00162732 0 0.0016272399999999998 0 0.00162734 3.3 0.00162726 3.3 0.00162736 0 0.0016272799999999998 0 0.0016273799999999999 3.3 0.0016273 3.3 0.0016274 0 0.0016273199999999998 0 0.0016274199999999999 3.3 0.00162734 3.3 0.00162744 0 0.00162736 0 0.00162746 3.3 0.0016273799999999999 3.3 0.00162748 0 0.0016274 0 0.0016275 3.3 0.0016274199999999999 3.3 0.00162752 0 0.00162744 0 0.00162754 3.3 0.0016274599999999998 3.3 0.00162756 0 0.00162748 0 0.00162758 3.3 0.0016274999999999998 3.3 0.0016275999999999999 0 0.00162752 0 0.00162762 3.3 0.0016275399999999998 3.3 0.0016276399999999999 0 0.00162756 0 0.00162766 3.3 0.00162758 3.3 0.00162768 0 0.0016275999999999999 0 0.0016277 3.3 0.00162762 3.3 0.00162772 0 0.0016276399999999999 0 0.00162774 3.3 0.00162766 3.3 0.00162776 0 0.0016276799999999998 0 0.00162778 3.3 0.0016277 3.3 0.0016278 0 0.0016277199999999998 0 0.0016278199999999999 3.3 0.00162774 3.3 0.00162784 0 0.00162776 0 0.00162786 3.3 0.00162778 3.3 0.00162788 0 0.0016278 0 0.0016279 3.3 0.0016278199999999999 3.3 0.00162792 0 0.00162784 0 0.00162794 3.3 0.0016278599999999999 3.3 0.00162796 0 0.00162788 0 0.00162798 3.3 0.0016278999999999998 3.3 0.0016279999999999999 0 0.00162792 0 0.00162802 3.3 0.0016279399999999998 3.3 0.0016280399999999999 0 0.00162796 0 0.00162806 3.3 0.00162798 3.3 0.00162808 0 0.0016279999999999999 0 0.0016281 3.3 0.00162802 3.3 0.00162812 0 0.0016280399999999999 0 0.00162814 3.3 0.00162806 3.3 0.00162816 0 0.0016280799999999998 0 0.00162818 3.3 0.0016281 3.3 0.0016282 0 0.0016281199999999998 0 0.0016282199999999999 3.3 0.00162814 3.3 0.00162824 0 0.0016281599999999998 0 0.0016282599999999999 3.3 0.00162818 3.3 0.00162828 0 0.0016282 0 0.0016283 3.3 0.0016282199999999999 3.3 0.00162832 0 0.00162824 0 0.00162834 3.3 0.0016282599999999999 3.3 0.00162836 0 0.00162828 0 0.00162838 3.3 0.0016282999999999998 3.3 0.0016284 0 0.00162832 0 0.00162842 3.3 0.0016283399999999998 3.3 0.0016284399999999999 0 0.00162836 0 0.00162846 3.3 0.00162838 3.3 0.00162848 0 0.0016284 0 0.0016285 3.3 0.00162842 3.3 0.00162852 0 0.0016284399999999999 0 0.00162854 3.3 0.00162846 3.3 0.00162856 0 0.0016284799999999999 0 0.00162858 3.3 0.0016285 3.3 0.0016286 0 0.0016285199999999998 0 0.00162862 3.3 0.00162854 3.3 0.00162864 0 0.0016285599999999998 0 0.0016286599999999999 3.3 0.00162858 3.3 0.00162868 0 0.0016286 0 0.0016287 3.3 0.00162862 3.3 0.00162872 0 0.00162864 0 0.00162874 3.3 0.0016286599999999999 3.3 0.00162876 0 0.00162868 0 0.00162878 3.3 0.0016286999999999999 3.3 0.0016288 0 0.00162872 0 0.00162882 3.3 0.0016287399999999998 3.3 0.0016288399999999999 0 0.00162876 0 0.00162886 3.3 0.0016287799999999998 3.3 0.0016288799999999999 0 0.0016288 0 0.0016289 3.3 0.00162882 3.3 0.00162892 0 0.0016288399999999999 0 0.00162894 3.3 0.00162886 3.3 0.00162896 0 0.0016288799999999999 0 0.00162898 3.3 0.0016289 3.3 0.001629 0 0.0016289199999999998 0 0.00162902 3.3 0.00162894 3.3 0.00162904 0 0.0016289599999999998 0 0.0016290599999999999 3.3 0.00162898 3.3 0.00162908 0 0.0016289999999999998 0 0.0016290999999999999 3.3 0.00162902 3.3 0.00162912 0 0.00162904 0 0.00162914 3.3 0.0016290599999999999 3.3 0.00162916 0 0.00162908 0 0.00162918 3.3 0.0016290999999999999 3.3 0.0016292 0 0.00162912 0 0.00162922 3.3 0.0016291399999999998 3.3 0.00162924 0 0.00162916 0 0.00162926 3.3 0.0016291799999999998 3.3 0.0016292799999999999 0 0.0016292 0 0.0016293 3.3 0.00162922 3.3 0.00162932 0 0.00162924 0 0.00162934 3.3 0.00162926 3.3 0.00162936 0 0.0016292799999999999 0 0.00162938 3.3 0.0016293 3.3 0.0016294 0 0.0016293199999999999 0 0.00162942 3.3 0.00162934 3.3 0.00162944 0 0.0016293599999999998 0 0.00162946 3.3 0.00162938 3.3 0.00162948 0 0.0016293999999999998 0 0.0016294999999999999 3.3 0.00162942 3.3 0.00162952 0 0.00162944 0 0.00162954 3.3 0.00162946 3.3 0.00162956 0 0.00162948 0 0.00162958 3.3 0.0016294999999999999 3.3 0.0016296 0 0.00162952 0 0.00162962 3.3 0.0016295399999999999 3.3 0.00162964 0 0.00162956 0 0.00162966 3.3 0.0016295799999999998 3.3 0.0016296799999999999 0 0.0016296 0 0.0016297 3.3 0.0016296199999999998 3.3 0.0016297199999999999 0 0.00162964 0 0.00162974 3.3 0.00162966 3.3 0.00162976 0 0.0016296799999999999 0 0.00162978 3.3 0.0016297 3.3 0.0016298 0 0.0016297199999999999 0 0.00162982 3.3 0.00162974 3.3 0.00162984 0 0.0016297599999999998 0 0.00162986 3.3 0.00162978 3.3 0.00162988 0 0.0016297999999999998 0 0.0016298999999999999 3.3 0.00162982 3.3 0.00162992 0 0.0016298399999999998 0 0.0016299399999999999 3.3 0.00162986 3.3 0.00162996 0 0.00162988 0 0.00162998 3.3 0.0016298999999999999 3.3 0.00163 0 0.00162992 0 0.00163002 3.3 0.0016299399999999999 3.3 0.00163004 0 0.00162996 0 0.00163006 3.3 0.0016299799999999998 3.3 0.00163008 0 0.00163 0 0.0016301 3.3 0.0016300199999999998 3.3 0.0016301199999999999 0 0.00163004 0 0.00163014 3.3 0.00163006 3.3 0.00163016 0 0.00163008 0 0.00163018 3.3 0.0016301 3.3 0.0016302 0 0.0016301199999999999 0 0.00163022 3.3 0.00163014 3.3 0.00163024 0 0.0016301599999999999 0 0.00163026 3.3 0.00163018 3.3 0.00163028 0 0.0016301999999999998 0 0.0016303 3.3 0.00163022 3.3 0.00163032 0 0.0016302399999999998 0 0.0016303399999999999 3.3 0.00163026 3.3 0.00163036 0 0.00163028 0 0.00163038 3.3 0.0016303 3.3 0.0016304 0 0.00163032 0 0.00163042 3.3 0.0016303399999999999 3.3 0.00163044 0 0.00163036 0 0.00163046 3.3 0.0016303799999999999 3.3 0.00163048 0 0.0016304 0 0.0016305 3.3 0.0016304199999999998 3.3 0.0016305199999999999 0 0.00163044 0 0.00163054 3.3 0.0016304599999999998 3.3 0.0016305599999999999 0 0.00163048 0 0.00163058 3.3 0.0016305 3.3 0.0016306 0 0.0016305199999999999 0 0.00163062 3.3 0.00163054 3.3 0.00163064 0 0.0016305599999999999 0 0.00163066 3.3 0.00163058 3.3 0.00163068 0 0.0016305999999999998 0 0.0016307 3.3 0.00163062 3.3 0.00163072 0 0.0016306399999999998 0 0.0016307399999999999 3.3 0.00163066 3.3 0.00163076 0 0.0016306799999999998 0 0.0016307799999999999 3.3 0.0016307 3.3 0.0016308 0 0.00163072 0 0.00163082 3.3 0.0016307399999999999 3.3 0.00163084 0 0.00163076 0 0.00163086 3.3 0.0016307799999999999 3.3 0.00163088 0 0.0016308 0 0.0016309 3.3 0.0016308199999999998 3.3 0.00163092 0 0.00163084 0 0.00163094 3.3 0.0016308599999999998 3.3 0.0016309599999999999 0 0.00163088 0 0.00163098 3.3 0.0016309 3.3 0.001631 0 0.00163092 0 0.00163102 3.3 0.00163094 3.3 0.00163104 0 0.0016309599999999999 0 0.00163106 3.3 0.00163098 3.3 0.00163108 0 0.0016309999999999999 0 0.0016311 3.3 0.00163102 3.3 0.00163112 0 0.0016310399999999998 0 0.0016311399999999999 3.3 0.00163106 3.3 0.00163116 0 0.0016310799999999998 0 0.0016311799999999999 3.3 0.0016311 3.3 0.0016312 0 0.00163112 0 0.00163122 3.3 0.0016311399999999999 3.3 0.00163124 0 0.00163116 0 0.00163126 3.3 0.0016311799999999999 3.3 0.00163128 0 0.0016312 0 0.0016313 3.3 0.0016312199999999998 3.3 0.00163132 0 0.00163124 0 0.00163134 3.3 0.0016312599999999998 3.3 0.0016313599999999999 0 0.00163128 0 0.00163138 3.3 0.0016312999999999998 3.3 0.0016313999999999999 0 0.00163132 0 0.00163142 3.3 0.00163134 3.3 0.00163144 0 0.0016313599999999999 0 0.00163146 3.3 0.00163138 3.3 0.00163148 0 0.0016313999999999999 0 0.0016315 3.3 0.00163142 3.3 0.00163152 0 0.0016314399999999998 0 0.00163154 3.3 0.00163146 3.3 0.00163156 0 0.0016314799999999998 0 0.0016315799999999999 3.3 0.0016315 3.3 0.0016316 0 0.00163152 0 0.00163162 3.3 0.00163154 3.3 0.00163164 0 0.00163156 0 0.00163166 3.3 0.0016315799999999999 3.3 0.00163168 0 0.0016316 0 0.0016317 3.3 0.0016316199999999999 3.3 0.00163172 0 0.00163164 0 0.00163174 3.3 0.0016316599999999998 3.3 0.00163176 0 0.00163168 0 0.00163178 3.3 0.0016316999999999998 3.3 0.0016317999999999999 0 0.00163172 0 0.00163182 3.3 0.00163174 3.3 0.00163184 0 0.00163176 0 0.00163186 3.3 0.00163178 3.3 0.00163188 0 0.0016317999999999999 0 0.0016319 3.3 0.00163182 3.3 0.00163192 0 0.0016318399999999999 0 0.00163194 3.3 0.00163186 3.3 0.00163196 0 0.0016318799999999998 0 0.0016319799999999999 3.3 0.0016319 3.3 0.001632 0 0.0016319199999999998 0 0.0016320199999999999 3.3 0.00163194 3.3 0.00163204 0 0.00163196 0 0.00163206 3.3 0.0016319799999999999 3.3 0.00163208 0 0.001632 0 0.0016321 3.3 0.0016320199999999999 3.3 0.00163212 0 0.00163204 0 0.00163214 3.3 0.0016320599999999998 3.3 0.00163216 0 0.00163208 0 0.00163218 3.3 0.0016320999999999998 3.3 0.0016321999999999999 0 0.00163212 0 0.00163222 3.3 0.0016321399999999998 3.3 0.0016322399999999999 0 0.00163216 0 0.00163226 3.3 0.00163218 3.3 0.00163228 0 0.0016321999999999999 0 0.0016323 3.3 0.00163222 3.3 0.00163232 0 0.0016322399999999999 0 0.00163234 3.3 0.00163226 3.3 0.00163236 0 0.0016322799999999998 0 0.00163238 3.3 0.0016323 3.3 0.0016324 0 0.0016323199999999998 0 0.0016324199999999999 3.3 0.00163234 3.3 0.00163244 0 0.00163236 0 0.00163246 3.3 0.00163238 3.3 0.00163248 0 0.0016324 0 0.0016325 3.3 0.0016324199999999999 3.3 0.00163252 0 0.00163244 0 0.00163254 3.3 0.0016324599999999999 3.3 0.00163256 0 0.00163248 0 0.00163258 3.3 0.0016324999999999998 3.3 0.0016326 0 0.00163252 0 0.00163262 3.3 0.0016325399999999998 3.3 0.0016326399999999999 0 0.00163256 0 0.00163266 3.3 0.00163258 3.3 0.00163268 0 0.0016326 0 0.0016327 3.3 0.00163262 3.3 0.00163272 0 0.0016326399999999999 0 0.00163274 3.3 0.00163266 3.3 0.00163276 0 0.0016326799999999999 0 0.00163278 3.3 0.0016327 3.3 0.0016328 0 0.0016327199999999998 0 0.0016328199999999999 3.3 0.00163274 3.3 0.00163284 0 0.0016327599999999998 0 0.0016328599999999999 3.3 0.00163278 3.3 0.00163288 0 0.0016328 0 0.0016329 3.3 0.0016328199999999999 3.3 0.00163292 0 0.00163284 0 0.00163294 3.3 0.0016328599999999999 3.3 0.00163296 0 0.00163288 0 0.00163298 3.3 0.0016328999999999998 3.3 0.001633 0 0.00163292 0 0.00163302 3.3 0.0016329399999999998 3.3 0.0016330399999999999 0 0.00163296 0 0.00163306 3.3 0.0016329799999999998 3.3 0.0016330799999999999 0 0.001633 0 0.0016331 3.3 0.00163302 3.3 0.00163312 0 0.0016330399999999999 0 0.00163314 3.3 0.00163306 3.3 0.00163316 0 0.0016330799999999999 0 0.00163318 3.3 0.0016331 3.3 0.0016332 0 0.0016331199999999998 0 0.00163322 3.3 0.00163314 3.3 0.00163324 0 0.0016331599999999998 0 0.0016332599999999999 3.3 0.00163318 3.3 0.00163328 0 0.0016332 0 0.0016333 3.3 0.00163322 3.3 0.00163332 0 0.00163324 0 0.00163334 3.3 0.0016332599999999999 3.3 0.00163336 0 0.00163328 0 0.00163338 3.3 0.0016332999999999999 3.3 0.0016334 0 0.00163332 0 0.00163342 3.3 0.0016333399999999998 3.3 0.00163344 0 0.00163336 0 0.00163346 3.3 0.0016333799999999998 3.3 0.0016334799999999999 0 0.0016334 0 0.0016335 3.3 0.00163342 3.3 0.00163352 0 0.00163344 0 0.00163354 3.3 0.00163346 3.3 0.00163356 0 0.0016334799999999999 0 0.00163358 3.3 0.0016335 3.3 0.0016336 0 0.0016335199999999999 0 0.00163362 3.3 0.00163354 3.3 0.00163364 0 0.0016335599999999998 0 0.0016336599999999999 3.3 0.00163358 3.3 0.00163368 0 0.0016335999999999998 0 0.0016336999999999999 3.3 0.00163362 3.3 0.00163372 0 0.00163364 0 0.00163374 3.3 0.0016336599999999999 3.3 0.00163376 0 0.00163368 0 0.00163378 3.3 0.0016336999999999999 3.3 0.0016338 0 0.00163372 0 0.00163382 3.3 0.0016337399999999998 3.3 0.00163384 0 0.00163376 0 0.00163386 3.3 0.0016337799999999998 3.3 0.0016338799999999999 0 0.0016338 0 0.0016339 3.3 0.0016338199999999998 3.3 0.0016339199999999999 0 0.00163384 0 0.00163394 3.3 0.00163386 3.3 0.00163396 0 0.0016338799999999999 0 0.00163398 3.3 0.0016339 3.3 0.001634 0 0.0016339199999999999 0 0.00163402 3.3 0.00163394 3.3 0.00163404 0 0.0016339599999999998 0 0.00163406 3.3 0.00163398 3.3 0.00163408 0 0.0016339999999999998 0 0.0016340999999999999 3.3 0.00163402 3.3 0.00163412 0 0.00163404 0 0.00163414 3.3 0.00163406 3.3 0.00163416 0 0.00163408 0 0.00163418 3.3 0.0016340999999999999 3.3 0.0016342 0 0.00163412 0 0.00163422 3.3 0.0016341399999999999 3.3 0.00163424 0 0.00163416 0 0.00163426 3.3 0.0016341799999999998 3.3 0.0016342799999999999 0 0.0016342 0 0.0016343 3.3 0.0016342199999999998 3.3 0.0016343199999999999 0 0.00163424 0 0.00163434 3.3 0.00163426 3.3 0.00163436 0 0.0016342799999999999 0 0.00163438 3.3 0.0016343 3.3 0.0016344 0 0.0016343199999999999 0 0.00163442 3.3 0.00163434 3.3 0.00163444 0 0.0016343599999999998 0 0.00163446 3.3 0.00163438 3.3 0.00163448 0 0.0016343999999999998 0 0.0016344999999999999 3.3 0.00163442 3.3 0.00163452 0 0.0016344399999999998 0 0.0016345399999999999 3.3 0.00163446 3.3 0.00163456 0 0.00163448 0 0.00163458 3.3 0.0016344999999999999 3.3 0.0016346 0 0.00163452 0 0.00163462 3.3 0.0016345399999999999 3.3 0.00163464 0 0.00163456 0 0.00163466 3.3 0.0016345799999999998 3.3 0.00163468 0 0.0016346 0 0.0016347 3.3 0.0016346199999999998 3.3 0.0016347199999999999 0 0.00163464 0 0.00163474 3.3 0.0016346599999999998 3.3 0.0016347599999999999 0 0.00163468 0 0.00163478 3.3 0.0016347 3.3 0.0016348 0 0.0016347199999999999 0 0.00163482 3.3 0.00163474 3.3 0.00163484 0 0.0016347599999999999 0 0.00163486 3.3 0.00163478 3.3 0.00163488 0 0.0016347999999999998 0 0.0016349 3.3 0.00163482 3.3 0.00163492 0 0.0016348399999999998 0 0.0016349399999999999 3.3 0.00163486 3.3 0.00163496 0 0.00163488 0 0.00163498 3.3 0.0016349 3.3 0.001635 0 0.00163492 0 0.00163502 3.3 0.0016349399999999999 3.3 0.00163504 0 0.00163496 0 0.00163506 3.3 0.0016349799999999999 3.3 0.00163508 0 0.001635 0 0.0016351 3.3 0.0016350199999999998 3.3 0.0016351199999999999 0 0.00163504 0 0.00163514 3.3 0.0016350599999999998 3.3 0.0016351599999999999 0 0.00163508 0 0.00163518 3.3 0.0016351 3.3 0.0016352 0 0.0016351199999999999 0 0.00163522 3.3 0.00163514 3.3 0.00163524 0 0.0016351599999999999 0 0.00163526 3.3 0.00163518 3.3 0.00163528 0 0.0016351999999999998 0 0.0016353 3.3 0.00163522 3.3 0.00163532 0 0.0016352399999999998 0 0.0016353399999999999 3.3 0.00163526 3.3 0.00163536 0 0.0016352799999999998 0 0.0016353799999999999 3.3 0.0016353 3.3 0.0016354 0 0.00163532 0 0.00163542 3.3 0.0016353399999999999 3.3 0.00163544 0 0.00163536 0 0.00163546 3.3 0.0016353799999999999 3.3 0.00163548 0 0.0016354 0 0.0016355 3.3 0.0016354199999999998 3.3 0.00163552 0 0.00163544 0 0.00163554 3.3 0.0016354599999999998 3.3 0.0016355599999999999 0 0.00163548 0 0.00163558 3.3 0.0016355 3.3 0.0016356 0 0.00163552 0 0.00163562 3.3 0.00163554 3.3 0.00163564 0 0.0016355599999999999 0 0.00163566 3.3 0.00163558 3.3 0.00163568 0 0.0016355999999999999 0 0.0016357 3.3 0.00163562 3.3 0.00163572 0 0.0016356399999999998 0 0.00163574 3.3 0.00163566 3.3 0.00163576 0 0.0016356799999999998 0 0.0016357799999999999 3.3 0.0016357 3.3 0.0016358 0 0.00163572 0 0.00163582 3.3 0.00163574 3.3 0.00163584 0 0.00163576 0 0.00163586 3.3 0.0016357799999999999 3.3 0.00163588 0 0.0016358 0 0.0016359 3.3 0.0016358199999999999 3.3 0.00163592 0 0.00163584 0 0.00163594 3.3 0.0016358599999999998 3.3 0.0016359599999999999 0 0.00163588 0 0.00163598 3.3 0.0016358999999999998 3.3 0.0016359999999999999 0 0.00163592 0 0.00163602 3.3 0.00163594 3.3 0.00163604 0 0.0016359599999999999 0 0.00163606 3.3 0.00163598 3.3 0.00163608 0 0.0016359999999999999 0 0.0016361 3.3 0.00163602 3.3 0.00163612 0 0.0016360399999999998 0 0.00163614 3.3 0.00163606 3.3 0.00163616 0 0.0016360799999999998 0 0.0016361799999999999 3.3 0.0016361 3.3 0.0016362 0 0.0016361199999999998 0 0.0016362199999999999 3.3 0.00163614 3.3 0.00163624 0 0.00163616 0 0.00163626 3.3 0.0016361799999999999 3.3 0.00163628 0 0.0016362 0 0.0016363 3.3 0.0016362199999999999 3.3 0.00163632 0 0.00163624 0 0.00163634 3.3 0.0016362599999999998 3.3 0.00163636 0 0.00163628 0 0.00163638 3.3 0.0016362999999999998 3.3 0.0016363999999999999 0 0.00163632 0 0.00163642 3.3 0.00163634 3.3 0.00163644 0 0.00163636 0 0.00163646 3.3 0.00163638 3.3 0.00163648 0 0.0016363999999999999 0 0.0016365 3.3 0.00163642 3.3 0.00163652 0 0.0016364399999999999 0 0.00163654 3.3 0.00163646 3.3 0.00163656 0 0.0016364799999999998 0 0.00163658 3.3 0.0016365 3.3 0.0016366 0 0.0016365199999999998 0 0.0016366199999999999 3.3 0.00163654 3.3 0.00163664 0 0.00163656 0 0.00163666 3.3 0.00163658 3.3 0.00163668 0 0.0016366 0 0.0016367 3.3 0.0016366199999999999 3.3 0.00163672 0 0.00163664 0 0.00163674 3.3 0.0016366599999999999 3.3 0.00163676 0 0.00163668 0 0.00163678 3.3 0.0016366999999999998 3.3 0.0016367999999999999 0 0.00163672 0 0.00163682 3.3 0.0016367399999999998 3.3 0.0016368399999999999 0 0.00163676 0 0.00163686 3.3 0.00163678 3.3 0.00163688 0 0.0016367999999999999 0 0.0016369 3.3 0.00163682 3.3 0.00163692 0 0.0016368399999999999 0 0.00163694 3.3 0.00163686 3.3 0.00163696 0 0.0016368799999999998 0 0.00163698 3.3 0.0016369 3.3 0.001637 0 0.0016369199999999998 0 0.0016370199999999999 3.3 0.00163694 3.3 0.00163704 0 0.0016369599999999998 0 0.0016370599999999999 3.3 0.00163698 3.3 0.00163708 0 0.001637 0 0.0016371 3.3 0.0016370199999999999 3.3 0.00163712 0 0.00163704 0 0.00163714 3.3 0.0016370599999999999 3.3 0.00163716 0 0.00163708 0 0.00163718 3.3 0.0016370999999999998 3.3 0.0016372 0 0.00163712 0 0.00163722 3.3 0.0016371399999999998 3.3 0.0016372399999999999 0 0.00163716 0 0.00163726 3.3 0.00163718 3.3 0.00163728 0 0.0016372 0 0.0016373 3.3 0.00163722 3.3 0.00163732 0 0.0016372399999999999 0 0.00163734 3.3 0.00163726 3.3 0.00163736 0 0.0016372799999999999 0 0.00163738 3.3 0.0016373 3.3 0.0016374 0 0.0016373199999999998 0 0.0016374199999999999 3.3 0.00163734 3.3 0.00163744 0 0.0016373599999999998 0 0.0016374599999999999 3.3 0.00163738 3.3 0.00163748 0 0.0016374 0 0.0016375 3.3 0.0016374199999999999 3.3 0.00163752 0 0.00163744 0 0.00163754 3.3 0.0016374599999999999 3.3 0.00163756 0 0.00163748 0 0.00163758 3.3 0.0016374999999999998 3.3 0.0016376 0 0.00163752 0 0.00163762 3.3 0.0016375399999999998 3.3 0.0016376399999999999 0 0.00163756 0 0.00163766 3.3 0.0016375799999999998 3.3 0.0016376799999999999 0 0.0016376 0 0.0016377 3.3 0.00163762 3.3 0.00163772 0 0.0016376399999999999 0 0.00163774 3.3 0.00163766 3.3 0.00163776 0 0.0016376799999999999 0 0.00163778 3.3 0.0016377 3.3 0.0016378 0 0.0016377199999999998 0 0.00163782 3.3 0.00163774 3.3 0.00163784 0 0.0016377599999999998 0 0.0016378599999999999 3.3 0.00163778 3.3 0.00163788 0 0.0016377999999999998 0 0.0016378999999999999 3.3 0.00163782 3.3 0.00163792 0 0.00163784 0 0.00163794 3.3 0.0016378599999999999 3.3 0.00163796 0 0.00163788 0 0.00163798 3.3 0.0016378999999999999 3.3 0.001638 0 0.00163792 0 0.00163802 3.3 0.0016379399999999998 3.3 0.00163804 0 0.00163796 0 0.00163806 3.3 0.0016379799999999998 3.3 0.0016380799999999999 0 0.001638 0 0.0016381 3.3 0.00163802 3.3 0.00163812 0 0.00163804 0 0.00163814 3.3 0.00163806 3.3 0.00163816 0 0.0016380799999999999 0 0.00163818 3.3 0.0016381 3.3 0.0016382 0 0.0016381199999999999 0 0.00163822 3.3 0.00163814 3.3 0.00163824 0 0.0016381599999999998 0 0.0016382599999999999 3.3 0.00163818 3.3 0.00163828 0 0.0016381999999999998 0 0.0016382999999999999 3.3 0.00163822 3.3 0.00163832 0 0.00163824 0 0.00163834 3.3 0.0016382599999999999 3.3 0.00163836 0 0.00163828 0 0.00163838 3.3 0.0016382999999999999 3.3 0.0016384 0 0.00163832 0 0.00163842 3.3 0.0016383399999999998 3.3 0.00163844 0 0.00163836 0 0.00163846 3.3 0.0016383799999999998 3.3 0.0016384799999999999 0 0.0016384 0 0.0016385 3.3 0.0016384199999999998 3.3 0.0016385199999999999 0 0.00163844 0 0.00163854 3.3 0.00163846 3.3 0.00163856 0 0.0016384799999999999 0 0.00163858 3.3 0.0016385 3.3 0.0016386 0 0.0016385199999999999 0 0.00163862 3.3 0.00163854 3.3 0.00163864 0 0.0016385599999999998 0 0.00163866 3.3 0.00163858 3.3 0.00163868 0 0.0016385999999999998 0 0.0016386999999999999 3.3 0.00163862 3.3 0.00163872 0 0.00163864 0 0.00163874 3.3 0.00163866 3.3 0.00163876 0 0.00163868 0 0.00163878 3.3 0.0016386999999999999 3.3 0.0016388 0 0.00163872 0 0.00163882 3.3 0.0016387399999999999 3.3 0.00163884 0 0.00163876 0 0.00163886 3.3 0.0016387799999999998 3.3 0.00163888 0 0.0016388 0 0.0016389 3.3 0.0016388199999999998 3.3 0.0016389199999999999 0 0.00163884 0 0.00163894 3.3 0.00163886 3.3 0.00163896 0 0.00163888 0 0.00163898 3.3 0.0016389 3.3 0.001639 0 0.0016389199999999999 0 0.00163902 3.3 0.00163894 3.3 0.00163904 0 0.0016389599999999999 0 0.00163906 3.3 0.00163898 3.3 0.00163908 0 0.0016389999999999998 0 0.0016390999999999999 3.3 0.00163902 3.3 0.00163912 0 0.0016390399999999998 0 0.0016391399999999999 3.3 0.00163906 3.3 0.00163916 0 0.00163908 0 0.00163918 3.3 0.0016390999999999999 3.3 0.0016392 0 0.00163912 0 0.00163922 3.3 0.0016391399999999999 3.3 0.00163924 0 0.00163916 0 0.00163926 3.3 0.0016391799999999998 3.3 0.00163928 0 0.0016392 0 0.0016393 3.3 0.0016392199999999998 3.3 0.0016393199999999999 0 0.00163924 0 0.00163934 3.3 0.0016392599999999998 3.3 0.0016393599999999999 0 0.00163928 0 0.00163938 3.3 0.0016393 3.3 0.0016394 0 0.0016393199999999999 0 0.00163942 3.3 0.00163934 3.3 0.00163944 0 0.0016393599999999999 0 0.00163946 3.3 0.00163938 3.3 0.00163948 0 0.0016393999999999998 0 0.0016395 3.3 0.00163942 3.3 0.00163952 0 0.0016394399999999998 0 0.0016395399999999999 3.3 0.00163946 3.3 0.00163956 0 0.00163948 0 0.00163958 3.3 0.0016395 3.3 0.0016396 0 0.00163952 0 0.00163962 3.3 0.0016395399999999999 3.3 0.00163964 0 0.00163956 0 0.00163966 3.3 0.0016395799999999999 3.3 0.00163968 0 0.0016396 0 0.0016397 3.3 0.0016396199999999998 3.3 0.00163972 0 0.00163964 0 0.00163974 3.3 0.0016396599999999998 3.3 0.0016397599999999999 0 0.00163968 0 0.00163978 3.3 0.0016397 3.3 0.0016398 0 0.00163972 0 0.00163982 3.3 0.00163974 3.3 0.00163984 0 0.0016397599999999999 0 0.00163986 3.3 0.00163978 3.3 0.00163988 0 0.0016397999999999999 0 0.0016399 3.3 0.00163982 3.3 0.00163992 0 0.0016398399999999998 0 0.0016399399999999999 3.3 0.00163986 3.3 0.00163996 0 0.0016398799999999998 0 0.0016399799999999999 3.3 0.0016399 3.3 0.00164 0 0.00163992 0 0.00164002 3.3 0.0016399399999999999 3.3 0.00164004 0 0.00163996 0 0.00164006 3.3 0.0016399799999999999 3.3 0.00164008 0 0.00164 0 0.0016401 3.3 0.0016400199999999998 3.3 0.00164012 0 0.00164004 0 0.00164014 3.3 0.0016400599999999998 3.3 0.0016401599999999999 0 0.00164008 0 0.00164018 3.3 0.0016400999999999998 3.3 0.0016401999999999999 0 0.00164012 0 0.00164022 3.3 0.00164014 3.3 0.00164024 0 0.0016401599999999999 0 0.00164026 3.3 0.00164018 3.3 0.00164028 0 0.0016401999999999999 0 0.0016403 3.3 0.00164022 3.3 0.00164032 0 0.0016402399999999998 0 0.00164034 3.3 0.00164026 3.3 0.00164036 0 0.0016402799999999998 0 0.0016403799999999999 3.3 0.0016403 3.3 0.0016404 0 0.00164032 0 0.00164042 3.3 0.00164034 3.3 0.00164044 0 0.00164036 0 0.00164046 3.3 0.0016403799999999999 3.3 0.00164048 0 0.0016404 0 0.0016405 3.3 0.0016404199999999999 3.3 0.00164052 0 0.00164044 0 0.00164054 3.3 0.0016404599999999998 3.3 0.00164056 0 0.00164048 0 0.00164058 3.3 0.0016404999999999998 3.3 0.0016405999999999999 0 0.00164052 0 0.00164062 3.3 0.00164054 3.3 0.00164064 0 0.00164056 0 0.00164066 3.3 0.00164058 3.3 0.00164068 0 0.0016405999999999999 0 0.0016407 3.3 0.00164062 3.3 0.00164072 0 0.0016406399999999999 0 0.00164074 3.3 0.00164066 3.3 0.00164076 0 0.0016406799999999998 0 0.0016407799999999999 3.3 0.0016407 3.3 0.0016408 0 0.0016407199999999998 0 0.0016408199999999999 3.3 0.00164074 3.3 0.00164084 0 0.00164076 0 0.00164086 3.3 0.0016407799999999999 3.3 0.00164088 0 0.0016408 0 0.0016409 3.3 0.0016408199999999999 3.3 0.00164092 0 0.00164084 0 0.00164094 3.3 0.0016408599999999998 3.3 0.00164096 0 0.00164088 0 0.00164098 3.3 0.0016408999999999998 3.3 0.0016409999999999999 0 0.00164092 0 0.00164102 3.3 0.0016409399999999998 3.3 0.0016410399999999999 0 0.00164096 0 0.00164106 3.3 0.00164098 3.3 0.00164108 0 0.0016409999999999999 0 0.0016411 3.3 0.00164102 3.3 0.00164112 0 0.0016410399999999999 0 0.00164114 3.3 0.00164106 3.3 0.00164116 0 0.0016410799999999998 0 0.00164118 3.3 0.0016411 3.3 0.0016412 0 0.0016411199999999998 0 0.0016412199999999999 3.3 0.00164114 3.3 0.00164124 0 0.00164116 0 0.00164126 3.3 0.00164118 3.3 0.00164128 0 0.0016412 0 0.0016413 3.3 0.0016412199999999999 3.3 0.00164132 0 0.00164124 0 0.00164134 3.3 0.0016412599999999999 3.3 0.00164136 0 0.00164128 0 0.00164138 3.3 0.0016412999999999998 3.3 0.0016413999999999999 0 0.00164132 0 0.00164142 3.3 0.0016413399999999998 3.3 0.0016414399999999999 0 0.00164136 0 0.00164146 3.3 0.00164138 3.3 0.00164148 0 0.0016413999999999999 0 0.0016415 3.3 0.00164142 3.3 0.00164152 0 0.0016414399999999999 0 0.00164154 3.3 0.00164146 3.3 0.00164156 0 0.0016414799999999998 0 0.00164158 3.3 0.0016415 3.3 0.0016416 0 0.0016415199999999998 0 0.0016416199999999999 3.3 0.00164154 3.3 0.00164164 0 0.0016415599999999998 0 0.0016416599999999999 3.3 0.00164158 3.3 0.00164168 0 0.0016416 0 0.0016417 3.3 0.0016416199999999999 3.3 0.00164172 0 0.00164164 0 0.00164174 3.3 0.0016416599999999999 3.3 0.00164176 0 0.00164168 0 0.00164178 3.3 0.0016416999999999998 3.3 0.0016418 0 0.00164172 0 0.00164182 3.3 0.0016417399999999998 3.3 0.0016418399999999999 0 0.00164176 0 0.00164186 3.3 0.0016417799999999998 3.3 0.0016418799999999999 0 0.0016418 0 0.0016419 3.3 0.00164182 3.3 0.00164192 0 0.0016418399999999999 0 0.00164194 3.3 0.00164186 3.3 0.00164196 0 0.0016418799999999999 0 0.00164198 3.3 0.0016419 3.3 0.001642 0 0.0016419199999999998 0 0.00164202 3.3 0.00164194 3.3 0.00164204 0 0.0016419599999999998 0 0.0016420599999999999 3.3 0.00164198 3.3 0.00164208 0 0.001642 0 0.0016421 3.3 0.00164202 3.3 0.00164212 0 0.00164204 0 0.00164214 3.3 0.0016420599999999999 3.3 0.00164216 0 0.00164208 0 0.00164218 3.3 0.0016420999999999999 3.3 0.0016422 0 0.00164212 0 0.00164222 3.3 0.0016421399999999998 3.3 0.0016422399999999999 0 0.00164216 0 0.00164226 3.3 0.0016421799999999998 3.3 0.0016422799999999999 0 0.0016422 0 0.0016423 3.3 0.00164222 3.3 0.00164232 0 0.0016422399999999999 0 0.00164234 3.3 0.00164226 3.3 0.00164236 0 0.0016422799999999999 0 0.00164238 3.3 0.0016423 3.3 0.0016424 0 0.0016423199999999998 0 0.00164242 3.3 0.00164234 3.3 0.00164244 0 0.0016423599999999998 0 0.0016424599999999999 3.3 0.00164238 3.3 0.00164248 0 0.0016423999999999998 0 0.0016424999999999999 3.3 0.00164242 3.3 0.00164252 0 0.00164244 0 0.00164254 3.3 0.0016424599999999999 3.3 0.00164256 0 0.00164248 0 0.00164258 3.3 0.0016424999999999999 3.3 0.0016426 0 0.00164252 0 0.00164262 3.3 0.0016425399999999998 3.3 0.00164264 0 0.00164256 0 0.00164266 3.3 0.0016425799999999998 3.3 0.0016426799999999999 0 0.0016426 0 0.0016427 3.3 0.00164262 3.3 0.00164272 0 0.00164264 0 0.00164274 3.3 0.00164266 3.3 0.00164276 0 0.0016426799999999999 0 0.00164278 3.3 0.0016427 3.3 0.0016428 0 0.0016427199999999999 0 0.00164282 3.3 0.00164274 3.3 0.00164284 0 0.0016427599999999998 0 0.00164286 3.3 0.00164278 3.3 0.00164288 0 0.0016427999999999998 0 0.0016428999999999999 3.3 0.00164282 3.3 0.00164292 0 0.00164284 0 0.00164294 3.3 0.00164286 3.3 0.00164296 0 0.00164288 0 0.00164298 3.3 0.0016428999999999999 3.3 0.001643 0 0.00164292 0 0.00164302 3.3 0.0016429399999999999 3.3 0.00164304 0 0.00164296 0 0.00164306 3.3 0.0016429799999999998 3.3 0.0016430799999999999 0 0.001643 0 0.0016431 3.3 0.0016430199999999998 3.3 0.0016431199999999999 0 0.00164304 0 0.00164314 3.3 0.00164306 3.3 0.00164316 0 0.0016430799999999999 0 0.00164318 3.3 0.0016431 3.3 0.0016432 0 0.0016431199999999999 0 0.00164322 3.3 0.00164314 3.3 0.00164324 0 0.0016431599999999998 0 0.00164326 3.3 0.00164318 3.3 0.00164328 0 0.0016431999999999998 0 0.0016432999999999999 3.3 0.00164322 3.3 0.00164332 0 0.0016432399999999998 0 0.0016433399999999999 3.3 0.00164326 3.3 0.00164336 0 0.00164328 0 0.00164338 3.3 0.0016432999999999999 3.3 0.0016434 0 0.00164332 0 0.00164342 3.3 0.0016433399999999999 3.3 0.00164344 0 0.00164336 0 0.00164346 3.3 0.0016433799999999998 3.3 0.00164348 0 0.0016434 0 0.0016435 3.3 0.0016434199999999998 3.3 0.0016435199999999999 0 0.00164344 0 0.00164354 3.3 0.00164346 3.3 0.00164356 0 0.00164348 0 0.00164358 3.3 0.0016435 3.3 0.0016436 0 0.0016435199999999999 0 0.00164362 3.3 0.00164354 3.3 0.00164364 0 0.0016435599999999999 0 0.00164366 3.3 0.00164358 3.3 0.00164368 0 0.0016435999999999998 0 0.0016437 3.3 0.00164362 3.3 0.00164372 0 0.0016436399999999998 0 0.0016437399999999999 3.3 0.00164366 3.3 0.00164376 0 0.00164368 0 0.00164378 3.3 0.0016437 3.3 0.0016438 0 0.00164372 0 0.00164382 3.3 0.0016437399999999999 3.3 0.00164384 0 0.00164376 0 0.00164386 3.3 0.0016437799999999999 3.3 0.00164388 0 0.0016438 0 0.0016439 3.3 0.0016438199999999998 3.3 0.0016439199999999999 0 0.00164384 0 0.00164394 3.3 0.0016438599999999998 3.3 0.0016439599999999999 0 0.00164388 0 0.00164398 3.3 0.0016439 3.3 0.001644 0 0.0016439199999999999 0 0.00164402 3.3 0.00164394 3.3 0.00164404 0 0.0016439599999999999 0 0.00164406 3.3 0.00164398 3.3 0.00164408 0 0.0016439999999999998 0 0.0016441 3.3 0.00164402 3.3 0.00164412 0 0.0016440399999999998 0 0.0016441399999999999 3.3 0.00164406 3.3 0.00164416 0 0.0016440799999999998 0 0.0016441799999999999 3.3 0.0016441 3.3 0.0016442 0 0.00164412 0 0.00164422 3.3 0.0016441399999999999 3.3 0.00164424 0 0.00164416 0 0.00164426 3.3 0.0016441799999999999 3.3 0.00164428 0 0.0016442 0 0.0016443 3.3 0.0016442199999999998 3.3 0.00164432 0 0.00164424 0 0.00164434 3.3 0.0016442599999999998 3.3 0.0016443599999999999 0 0.00164428 0 0.00164438 3.3 0.0016443 3.3 0.0016444 0 0.00164432 0 0.00164442 3.3 0.00164434 3.3 0.00164444 0 0.0016443599999999999 0 0.00164446 3.3 0.00164438 3.3 0.00164448 0 0.0016443999999999999 0 0.0016445 3.3 0.00164442 3.3 0.00164452 0 0.0016444399999999998 0 0.0016445399999999999 3.3 0.00164446 3.3 0.00164456 0 0.0016444799999999998 0 0.0016445799999999999 3.3 0.0016445 3.3 0.0016446 0 0.00164452 0 0.00164462 3.3 0.0016445399999999999 3.3 0.00164464 0 0.00164456 0 0.00164466 3.3 0.0016445799999999999 3.3 0.00164468 0 0.0016446 0 0.0016447 3.3 0.0016446199999999998 3.3 0.00164472 0 0.00164464 0 0.00164474 3.3 0.0016446599999999998 3.3 0.0016447599999999999 0 0.00164468 0 0.00164478 3.3 0.0016446999999999998 3.3 0.0016447999999999999 0 0.00164472 0 0.00164482 3.3 0.00164474 3.3 0.00164484 0 0.0016447599999999999 0 0.00164486 3.3 0.00164478 3.3 0.00164488 0 0.0016447999999999999 0 0.0016449 3.3 0.00164482 3.3 0.00164492 0 0.0016448399999999998 0 0.00164494 3.3 0.00164486 3.3 0.00164496 0 0.0016448799999999998 0 0.0016449799999999999 3.3 0.0016449 3.3 0.001645 0 0.0016449199999999998 0 0.0016450199999999999 3.3 0.00164494 3.3 0.00164504 0 0.00164496 0 0.00164506 3.3 0.0016449799999999999 3.3 0.00164508 0 0.001645 0 0.0016451 3.3 0.0016450199999999999 3.3 0.00164512 0 0.00164504 0 0.00164514 3.3 0.0016450599999999998 3.3 0.00164516 0 0.00164508 0 0.00164518 3.3 0.0016450999999999998 3.3 0.0016451999999999999 0 0.00164512 0 0.00164522 3.3 0.00164514 3.3 0.00164524 0 0.00164516 0 0.00164526 3.3 0.00164518 3.3 0.00164528 0 0.0016451999999999999 0 0.0016453 3.3 0.00164522 3.3 0.00164532 0 0.0016452399999999999 0 0.00164534 3.3 0.00164526 3.3 0.00164536 0 0.0016452799999999998 0 0.0016453799999999999 3.3 0.0016453 3.3 0.0016454 0 0.0016453199999999998 0 0.0016454199999999999 3.3 0.00164534 3.3 0.00164544 0 0.00164536 0 0.00164546 3.3 0.0016453799999999999 3.3 0.00164548 0 0.0016454 0 0.0016455 3.3 0.0016454199999999999 3.3 0.00164552 0 0.00164544 0 0.00164554 3.3 0.0016454599999999998 3.3 0.00164556 0 0.00164548 0 0.00164558 3.3 0.0016454999999999998 3.3 0.0016455999999999999 0 0.00164552 0 0.00164562 3.3 0.0016455399999999998 3.3 0.0016456399999999999 0 0.00164556 0 0.00164566 3.3 0.00164558 3.3 0.00164568 0 0.0016455999999999999 0 0.0016457 3.3 0.00164562 3.3 0.00164572 0 0.0016456399999999999 0 0.00164574 3.3 0.00164566 3.3 0.00164576 0 0.0016456799999999998 0 0.00164578 3.3 0.0016457 3.3 0.0016458 0 0.0016457199999999998 0 0.0016458199999999999 3.3 0.00164574 3.3 0.00164584 0 0.00164576 0 0.00164586 3.3 0.00164578 3.3 0.00164588 0 0.0016458 0 0.0016459 3.3 0.0016458199999999999 3.3 0.00164592 0 0.00164584 0 0.00164594 3.3 0.0016458599999999999 3.3 0.00164596 0 0.00164588 0 0.00164598 3.3 0.0016458999999999998 3.3 0.001646 0 0.00164592 0 0.00164602 3.3 0.0016459399999999998 3.3 0.0016460399999999999 0 0.00164596 0 0.00164606 3.3 0.00164598 3.3 0.00164608 0 0.001646 0 0.0016461 3.3 0.00164602 3.3 0.00164612 0 0.0016460399999999999 0 0.00164614 3.3 0.00164606 3.3 0.00164616 0 0.0016460799999999999 0 0.00164618 3.3 0.0016461 3.3 0.0016462 0 0.0016461199999999998 0 0.0016462199999999999 3.3 0.00164614 3.3 0.00164624 0 0.0016461599999999998 0 0.0016462599999999999 3.3 0.00164618 3.3 0.00164628 0 0.0016462 0 0.0016463 3.3 0.0016462199999999999 3.3 0.00164632 0 0.00164624 0 0.00164634 3.3 0.0016462599999999999 3.3 0.00164636 0 0.00164628 0 0.00164638 3.3 0.0016462999999999998 3.3 0.0016464 0 0.00164632 0 0.00164642 3.3 0.0016463399999999998 3.3 0.0016464399999999999 0 0.00164636 0 0.00164646 3.3 0.0016463799999999998 3.3 0.0016464799999999999 0 0.0016464 0 0.0016465 3.3 0.00164642 3.3 0.00164652 0 0.0016464399999999999 0 0.00164654 3.3 0.00164646 3.3 0.00164656 0 0.0016464799999999999 0 0.00164658 3.3 0.0016465 3.3 0.0016466 0 0.0016465199999999998 0 0.00164662 3.3 0.00164654 3.3 0.00164664 0 0.0016465599999999998 0 0.0016466599999999999 3.3 0.00164658 3.3 0.00164668 0 0.0016466 0 0.0016467 3.3 0.00164662 3.3 0.00164672 0 0.00164664 0 0.00164674 3.3 0.0016466599999999999 3.3 0.00164676 0 0.00164668 0 0.00164678 3.3 0.0016466999999999999 3.3 0.0016468 0 0.00164672 0 0.00164682 3.3 0.0016467399999999998 3.3 0.00164684 0 0.00164676 0 0.00164686 3.3 0.0016467799999999998 3.3 0.0016468799999999999 0 0.0016468 0 0.0016469 3.3 0.00164682 3.3 0.00164692 0 0.00164684 0 0.00164694 3.3 0.00164686 3.3 0.00164696 0 0.0016468799999999999 0 0.00164698 3.3 0.0016469 3.3 0.001647 0 0.0016469199999999999 0 0.00164702 3.3 0.00164694 3.3 0.00164704 0 0.0016469599999999998 0 0.0016470599999999999 3.3 0.00164698 3.3 0.00164708 0 0.0016469999999999998 0 0.0016470999999999999 3.3 0.00164702 3.3 0.00164712 0 0.00164704 0 0.00164714 3.3 0.0016470599999999999 3.3 0.00164716 0 0.00164708 0 0.00164718 3.3 0.0016470999999999999 3.3 0.0016472 0 0.00164712 0 0.00164722 3.3 0.0016471399999999998 3.3 0.00164724 0 0.00164716 0 0.00164726 3.3 0.0016471799999999998 3.3 0.0016472799999999999 0 0.0016472 0 0.0016473 3.3 0.0016472199999999998 3.3 0.0016473199999999999 0 0.00164724 0 0.00164734 3.3 0.00164726 3.3 0.00164736 0 0.0016472799999999999 0 0.00164738 3.3 0.0016473 3.3 0.0016474 0 0.0016473199999999999 0 0.00164742 3.3 0.00164734 3.3 0.00164744 0 0.0016473599999999998 0 0.00164746 3.3 0.00164738 3.3 0.00164748 0 0.0016473999999999998 0 0.0016474999999999999 3.3 0.00164742 3.3 0.00164752 0 0.00164744 0 0.00164754 3.3 0.00164746 3.3 0.00164756 0 0.00164748 0 0.00164758 3.3 0.0016474999999999999 3.3 0.0016476 0 0.00164752 0 0.00164762 3.3 0.0016475399999999999 3.3 0.00164764 0 0.00164756 0 0.00164766 3.3 0.0016475799999999998 3.3 0.0016476799999999999 0 0.0016476 0 0.0016477 3.3 0.0016476199999999998 3.3 0.0016477199999999999 0 0.00164764 0 0.00164774 3.3 0.00164766 3.3 0.00164776 0 0.0016476799999999999 0 0.00164778 3.3 0.0016477 3.3 0.0016478 0 0.0016477199999999999 0 0.00164782 3.3 0.00164774 3.3 0.00164784 0 0.0016477599999999998 0 0.00164786 3.3 0.00164778 3.3 0.00164788 0 0.0016477999999999998 0 0.0016478999999999999 3.3 0.00164782 3.3 0.00164792 0 0.0016478399999999998 0 0.0016479399999999999 3.3 0.00164786 3.3 0.00164796 0 0.00164788 0 0.00164798 3.3 0.0016478999999999999 3.3 0.001648 0 0.00164792 0 0.00164802 3.3 0.0016479399999999999 3.3 0.00164804 0 0.00164796 0 0.00164806 3.3 0.0016479799999999998 3.3 0.00164808 0 0.001648 0 0.0016481 3.3 0.0016480199999999998 3.3 0.0016481199999999999 0 0.00164804 0 0.00164814 3.3 0.0016480599999999998 3.3 0.0016481599999999999 0 0.00164808 0 0.00164818 3.3 0.0016481 3.3 0.0016482 0 0.0016481199999999999 0 0.00164822 3.3 0.00164814 3.3 0.00164824 0 0.0016481599999999999 0 0.00164826 3.3 0.00164818 3.3 0.00164828 0 0.0016481999999999998 0 0.0016483 3.3 0.00164822 3.3 0.00164832 0 0.0016482399999999998 0 0.0016483399999999999 3.3 0.00164826 3.3 0.00164836 0 0.00164828 0 0.00164838 3.3 0.0016483 3.3 0.0016484 0 0.00164832 0 0.00164842 3.3 0.0016483399999999999 3.3 0.00164844 0 0.00164836 0 0.00164846 3.3 0.0016483799999999999 3.3 0.00164848 0 0.0016484 0 0.0016485 3.3 0.0016484199999999998 3.3 0.0016485199999999999 0 0.00164844 0 0.00164854 3.3 0.0016484599999999998 3.3 0.0016485599999999999 0 0.00164848 0 0.00164858 3.3 0.0016485 3.3 0.0016486 0 0.0016485199999999999 0 0.00164862 3.3 0.00164854 3.3 0.00164864 0 0.0016485599999999999 0 0.00164866 3.3 0.00164858 3.3 0.00164868 0 0.0016485999999999998 0 0.0016487 3.3 0.00164862 3.3 0.00164872 0 0.0016486399999999998 0 0.0016487399999999999 3.3 0.00164866 3.3 0.00164876 0 0.0016486799999999998 0 0.0016487799999999999 3.3 0.0016487 3.3 0.0016488 0 0.00164872 0 0.00164882 3.3 0.0016487399999999999 3.3 0.00164884 0 0.00164876 0 0.00164886 3.3 0.0016487799999999999 3.3 0.00164888 0 0.0016488 0 0.0016489 3.3 0.0016488199999999998 3.3 0.00164892 0 0.00164884 0 0.00164894 3.3 0.0016488599999999998 3.3 0.0016489599999999999 0 0.00164888 0 0.00164898 3.3 0.0016489 3.3 0.001649 0 0.00164892 0 0.00164902 3.3 0.00164894 3.3 0.00164904 0 0.0016489599999999999 0 0.00164906 3.3 0.00164898 3.3 0.00164908 0 0.0016489999999999999 0 0.0016491 3.3 0.00164902 3.3 0.00164912 0 0.0016490399999999998 0 0.00164914 3.3 0.00164906 3.3 0.00164916 0 0.0016490799999999998 0 0.0016491799999999999 3.3 0.0016491 3.3 0.0016492 0 0.00164912 0 0.00164922 3.3 0.00164914 3.3 0.00164924 0 0.00164916 0 0.00164926 3.3 0.0016491799999999999 3.3 0.00164928 0 0.0016492 0 0.0016493 3.3 0.0016492199999999999 3.3 0.00164932 0 0.00164924 0 0.00164934 3.3 0.0016492599999999998 3.3 0.0016493599999999999 0 0.00164928 0 0.00164938 3.3 0.0016492999999999998 3.3 0.0016493999999999999 0 0.00164932 0 0.00164942 3.3 0.00164934 3.3 0.00164944 0 0.0016493599999999999 0 0.00164946 3.3 0.00164938 3.3 0.00164948 0 0.0016493999999999999 0 0.0016495 3.3 0.00164942 3.3 0.00164952 0 0.0016494399999999998 0 0.00164954 3.3 0.00164946 3.3 0.00164956 0 0.0016494799999999998 0 0.0016495799999999999 3.3 0.0016495 3.3 0.0016496 0 0.0016495199999999998 0 0.0016496199999999999 3.3 0.00164954 3.3 0.00164964 0 0.00164956 0 0.00164966 3.3 0.0016495799999999999 3.3 0.00164968 0 0.0016496 0 0.0016497 3.3 0.0016496199999999999 3.3 0.00164972 0 0.00164964 0 0.00164974 3.3 0.0016496599999999998 3.3 0.00164976 0 0.00164968 0 0.00164978 3.3 0.0016496999999999998 3.3 0.0016497999999999999 0 0.00164972 0 0.00164982 3.3 0.00164974 3.3 0.00164984 0 0.00164976 0 0.00164986 3.3 0.00164978 3.3 0.00164988 0 0.0016497999999999999 0 0.0016499 3.3 0.00164982 3.3 0.00164992 0 0.0016498399999999999 0 0.00164994 3.3 0.00164986 3.3 0.00164996 0 0.0016498799999999998 0 0.00164998 3.3 0.0016499 3.3 0.00165 0 0.0016499199999999998 0 0.0016500199999999999 3.3 0.00164994 3.3 0.00165004 0 0.00164996 0 0.00165006 3.3 0.00164998 3.3 0.00165008 0 0.00165 0 0.0016501 3.3 0.0016500199999999999 3.3 0.00165012 0 0.00165004 0 0.00165014 3.3 0.0016500599999999999 3.3 0.00165016 0 0.00165008 0 0.00165018 3.3 0.0016500999999999998 3.3 0.0016501999999999999 0 0.00165012 0 0.00165022 3.3 0.0016501399999999998 3.3 0.0016502399999999999 0 0.00165016 0 0.00165026 3.3 0.00165018 3.3 0.00165028 0 0.0016501999999999999 0 0.0016503 3.3 0.00165022 3.3 0.00165032 0 0.0016502399999999999 0 0.00165034 3.3 0.00165026 3.3 0.00165036 0 0.0016502799999999998 0 0.00165038 3.3 0.0016503 3.3 0.0016504 0 0.0016503199999999998 0 0.0016504199999999999 3.3 0.00165034 3.3 0.00165044 0 0.0016503599999999998 0 0.0016504599999999999 3.3 0.00165038 3.3 0.00165048 0 0.0016504 0 0.0016505 3.3 0.0016504199999999999 3.3 0.00165052 0 0.00165044 0 0.00165054 3.3 0.0016504599999999999 3.3 0.00165056 0 0.00165048 0 0.00165058 3.3 0.0016504999999999998 3.3 0.0016506 0 0.00165052 0 0.00165062 3.3 0.0016505399999999998 3.3 0.0016506399999999999 0 0.00165056 0 0.00165066 3.3 0.00165058 3.3 0.00165068 0 0.0016506 0 0.0016507 3.3 0.00165062 3.3 0.00165072 0 0.0016506399999999999 0 0.00165074 3.3 0.00165066 3.3 0.00165076 0 0.0016506799999999999 0 0.00165078 3.3 0.0016507 3.3 0.0016508 0 0.0016507199999999998 0 0.00165082 3.3 0.00165074 3.3 0.00165084 0 0.0016507599999999998 0 0.0016508599999999999 3.3 0.00165078 3.3 0.00165088 0 0.0016508 0 0.0016509 3.3 0.00165082 3.3 0.00165092 0 0.00165084 0 0.00165094 3.3 0.0016508599999999999 3.3 0.00165096 0 0.00165088 0 0.00165098 3.3 0.0016508999999999999 3.3 0.001651 0 0.00165092 0 0.00165102 3.3 0.0016509399999999998 3.3 0.0016510399999999999 0 0.00165096 0 0.00165106 3.3 0.0016509799999999998 3.3 0.0016510799999999999 0 0.001651 0 0.0016511 3.3 0.00165102 3.3 0.00165112 0 0.0016510399999999999 0 0.00165114 3.3 0.00165106 3.3 0.00165116 0 0.0016510799999999999 0 0.00165118 3.3 0.0016511 3.3 0.0016512 0 0.0016511199999999998 0 0.00165122 3.3 0.00165114 3.3 0.00165124 0 0.0016511599999999998 0 0.0016512599999999999 3.3 0.00165118 3.3 0.00165128 0 0.0016511999999999998 0 0.0016512999999999999 3.3 0.00165122 3.3 0.00165132 0 0.00165124 0 0.00165134 3.3 0.0016512599999999999 3.3 0.00165136 0 0.00165128 0 0.00165138 3.3 0.0016512999999999999 3.3 0.0016514 0 0.00165132 0 0.00165142 3.3 0.0016513399999999998 3.3 0.00165144 0 0.00165136 0 0.00165146 3.3 0.0016513799999999998 3.3 0.0016514799999999999 0 0.0016514 0 0.0016515 3.3 0.00165142 3.3 0.00165152 0 0.00165144 0 0.00165154 3.3 0.00165146 3.3 0.00165156 0 0.0016514799999999999 0 0.00165158 3.3 0.0016515 3.3 0.0016516 0 0.0016515199999999999 0 0.00165162 3.3 0.00165154 3.3 0.00165164 0 0.0016515599999999998 0 0.0016516599999999999 3.3 0.00165158 3.3 0.00165168 0 0.0016515999999999998 0 0.0016516999999999999 3.3 0.00165162 3.3 0.00165172 0 0.00165164 0 0.00165174 3.3 0.0016516599999999999 3.3 0.00165176 0 0.00165168 0 0.00165178 3.3 0.0016516999999999999 3.3 0.0016518 0 0.00165172 0 0.00165182 3.3 0.0016517399999999998 3.3 0.00165184 0 0.00165176 0 0.00165186 3.3 0.0016517799999999998 3.3 0.0016518799999999999 0 0.0016518 0 0.0016519 3.3 0.0016518199999999998 3.3 0.0016519199999999999 0 0.00165184 0 0.00165194 3.3 0.00165186 3.3 0.00165196 0 0.0016518799999999999 0 0.00165198 3.3 0.0016519 3.3 0.001652 0 0.0016519199999999999 0 0.00165202 3.3 0.00165194 3.3 0.00165204 0 0.0016519599999999998 0 0.00165206 3.3 0.00165198 3.3 0.00165208 0 0.0016519999999999998 0 0.0016520999999999999 3.3 0.00165202 3.3 0.00165212 0 0.0016520399999999998 0 0.0016521399999999999 3.3 0.00165206 3.3 0.00165216 0 0.00165208 0 0.00165218 3.3 0.0016520999999999999 3.3 0.0016522 0 0.00165212 0 0.00165222 3.3 0.0016521399999999999 3.3 0.00165224 0 0.00165216 0 0.00165226 3.3 0.0016521799999999998 3.3 0.00165228 0 0.0016522 0 0.0016523 3.3 0.0016522199999999998 3.3 0.0016523199999999999 0 0.00165224 0 0.00165234 3.3 0.00165226 3.3 0.00165236 0 0.00165228 0 0.00165238 3.3 0.0016523 3.3 0.0016524 0 0.0016523199999999999 0 0.00165242 3.3 0.00165234 3.3 0.00165244 0 0.0016523599999999999 0 0.00165246 3.3 0.00165238 3.3 0.00165248 0 0.0016523999999999998 0 0.0016524999999999999 3.3 0.00165242 3.3 0.00165252 0 0.0016524399999999998 0 0.0016525399999999999 3.3 0.00165246 3.3 0.00165256 0 0.00165248 0 0.00165258 3.3 0.0016524999999999999 3.3 0.0016526 0 0.00165252 0 0.00165262 3.3 0.0016525399999999999 3.3 0.00165264 0 0.00165256 0 0.00165266 3.3 0.0016525799999999998 3.3 0.00165268 0 0.0016526 0 0.0016527 3.3 0.0016526199999999998 3.3 0.0016527199999999999 0 0.00165264 0 0.00165274 3.3 0.0016526599999999998 3.3 0.0016527599999999999 0 0.00165268 0 0.00165278 3.3 0.0016527 3.3 0.0016528 0 0.0016527199999999999 0 0.00165282 3.3 0.00165274 3.3 0.00165284 0 0.0016527599999999999 0 0.00165286 3.3 0.00165278 3.3 0.00165288 0 0.0016527999999999998 0 0.0016529 3.3 0.00165282 3.3 0.00165292 0 0.0016528399999999998 0 0.0016529399999999999 3.3 0.00165286 3.3 0.00165296 0 0.00165288 0 0.00165298 3.3 0.0016529 3.3 0.001653 0 0.00165292 0 0.00165302 3.3 0.0016529399999999999 3.3 0.00165304 0 0.00165296 0 0.00165306 3.3 0.0016529799999999999 3.3 0.00165308 0 0.001653 0 0.0016531 3.3 0.0016530199999999998 3.3 0.00165312 0 0.00165304 0 0.00165314 3.3 0.0016530599999999998 3.3 0.0016531599999999999 0 0.00165308 0 0.00165318 3.3 0.0016531 3.3 0.0016532 0 0.00165312 0 0.00165322 3.3 0.00165314 3.3 0.00165324 0 0.0016531599999999999 0 0.00165326 3.3 0.00165318 3.3 0.00165328 0 0.0016531999999999999 0 0.0016533 3.3 0.00165322 3.3 0.00165332 0 0.0016532399999999998 0 0.0016533399999999999 3.3 0.00165326 3.3 0.00165336 0 0.0016532799999999998 0 0.0016533799999999999 3.3 0.0016533 3.3 0.0016534 0 0.00165332 0 0.00165342 3.3 0.0016533399999999999 3.3 0.00165344 0 0.00165336 0 0.00165346 3.3 0.0016533799999999999 3.3 0.00165348 0 0.0016534 0 0.0016535 3.3 0.0016534199999999998 3.3 0.00165352 0 0.00165344 0 0.00165354 3.3 0.0016534599999999998 3.3 0.0016535599999999999 0 0.00165348 0 0.00165358 3.3 0.0016534999999999998 3.3 0.0016535999999999999 0 0.00165352 0 0.00165362 3.3 0.00165354 3.3 0.00165364 0 0.0016535599999999999 0 0.00165366 3.3 0.00165358 3.3 0.00165368 0 0.0016535999999999999 0 0.0016537 3.3 0.00165362 3.3 0.00165372 0 0.0016536399999999998 0 0.00165374 3.3 0.00165366 3.3 0.00165376 0 0.0016536799999999998 0 0.0016537799999999999 3.3 0.0016537 3.3 0.0016538 0 0.00165372 0 0.00165382 3.3 0.00165374 3.3 0.00165384 0 0.00165376 0 0.00165386 3.3 0.0016537799999999999 3.3 0.00165388 0 0.0016538 0 0.0016539 3.3 0.0016538199999999999 3.3 0.00165392 0 0.00165384 0 0.00165394 3.3 0.0016538599999999998 3.3 0.00165396 0 0.00165388 0 0.00165398 3.3 0.0016538999999999998 3.3 0.0016539999999999999 0 0.00165392 0 0.00165402 3.3 0.00165394 3.3 0.00165404 0 0.00165396 0 0.00165406 3.3 0.00165398 3.3 0.00165408 0 0.0016539999999999999 0 0.0016541 3.3 0.00165402 3.3 0.00165412 0 0.0016540399999999999 0 0.00165414 3.3 0.00165406 3.3 0.00165416 0 0.0016540799999999998 0 0.0016541799999999999 3.3 0.0016541 3.3 0.0016542 0 0.0016541199999999998 0 0.0016542199999999999 3.3 0.00165414 3.3 0.00165424 0 0.00165416 0 0.00165426 3.3 0.0016541799999999999 3.3 0.00165428 0 0.0016542 0 0.0016543 3.3 0.0016542199999999999 3.3 0.00165432 0 0.00165424 0 0.00165434 3.3 0.0016542599999999998 3.3 0.00165436 0 0.00165428 0 0.00165438 3.3 0.0016542999999999998 3.3 0.0016543999999999999 0 0.00165432 0 0.00165442 3.3 0.0016543399999999998 3.3 0.0016544399999999999 0 0.00165436 0 0.00165446 3.3 0.00165438 3.3 0.00165448 0 0.0016543999999999999 0 0.0016545 3.3 0.00165442 3.3 0.00165452 0 0.0016544399999999999 0 0.00165454 3.3 0.00165446 3.3 0.00165456 0 0.0016544799999999998 0 0.00165458 3.3 0.0016545 3.3 0.0016546 0 0.0016545199999999998 0 0.0016546199999999999 3.3 0.00165454 3.3 0.00165464 0 0.00165456 0 0.00165466 3.3 0.00165458 3.3 0.00165468 0 0.0016546 0 0.0016547 3.3 0.0016546199999999999 3.3 0.00165472 0 0.00165464 0 0.00165474 3.3 0.0016546599999999999 3.3 0.00165476 0 0.00165468 0 0.00165478 3.3 0.0016546999999999998 3.3 0.0016547999999999999 0 0.00165472 0 0.00165482 3.3 0.0016547399999999998 3.3 0.0016548399999999999 0 0.00165476 0 0.00165486 3.3 0.00165478 3.3 0.00165488 0 0.0016547999999999999 0 0.0016549 3.3 0.00165482 3.3 0.00165492 0 0.0016548399999999999 0 0.00165494 3.3 0.00165486 3.3 0.00165496 0 0.0016548799999999998 0 0.00165498 3.3 0.0016549 3.3 0.001655 0 0.0016549199999999998 0 0.0016550199999999999 3.3 0.00165494 3.3 0.00165504 0 0.0016549599999999998 0 0.0016550599999999999 3.3 0.00165498 3.3 0.00165508 0 0.001655 0 0.0016551 3.3 0.0016550199999999999 3.3 0.00165512 0 0.00165504 0 0.00165514 3.3 0.0016550599999999999 3.3 0.00165516 0 0.00165508 0 0.00165518 3.3 0.0016550999999999998 3.3 0.0016552 0 0.00165512 0 0.00165522 3.3 0.0016551399999999998 3.3 0.0016552399999999999 0 0.00165516 0 0.00165526 3.3 0.0016551799999999998 3.3 0.0016552799999999999 0 0.0016552 0 0.0016553 3.3 0.00165522 3.3 0.00165532 0 0.0016552399999999999 0 0.00165534 3.3 0.00165526 3.3 0.00165536 0 0.0016552799999999999 0 0.00165538 3.3 0.0016553 3.3 0.0016554 0 0.0016553199999999998 0 0.00165542 3.3 0.00165534 3.3 0.00165544 0 0.0016553599999999998 0 0.0016554599999999999 3.3 0.00165538 3.3 0.00165548 0 0.0016554 0 0.0016555 3.3 0.00165542 3.3 0.00165552 0 0.00165544 0 0.00165554 3.3 0.0016554599999999999 3.3 0.00165556 0 0.00165548 0 0.00165558 3.3 0.0016554999999999999 3.3 0.0016556 0 0.00165552 0 0.00165562 3.3 0.0016555399999999998 3.3 0.0016556399999999999 0 0.00165556 0 0.00165566 3.3 0.0016555799999999998 3.3 0.0016556799999999999 0 0.0016556 0 0.0016557 3.3 0.00165562 3.3 0.00165572 0 0.0016556399999999999 0 0.00165574 3.3 0.00165566 3.3 0.00165576 0 0.0016556799999999999 0 0.00165578 3.3 0.0016557 3.3 0.0016558 0 0.0016557199999999998 0 0.00165582 3.3 0.00165574 3.3 0.00165584 0 0.0016557599999999998 0 0.0016558599999999999 3.3 0.00165578 3.3 0.00165588 0 0.0016557999999999998 0 0.0016558999999999999 3.3 0.00165582 3.3 0.00165592 0 0.00165584 0 0.00165594 3.3 0.0016558599999999999 3.3 0.00165596 0 0.00165588 0 0.00165598 3.3 0.0016558999999999999 3.3 0.001656 0 0.00165592 0 0.00165602 3.3 0.0016559399999999998 3.3 0.00165604 0 0.00165596 0 0.00165606 3.3 0.0016559799999999998 3.3 0.0016560799999999999 0 0.001656 0 0.0016561 3.3 0.00165602 3.3 0.00165612 0 0.00165604 0 0.00165614 3.3 0.00165606 3.3 0.00165616 0 0.0016560799999999999 0 0.00165618 3.3 0.0016561 3.3 0.0016562 0 0.0016561199999999999 0 0.00165622 3.3 0.00165614 3.3 0.00165624 0 0.0016561599999999998 0 0.00165626 3.3 0.00165618 3.3 0.00165628 0 0.0016561999999999998 0 0.0016562999999999999 3.3 0.00165622 3.3 0.00165632 0 0.00165624 0 0.00165634 3.3 0.00165626 3.3 0.00165636 0 0.00165628 0 0.00165638 3.3 0.0016562999999999999 3.3 0.0016564 0 0.00165632 0 0.00165642 3.3 0.0016563399999999999 3.3 0.00165644 0 0.00165636 0 0.00165646 3.3 0.0016563799999999998 3.3 0.0016564799999999999 0 0.0016564 0 0.0016565 3.3 0.0016564199999999998 3.3 0.0016565199999999999 0 0.00165644 0 0.00165654 3.3 0.00165646 3.3 0.00165656 0 0.0016564799999999999 0 0.00165658 3.3 0.0016565 3.3 0.0016566 0 0.0016565199999999999 0 0.00165662 3.3 0.00165654 3.3 0.00165664 0 0.0016565599999999998 0 0.00165666 3.3 0.00165658 3.3 0.00165668 0 0.0016565999999999998 0 0.0016566999999999999 3.3 0.00165662 3.3 0.00165672 0 0.0016566399999999998 0 0.0016567399999999999 3.3 0.00165666 3.3 0.00165676 0 0.00165668 0 0.00165678 3.3 0.0016566999999999999 3.3 0.0016568 0 0.00165672 0 0.00165682 3.3 0.0016567399999999999 3.3 0.00165684 0 0.00165676 0 0.00165686 3.3 0.0016567799999999998 3.3 0.00165688 0 0.0016568 0 0.0016569 3.3 0.0016568199999999998 3.3 0.0016569199999999999 0 0.00165684 0 0.00165694 3.3 0.00165686 3.3 0.00165696 0 0.00165688 0 0.00165698 3.3 0.0016569 3.3 0.001657 0 0.0016569199999999999 0 0.00165702 3.3 0.00165694 3.3 0.00165704 0 0.0016569599999999999 0 0.00165706 3.3 0.00165698 3.3 0.00165708 0 0.0016569999999999998 0 0.0016571 3.3 0.00165702 3.3 0.00165712 0 0.0016570399999999998 0 0.0016571399999999999 3.3 0.00165706 3.3 0.00165716 0 0.00165708 0 0.00165718 3.3 0.0016571 3.3 0.0016572 0 0.00165712 0 0.00165722 3.3 0.0016571399999999999 3.3 0.00165724 0 0.00165716 0 0.00165726 3.3 0.0016571799999999999 3.3 0.00165728 0 0.0016572 0 0.0016573 3.3 0.0016572199999999998 3.3 0.0016573199999999999 0 0.00165724 0 0.00165734 3.3 0.0016572599999999998 3.3 0.0016573599999999999 0 0.00165728 0 0.00165738 3.3 0.0016573 3.3 0.0016574 0 0.0016573199999999999 0 0.00165742 3.3 0.00165734 3.3 0.00165744 0 0.0016573599999999999 0 0.00165746 3.3 0.00165738 3.3 0.00165748 0 0.0016573999999999998 0 0.0016575 3.3 0.00165742 3.3 0.00165752 0 0.0016574399999999998 0 0.0016575399999999999 3.3 0.00165746 3.3 0.00165756 0 0.0016574799999999998 0 0.0016575799999999999 3.3 0.0016575 3.3 0.0016576 0 0.00165752 0 0.00165762 3.3 0.0016575399999999999 3.3 0.00165764 0 0.00165756 0 0.00165766 3.3 0.0016575799999999999 3.3 0.00165768 0 0.0016576 0 0.0016577 3.3 0.0016576199999999998 3.3 0.00165772 0 0.00165764 0 0.00165774 3.3 0.0016576599999999998 3.3 0.0016577599999999999 0 0.00165768 0 0.00165778 3.3 0.0016577 3.3 0.0016578 0 0.00165772 0 0.00165782 3.3 0.00165774 3.3 0.00165784 0 0.0016577599999999999 0 0.00165786 3.3 0.00165778 3.3 0.00165788 0 0.0016577999999999999 0 0.0016579 3.3 0.00165782 3.3 0.00165792 0 0.0016578399999999998 0 0.0016579399999999999 3.3 0.00165786 3.3 0.00165796 0 0.0016578799999999998 0 0.0016579799999999999 3.3 0.0016579 3.3 0.001658 0 0.00165792 0 0.00165802 3.3 0.0016579399999999999 3.3 0.00165804 0 0.00165796 0 0.00165806 3.3 0.0016579799999999999 3.3 0.00165808 0 0.001658 0 0.0016581 3.3 0.0016580199999999998 3.3 0.00165812 0 0.00165804 0 0.00165814 3.3 0.0016580599999999998 3.3 0.0016581599999999999 0 0.00165808 0 0.00165818 3.3 0.0016580999999999998 3.3 0.0016581999999999999 0 0.00165812 0 0.00165822 3.3 0.00165814 3.3 0.00165824 0 0.0016581599999999999 0 0.00165826 3.3 0.00165818 3.3 0.00165828 0 0.0016581999999999999 0 0.0016583 3.3 0.00165822 3.3 0.00165832 0 0.0016582399999999998 0 0.00165834 3.3 0.00165826 3.3 0.00165836 0 0.0016582799999999998 0 0.0016583799999999999 3.3 0.0016583 3.3 0.0016584 0 0.0016583199999999998 0 0.0016584199999999999 3.3 0.00165834 3.3 0.00165844 0 0.00165836 0 0.00165846 3.3 0.0016583799999999999 3.3 0.00165848 0 0.0016584 0 0.0016585 3.3 0.0016584199999999999 3.3 0.00165852 0 0.00165844 0 0.00165854 3.3 0.0016584599999999998 3.3 0.00165856 0 0.00165848 0 0.00165858 3.3 0.0016584999999999998 3.3 0.0016585999999999999 0 0.00165852 0 0.00165862 3.3 0.00165854 3.3 0.00165864 0 0.00165856 0 0.00165866 3.3 0.00165858 3.3 0.00165868 0 0.0016585999999999999 0 0.0016587 3.3 0.00165862 3.3 0.00165872 0 0.0016586399999999999 0 0.00165874 3.3 0.00165866 3.3 0.00165876 0 0.0016586799999999998 0 0.0016587799999999999 3.3 0.0016587 3.3 0.0016588 0 0.0016587199999999998 0 0.0016588199999999999 3.3 0.00165874 3.3 0.00165884 0 0.00165876 0 0.00165886 3.3 0.0016587799999999999 3.3 0.00165888 0 0.0016588 0 0.0016589 3.3 0.0016588199999999999 3.3 0.00165892 0 0.00165884 0 0.00165894 3.3 0.0016588599999999998 3.3 0.00165896 0 0.00165888 0 0.00165898 3.3 0.0016588999999999998 3.3 0.0016589999999999999 0 0.00165892 0 0.00165902 3.3 0.0016589399999999998 3.3 0.0016590399999999999 0 0.00165896 0 0.00165906 3.3 0.00165898 3.3 0.00165908 0 0.0016589999999999999 0 0.0016591 3.3 0.00165902 3.3 0.00165912 0 0.0016590399999999999 0 0.00165914 3.3 0.00165906 3.3 0.00165916 0 0.0016590799999999998 0 0.00165918 3.3 0.0016591 3.3 0.0016592 0 0.0016591199999999998 0 0.0016592199999999999 3.3 0.00165914 3.3 0.00165924 0 0.0016591599999999998 0 0.0016592599999999999 3.3 0.00165918 3.3 0.00165928 0 0.0016592 0 0.0016593 3.3 0.0016592199999999999 3.3 0.00165932 0 0.00165924 0 0.00165934 3.3 0.0016592599999999999 3.3 0.00165936 0 0.00165928 0 0.00165938 3.3 0.0016592999999999998 3.3 0.0016594 0 0.00165932 0 0.00165942 3.3 0.0016593399999999998 3.3 0.0016594399999999999 0 0.00165936 0 0.00165946 3.3 0.00165938 3.3 0.00165948 0 0.0016594 0 0.0016595 3.3 0.00165942 3.3 0.00165952 0 0.0016594399999999999 0 0.00165954 3.3 0.00165946 3.3 0.00165956 0 0.0016594799999999999 0 0.00165958 3.3 0.0016595 3.3 0.0016596 0 0.0016595199999999998 0 0.0016596199999999999 3.3 0.00165954 3.3 0.00165964 0 0.0016595599999999998 0 0.0016596599999999999 3.3 0.00165958 3.3 0.00165968 0 0.0016596 0 0.0016597 3.3 0.0016596199999999999 3.3 0.00165972 0 0.00165964 0 0.00165974 3.3 0.0016596599999999999 3.3 0.00165976 0 0.00165968 0 0.00165978 3.3 0.0016596999999999998 3.3 0.0016598 0 0.00165972 0 0.00165982 3.3 0.0016597399999999998 3.3 0.0016598399999999999 0 0.00165976 0 0.00165986 3.3 0.0016597799999999998 3.3 0.0016598799999999999 0 0.0016598 0 0.0016599 3.3 0.00165982 3.3 0.00165992 0 0.0016598399999999999 0 0.00165994 3.3 0.00165986 3.3 0.00165996 0 0.0016598799999999999 0 0.00165998 3.3 0.0016599 3.3 0.00166 0 0.0016599199999999998 0 0.00166002 3.3 0.00165994 3.3 0.00166004 0 0.0016599599999999998 0 0.0016600599999999999 3.3 0.00165998 3.3 0.00166008 0 0.00166 0 0.0016601 3.3 0.00166002 3.3 0.00166012 0 0.00166004 0 0.00166014 3.3 0.0016600599999999999 3.3 0.00166016 0 0.00166008 0 0.00166018 3.3 0.0016600999999999999 3.3 0.0016602 0 0.00166012 0 0.00166022 3.3 0.0016601399999999998 3.3 0.00166024 0 0.00166016 0 0.00166026 3.3 0.0016601799999999998 3.3 0.0016602799999999999 0 0.0016602 0 0.0016603 3.3 0.00166022 3.3 0.00166032 0 0.00166024 0 0.00166034 3.3 0.00166026 3.3 0.00166036 0 0.0016602799999999999 0 0.00166038 3.3 0.0016603 3.3 0.0016604 0 0.0016603199999999999 0 0.00166042 3.3 0.00166034 3.3 0.00166044 0 0.0016603599999999998 0 0.0016604599999999999 3.3 0.00166038 3.3 0.00166048 0 0.0016603999999999998 0 0.0016604999999999999 3.3 0.00166042 3.3 0.00166052 0 0.00166044 0 0.00166054 3.3 0.0016604599999999999 3.3 0.00166056 0 0.00166048 0 0.00166058 3.3 0.0016604999999999999 3.3 0.0016606 0 0.00166052 0 0.00166062 3.3 0.0016605399999999998 3.3 0.00166064 0 0.00166056 0 0.00166066 3.3 0.0016605799999999998 3.3 0.0016606799999999999 0 0.0016606 0 0.0016607 3.3 0.0016606199999999998 3.3 0.0016607199999999999 0 0.00166064 0 0.00166074 3.3 0.00166066 3.3 0.00166076 0 0.0016606799999999999 0 0.00166078 3.3 0.0016607 3.3 0.0016608 0 0.0016607199999999999 0 0.00166082 3.3 0.00166074 3.3 0.00166084 0 0.0016607599999999998 0 0.00166086 3.3 0.00166078 3.3 0.00166088 0 0.0016607999999999998 0 0.0016608999999999999 3.3 0.00166082 3.3 0.00166092 0 0.00166084 0 0.00166094 3.3 0.00166086 3.3 0.00166096 0 0.00166088 0 0.00166098 3.3 0.0016608999999999999 3.3 0.001661 0 0.00166092 0 0.00166102 3.3 0.0016609399999999999 3.3 0.00166104 0 0.00166096 0 0.00166106 3.3 0.0016609799999999998 3.3 0.00166108 0 0.001661 0 0.0016611 3.3 0.0016610199999999998 3.3 0.0016611199999999999 0 0.00166104 0 0.00166114 3.3 0.00166106 3.3 0.00166116 0 0.00166108 0 0.00166118 3.3 0.0016611 3.3 0.0016612 0 0.0016611199999999999 0 0.00166122 3.3 0.00166114 3.3 0.00166124 0 0.0016611599999999999 0 0.00166126 3.3 0.00166118 3.3 0.00166128 0 0.0016611999999999998 0 0.0016612999999999999 3.3 0.00166122 3.3 0.00166132 0 0.0016612399999999998 0 0.0016613399999999999 3.3 0.00166126 3.3 0.00166136 0 0.00166128 0 0.00166138 3.3 0.0016612999999999999 3.3 0.0016614 0 0.00166132 0 0.00166142 3.3 0.0016613399999999999 3.3 0.00166144 0 0.00166136 0 0.00166146 3.3 0.0016613799999999998 3.3 0.00166148 0 0.0016614 0 0.0016615 3.3 0.0016614199999999998 3.3 0.0016615199999999999 0 0.00166144 0 0.00166154 3.3 0.0016614599999999998 3.3 0.0016615599999999999 0 0.00166148 0 0.00166158 3.3 0.0016615 3.3 0.0016616 0 0.0016615199999999999 0 0.00166162 3.3 0.00166154 3.3 0.00166164 0 0.0016615599999999999 0 0.00166166 3.3 0.00166158 3.3 0.00166168 0 0.0016615999999999998 0 0.0016617 3.3 0.00166162 3.3 0.00166172 0 0.0016616399999999998 0 0.0016617399999999999 3.3 0.00166166 3.3 0.00166176 0 0.00166168 0 0.00166178 3.3 0.0016617 3.3 0.0016618 0 0.00166172 0 0.00166182 3.3 0.0016617399999999999 3.3 0.00166184 0 0.00166176 0 0.00166186 3.3 0.0016617799999999999 3.3 0.00166188 0 0.0016618 0 0.0016619 3.3 0.0016618199999999998 3.3 0.0016619199999999999 0 0.00166184 0 0.00166194 3.3 0.0016618599999999998 3.3 0.0016619599999999999 0 0.00166188 0 0.00166198 3.3 0.0016619 3.3 0.001662 0 0.0016619199999999999 0 0.00166202 3.3 0.00166194 3.3 0.00166204 0 0.0016619599999999999 0 0.00166206 3.3 0.00166198 3.3 0.00166208 0 0.0016619999999999998 0 0.0016621 3.3 0.00166202 3.3 0.00166212 0 0.0016620399999999998 0 0.0016621399999999999 3.3 0.00166206 3.3 0.00166216 0 0.0016620799999999998 0 0.0016621799999999999 3.3 0.0016621 3.3 0.0016622 0 0.00166212 0 0.00166222 3.3 0.0016621399999999999 3.3 0.00166224 0 0.00166216 0 0.00166226 3.3 0.0016621799999999999 3.3 0.00166228 0 0.0016622 0 0.0016623 3.3 0.0016622199999999998 3.3 0.00166232 0 0.00166224 0 0.00166234 3.3 0.0016622599999999998 3.3 0.0016623599999999999 0 0.00166228 0 0.00166238 3.3 0.0016622999999999998 3.3 0.0016623999999999999 0 0.00166232 0 0.00166242 3.3 0.00166234 3.3 0.00166244 0 0.0016623599999999999 0 0.00166246 3.3 0.00166238 3.3 0.00166248 0 0.0016623999999999999 0 0.0016625 3.3 0.00166242 3.3 0.00166252 0 0.0016624399999999998 0 0.00166254 3.3 0.00166246 3.3 0.00166256 0 0.0016624799999999998 0 0.0016625799999999999 3.3 0.0016625 3.3 0.0016626 0 0.00166252 0 0.00166262 3.3 0.00166254 3.3 0.00166264 0 0.00166256 0 0.00166266 3.3 0.0016625799999999999 3.3 0.00166268 0 0.0016626 0 0.0016627 3.3 0.0016626199999999999 3.3 0.00166272 0 0.00166264 0 0.00166274 3.3 0.0016626599999999998 3.3 0.0016627599999999999 0 0.00166268 0 0.00166278 3.3 0.0016626999999999998 3.3 0.0016627999999999999 0 0.00166272 0 0.00166282 3.3 0.00166274 3.3 0.00166284 0 0.0016627599999999999 0 0.00166286 3.3 0.00166278 3.3 0.00166288 0 0.0016627999999999999 0 0.0016629 3.3 0.00166282 3.3 0.00166292 0 0.0016628399999999998 0 0.00166294 3.3 0.00166286 3.3 0.00166296 0 0.0016628799999999998 0 0.0016629799999999999 3.3 0.0016629 3.3 0.001663 0 0.0016629199999999998 0 0.0016630199999999999 3.3 0.00166294 3.3 0.00166304 0 0.00166296 0 0.00166306 3.3 0.0016629799999999999 3.3 0.00166308 0 0.001663 0 0.0016631 3.3 0.0016630199999999999 3.3 0.00166312 0 0.00166304 0 0.00166314 3.3 0.0016630599999999998 3.3 0.00166316 0 0.00166308 0 0.00166318 3.3 0.0016630999999999998 3.3 0.0016631999999999999 0 0.00166312 0 0.00166322 3.3 0.00166314 3.3 0.00166324 0 0.00166316 0 0.00166326 3.3 0.00166318 3.3 0.00166328 0 0.0016631999999999999 0 0.0016633 3.3 0.00166322 3.3 0.00166332 0 0.0016632399999999999 0 0.00166334 3.3 0.00166326 3.3 0.00166336 0 0.0016632799999999998 0 0.00166338 3.3 0.0016633 3.3 0.0016634 0 0.0016633199999999998 0 0.0016634199999999999 3.3 0.00166334 3.3 0.00166344 0 0.00166336 0 0.00166346 3.3 0.00166338 3.3 0.00166348 0 0.0016634 0 0.0016635 3.3 0.0016634199999999999 3.3 0.00166352 0 0.00166344 0 0.00166354 3.3 0.0016634599999999999 3.3 0.00166356 0 0.00166348 0 0.00166358 3.3 0.0016634999999999998 3.3 0.0016635999999999999 0 0.00166352 0 0.00166362 3.3 0.0016635399999999998 3.3 0.0016636399999999999 0 0.00166356 0 0.00166366 3.3 0.00166358 3.3 0.00166368 0 0.0016635999999999999 0 0.0016637 3.3 0.00166362 3.3 0.00166372 0 0.0016636399999999999 0 0.00166374 3.3 0.00166366 3.3 0.00166376 0 0.0016636799999999998 0 0.00166378 3.3 0.0016637 3.3 0.0016638 0 0.0016637199999999998 0 0.0016638199999999999 3.3 0.00166374 3.3 0.00166384 0 0.0016637599999999998 0 0.0016638599999999999 3.3 0.00166378 3.3 0.00166388 0 0.0016638 0 0.0016639 3.3 0.0016638199999999999 3.3 0.00166392 0 0.00166384 0 0.00166394 3.3 0.0016638599999999999 3.3 0.00166396 0 0.00166388 0 0.00166398 3.3 0.0016638999999999998 3.3 0.001664 0 0.00166392 0 0.00166402 3.3 0.0016639399999999998 3.3 0.0016640399999999999 0 0.00166396 0 0.00166406 3.3 0.00166398 3.3 0.00166408 0 0.001664 0 0.0016641 3.3 0.00166402 3.3 0.00166412 0 0.0016640399999999999 0 0.00166414 3.3 0.00166406 3.3 0.00166416 0 0.0016640799999999999 0 0.00166418 3.3 0.0016641 3.3 0.0016642 0 0.0016641199999999998 0 0.00166422 3.3 0.00166414 3.3 0.00166424 0 0.0016641599999999998 0 0.0016642599999999999 3.3 0.00166418 3.3 0.00166428 0 0.0016642 0 0.0016643 3.3 0.00166422 3.3 0.00166432 0 0.00166424 0 0.00166434 3.3 0.0016642599999999999 3.3 0.00166436 0 0.00166428 0 0.00166438 3.3 0.0016642999999999999 3.3 0.0016644 0 0.00166432 0 0.00166442 3.3 0.0016643399999999998 3.3 0.0016644399999999999 0 0.00166436 0 0.00166446 3.3 0.0016643799999999998 3.3 0.0016644799999999999 0 0.0016644 0 0.0016645 3.3 0.00166442 3.3 0.00166452 0 0.0016644399999999999 0 0.00166454 3.3 0.00166446 3.3 0.00166456 0 0.0016644799999999999 0 0.00166458 3.3 0.0016645 3.3 0.0016646 0 0.0016645199999999998 0 0.00166462 3.3 0.00166454 3.3 0.00166464 0 0.0016645599999999998 0 0.0016646599999999999 3.3 0.00166458 3.3 0.00166468 0 0.0016645999999999998 0 0.0016646999999999999 3.3 0.00166462 3.3 0.00166472 0 0.00166464 0 0.00166474 3.3 0.0016646599999999999 3.3 0.00166476 0 0.00166468 0 0.00166478 3.3 0.0016646999999999999 3.3 0.0016648 0 0.00166472 0 0.00166482 3.3 0.0016647399999999998 3.3 0.00166484 0 0.00166476 0 0.00166486 3.3 0.0016647799999999998 3.3 0.0016648799999999999 0 0.0016648 0 0.0016649 3.3 0.00166482 3.3 0.00166492 0 0.00166484 0 0.00166494 3.3 0.00166486 3.3 0.00166496 0 0.0016648799999999999 0 0.00166498 3.3 0.0016649 3.3 0.001665 0 0.0016649199999999999 0 0.00166502 3.3 0.00166494 3.3 0.00166504 0 0.0016649599999999998 0 0.0016650599999999999 3.3 0.00166498 3.3 0.00166508 0 0.0016649999999999998 0 0.0016650999999999999 3.3 0.00166502 3.3 0.00166512 0 0.00166504 0 0.00166514 3.3 0.0016650599999999999 3.3 0.00166516 0 0.00166508 0 0.00166518 3.3 0.0016650999999999999 3.3 0.0016652 0 0.00166512 0 0.00166522 3.3 0.0016651399999999998 3.3 0.00166524 0 0.00166516 0 0.00166526 3.3 0.0016651799999999998 3.3 0.0016652799999999999 0 0.0016652 0 0.0016653 3.3 0.0016652199999999998 3.3 0.0016653199999999999 0 0.00166524 0 0.00166534 3.3 0.00166526 3.3 0.00166536 0 0.0016652799999999999 0 0.00166538 3.3 0.0016653 3.3 0.0016654 0 0.0016653199999999999 0 0.00166542 3.3 0.00166534 3.3 0.00166544 0 0.0016653599999999998 0 0.00166546 3.3 0.00166538 3.3 0.00166548 0 0.0016653999999999998 0 0.0016654999999999999 3.3 0.00166542 3.3 0.00166552 0 0.0016654399999999998 0 0.0016655399999999999 3.3 0.00166546 3.3 0.00166556 0 0.00166548 0 0.00166558 3.3 0.0016654999999999999 3.3 0.0016656 0 0.00166552 0 0.00166562 3.3 0.0016655399999999999 3.3 0.00166564 0 0.00166556 0 0.00166566 3.3 0.0016655799999999998 3.3 0.00166568 0 0.0016656 0 0.0016657 3.3 0.0016656199999999998 3.3 0.0016657199999999999 0 0.00166564 0 0.00166574 3.3 0.00166566 3.3 0.00166576 0 0.00166568 0 0.00166578 3.3 0.0016657 3.3 0.0016658 0 0.0016657199999999999 0 0.00166582 3.3 0.00166574 3.3 0.00166584 0 0.0016657599999999999 0 0.00166586 3.3 0.00166578 3.3 0.00166588 0 0.0016657999999999998 0 0.0016658999999999999 3.3 0.00166582 3.3 0.00166592 0 0.0016658399999999998 0 0.0016659399999999999 3.3 0.00166586 3.3 0.00166596 0 0.00166588 0 0.00166598 3.3 0.0016658999999999999 3.3 0.001666 0 0.00166592 0 0.00166602 3.3 0.0016659399999999999 3.3 0.00166604 0 0.00166596 0 0.00166606 3.3 0.0016659799999999998 3.3 0.00166608 0 0.001666 0 0.0016661 3.3 0.0016660199999999998 3.3 0.0016661199999999999 0 0.00166604 0 0.00166614 3.3 0.0016660599999999998 3.3 0.0016661599999999999 0 0.00166608 0 0.00166618 3.3 0.0016661 3.3 0.0016662 0 0.0016661199999999999 0 0.00166622 3.3 0.00166614 3.3 0.00166624 0 0.0016661599999999999 0 0.00166626 3.3 0.00166618 3.3 0.00166628 0 0.0016661999999999998 0 0.0016663 3.3 0.00166622 3.3 0.00166632 0 0.0016662399999999998 0 0.0016663399999999999 3.3 0.00166626 3.3 0.00166636 0 0.00166628 0 0.00166638 3.3 0.0016663 3.3 0.0016664 0 0.00166632 0 0.00166642 3.3 0.0016663399999999999 3.3 0.00166644 0 0.00166636 0 0.00166646 3.3 0.0016663799999999999 3.3 0.00166648 0 0.0016664 0 0.0016665 3.3 0.0016664199999999998 3.3 0.00166652 0 0.00166644 0 0.00166654 3.3 0.0016664599999999998 3.3 0.0016665599999999999 0 0.00166648 0 0.00166658 3.3 0.0016665 3.3 0.0016666 0 0.00166652 0 0.00166662 3.3 0.00166654 3.3 0.00166664 0 0.0016665599999999999 0 0.00166666 3.3 0.00166658 3.3 0.00166668 0 0.0016665999999999999 0 0.0016667 3.3 0.00166662 3.3 0.00166672 0 0.0016666399999999998 0 0.0016667399999999999 3.3 0.00166666 3.3 0.00166676 0 0.0016666799999999998 0 0.0016667799999999999 3.3 0.0016667 3.3 0.0016668 0 0.00166672 0 0.00166682 3.3 0.0016667399999999999 3.3 0.00166684 0 0.00166676 0 0.00166686 3.3 0.0016667799999999999 3.3 0.00166688 0 0.0016668 0 0.0016669 3.3 0.0016668199999999998 3.3 0.00166692 0 0.00166684 0 0.00166694 3.3 0.0016668599999999998 3.3 0.0016669599999999999 0 0.00166688 0 0.00166698 3.3 0.0016668999999999998 3.3 0.0016669999999999999 0 0.00166692 0 0.00166702 3.3 0.00166694 3.3 0.00166704 0 0.0016669599999999999 0 0.00166706 3.3 0.00166698 3.3 0.00166708 0 0.0016669999999999999 0 0.0016671 3.3 0.00166702 3.3 0.00166712 0 0.0016670399999999998 0 0.00166714 3.3 0.00166706 3.3 0.00166716 0 0.0016670799999999998 0 0.0016671799999999999 3.3 0.0016671 3.3 0.0016672 0 0.00166712 0 0.00166722 3.3 0.00166714 3.3 0.00166724 0 0.00166716 0 0.00166726 3.3 0.0016671799999999999 3.3 0.00166728 0 0.0016672 0 0.0016673 3.3 0.0016672199999999999 3.3 0.00166732 0 0.00166724 0 0.00166734 3.3 0.0016672599999999998 3.3 0.00166736 0 0.00166728 0 0.00166738 3.3 0.0016672999999999998 3.3 0.0016673999999999999 0 0.00166732 0 0.00166742 3.3 0.00166734 3.3 0.00166744 0 0.00166736 0 0.00166746 3.3 0.00166738 3.3 0.00166748 0 0.0016673999999999999 0 0.0016675 3.3 0.00166742 3.3 0.00166752 0 0.0016674399999999999 0 0.00166754 3.3 0.00166746 3.3 0.00166756 0 0.0016674799999999998 0 0.0016675799999999999 3.3 0.0016675 3.3 0.0016676 0 0.0016675199999999998 0 0.0016676199999999999 3.3 0.00166754 3.3 0.00166764 0 0.00166756 0 0.00166766 3.3 0.0016675799999999999 3.3 0.00166768 0 0.0016676 0 0.0016677 3.3 0.0016676199999999999 3.3 0.00166772 0 0.00166764 0 0.00166774 3.3 0.0016676599999999998 3.3 0.00166776 0 0.00166768 0 0.00166778 3.3 0.0016676999999999998 3.3 0.0016677999999999999 0 0.00166772 0 0.00166782 3.3 0.0016677399999999998 3.3 0.0016678399999999999 0 0.00166776 0 0.00166786 3.3 0.00166778 3.3 0.00166788 0 0.0016677999999999999 0 0.0016679 3.3 0.00166782 3.3 0.00166792 0 0.0016678399999999999 0 0.00166794 3.3 0.00166786 3.3 0.00166796 0 0.0016678799999999998 0 0.00166798 3.3 0.0016679 3.3 0.001668 0 0.0016679199999999998 0 0.0016680199999999999 3.3 0.00166794 3.3 0.00166804 0 0.00166796 0 0.00166806 3.3 0.00166798 3.3 0.00166808 0 0.001668 0 0.0016681 3.3 0.0016680199999999999 3.3 0.00166812 0 0.00166804 0 0.00166814 3.3 0.0016680599999999999 3.3 0.00166816 0 0.00166808 0 0.00166818 3.3 0.0016680999999999998 3.3 0.0016681999999999999 0 0.00166812 0 0.00166822 3.3 0.0016681399999999998 3.3 0.0016682399999999999 0 0.00166816 0 0.00166826 3.3 0.00166818 3.3 0.00166828 0 0.0016681999999999999 0 0.0016683 3.3 0.00166822 3.3 0.00166832 0 0.0016682399999999999 0 0.00166834 3.3 0.00166826 3.3 0.00166836 0 0.0016682799999999998 0 0.00166838 3.3 0.0016683 3.3 0.0016684 0 0.0016683199999999998 0 0.0016684199999999999 3.3 0.00166834 3.3 0.00166844 0 0.0016683599999999998 0 0.0016684599999999999 3.3 0.00166838 3.3 0.00166848 0 0.0016684 0 0.0016685 3.3 0.0016684199999999999 3.3 0.00166852 0 0.00166844 0 0.00166854 3.3 0.0016684599999999999 3.3 0.00166856 0 0.00166848 0 0.00166858 3.3 0.0016684999999999998 3.3 0.0016686 0 0.00166852 0 0.00166862 3.3 0.0016685399999999998 3.3 0.0016686399999999999 0 0.00166856 0 0.00166866 3.3 0.0016685799999999998 3.3 0.0016686799999999999 0 0.0016686 0 0.0016687 3.3 0.00166862 3.3 0.00166872 0 0.0016686399999999999 0 0.00166874 3.3 0.00166866 3.3 0.00166876 0 0.0016686799999999999 0 0.00166878 3.3 0.0016687 3.3 0.0016688 0 0.0016687199999999998 0 0.00166882 3.3 0.00166874 3.3 0.00166884 0 0.0016687599999999998 0 0.0016688599999999999 3.3 0.00166878 3.3 0.00166888 0 0.0016688 0 0.0016689 3.3 0.00166882 3.3 0.00166892 0 0.00166884 0 0.00166894 3.3 0.0016688599999999999 3.3 0.00166896 0 0.00166888 0 0.00166898 3.3 0.0016688999999999999 3.3 0.001669 0 0.00166892 0 0.00166902 3.3 0.0016689399999999998 3.3 0.0016690399999999999 0 0.00166896 0 0.00166906 3.3 0.0016689799999999998 3.3 0.0016690799999999999 0 0.001669 0 0.0016691 3.3 0.00166902 3.3 0.00166912 0 0.0016690399999999999 0 0.00166914 3.3 0.00166906 3.3 0.00166916 0 0.0016690799999999999 0 0.00166918 3.3 0.0016691 3.3 0.0016692 0 0.0016691199999999998 0 0.00166922 3.3 0.00166914 3.3 0.00166924 0 0.0016691599999999998 0 0.0016692599999999999 3.3 0.00166918 3.3 0.00166928 0 0.0016691999999999998 0 0.0016692999999999999 3.3 0.00166922 3.3 0.00166932 0 0.00166924 0 0.00166934 3.3 0.0016692599999999999 3.3 0.00166936 0 0.00166928 0 0.00166938 3.3 0.0016692999999999999 3.3 0.0016694 0 0.00166932 0 0.00166942 3.3 0.0016693399999999998 3.3 0.00166944 0 0.00166936 0 0.00166946 3.3 0.0016693799999999998 3.3 0.0016694799999999999 0 0.0016694 0 0.0016695 3.3 0.0016694199999999998 3.3 0.0016695199999999999 0 0.00166944 0 0.00166954 3.3 0.00166946 3.3 0.00166956 0 0.0016694799999999999 0 0.00166958 3.3 0.0016695 3.3 0.0016696 0 0.0016695199999999999 0 0.00166962 3.3 0.00166954 3.3 0.00166964 0 0.0016695599999999998 0 0.00166966 3.3 0.00166958 3.3 0.00166968 0 0.0016695999999999998 0 0.0016696999999999999 3.3 0.00166962 3.3 0.00166972 0 0.00166964 0 0.00166974 3.3 0.00166966 3.3 0.00166976 0 0.00166968 0 0.00166978 3.3 0.0016696999999999999 3.3 0.0016698 0 0.00166972 0 0.00166982 3.3 0.0016697399999999999 3.3 0.00166984 0 0.00166976 0 0.00166986 3.3 0.0016697799999999998 3.3 0.0016698799999999999 0 0.0016698 0 0.0016699 3.3 0.0016698199999999998 3.3 0.0016699199999999999 0 0.00166984 0 0.00166994 3.3 0.00166986 3.3 0.00166996 0 0.0016698799999999999 0 0.00166998 3.3 0.0016699 3.3 0.00167 0 0.0016699199999999999 0 0.00167002 3.3 0.00166994 3.3 0.00167004 0 0.0016699599999999998 0 0.00167006 3.3 0.00166998 3.3 0.00167008 0 0.0016699999999999998 0 0.0016700999999999999 3.3 0.00167002 3.3 0.00167012 0 0.0016700399999999998 0 0.0016701399999999999 3.3 0.00167006 3.3 0.00167016 0 0.00167008 0 0.00167018 3.3 0.0016700999999999999 3.3 0.0016702 0 0.00167012 0 0.00167022 3.3 0.0016701399999999999 3.3 0.00167024 0 0.00167016 0 0.00167026 3.3 0.0016701799999999998 3.3 0.00167028 0 0.0016702 0 0.0016703 3.3 0.0016702199999999998 3.3 0.0016703199999999999 0 0.00167024 0 0.00167034 3.3 0.00167026 3.3 0.00167036 0 0.00167028 0 0.00167038 3.3 0.0016703 3.3 0.0016704 0 0.0016703199999999999 0 0.00167042 3.3 0.00167034 3.3 0.00167044 0 0.0016703599999999999 0 0.00167046 3.3 0.00167038 3.3 0.00167048 0 0.0016703999999999998 0 0.0016705 3.3 0.00167042 3.3 0.00167052 0 0.0016704399999999998 0 0.0016705399999999999 3.3 0.00167046 3.3 0.00167056 0 0.00167048 0 0.00167058 3.3 0.0016705 3.3 0.0016706 0 0.00167052 0 0.00167062 3.3 0.0016705399999999999 3.3 0.00167064 0 0.00167056 0 0.00167066 3.3 0.0016705799999999999 3.3 0.00167068 0 0.0016706 0 0.0016707 3.3 0.0016706199999999998 3.3 0.0016707199999999999 0 0.00167064 0 0.00167074 3.3 0.0016706599999999998 3.3 0.0016707599999999999 0 0.00167068 0 0.00167078 3.3 0.0016707 3.3 0.0016708 0 0.0016707199999999999 0 0.00167082 3.3 0.00167074 3.3 0.00167084 0 0.0016707599999999999 0 0.00167086 3.3 0.00167078 3.3 0.00167088 0 0.0016707999999999998 0 0.0016709 3.3 0.00167082 3.3 0.00167092 0 0.0016708399999999998 0 0.0016709399999999999 3.3 0.00167086 3.3 0.00167096 0 0.0016708799999999998 0 0.0016709799999999999 3.3 0.0016709 3.3 0.001671 0 0.00167092 0 0.00167102 3.3 0.0016709399999999999 3.3 0.00167104 0 0.00167096 0 0.00167106 3.3 0.0016709799999999999 3.3 0.00167108 0 0.001671 0 0.0016711 3.3 0.0016710199999999998 3.3 0.00167112 0 0.00167104 0 0.00167114 3.3 0.0016710599999999998 3.3 0.0016711599999999999 0 0.00167108 0 0.00167118 3.3 0.0016711 3.3 0.0016712 0 0.00167112 0 0.00167122 3.3 0.00167114 3.3 0.00167124 0 0.0016711599999999999 0 0.00167126 3.3 0.00167118 3.3 0.00167128 0 0.0016711999999999999 0 0.0016713 3.3 0.00167122 3.3 0.00167132 0 0.0016712399999999998 0 0.00167134 3.3 0.00167126 3.3 0.00167136 0 0.0016712799999999998 0 0.0016713799999999999 3.3 0.0016713 3.3 0.0016714 0 0.00167132 0 0.00167142 3.3 0.00167134 3.3 0.00167144 0 0.00167136 0 0.00167146 3.3 0.0016713799999999999 3.3 0.00167148 0 0.0016714 0 0.0016715 3.3 0.0016714199999999999 3.3 0.00167152 0 0.00167144 0 0.00167154 3.3 0.0016714599999999998 3.3 0.0016715599999999999 0 0.00167148 0 0.00167158 3.3 0.0016714999999999998 3.3 0.0016715999999999999 0 0.00167152 0 0.00167162 3.3 0.00167154 3.3 0.00167164 0 0.0016715599999999999 0 0.00167166 3.3 0.00167158 3.3 0.00167168 0 0.0016715999999999999 0 0.0016717 3.3 0.00167162 3.3 0.00167172 0 0.0016716399999999998 0 0.00167174 3.3 0.00167166 3.3 0.00167176 0 0.0016716799999999998 0 0.0016717799999999999 3.3 0.0016717 3.3 0.0016718 0 0.0016717199999999998 0 0.0016718199999999999 3.3 0.00167174 3.3 0.00167184 0 0.00167176 0 0.00167186 3.3 0.0016717799999999999 3.3 0.00167188 0 0.0016718 0 0.0016719 3.3 0.0016718199999999999 3.3 0.00167192 0 0.00167184 0 0.00167194 3.3 0.0016718599999999998 3.3 0.00167196 0 0.00167188 0 0.00167198 3.3 0.0016718999999999998 3.3 0.0016719999999999999 0 0.00167192 0 0.00167202 3.3 0.00167194 3.3 0.00167204 0 0.00167196 0 0.00167206 3.3 0.00167198 3.3 0.00167208 0 0.0016719999999999999 0 0.0016721 3.3 0.00167202 3.3 0.00167212 0 0.0016720399999999999 0 0.00167214 3.3 0.00167206 3.3 0.00167216 0 0.0016720799999999998 0 0.0016721799999999999 3.3 0.0016721 3.3 0.0016722 0 0.0016721199999999998 0 0.0016722199999999999 3.3 0.00167214 3.3 0.00167224 0 0.00167216 0 0.00167226 3.3 0.0016721799999999999 3.3 0.00167228 0 0.0016722 0 0.0016723 3.3 0.0016722199999999999 3.3 0.00167232 0 0.00167224 0 0.00167234 3.3 0.0016722599999999998 3.3 0.00167236 0 0.00167228 0 0.00167238 3.3 0.0016722999999999998 3.3 0.0016723999999999999 0 0.00167232 0 0.00167242 3.3 0.0016723399999999998 3.3 0.0016724399999999999 0 0.00167236 0 0.00167246 3.3 0.00167238 3.3 0.00167248 0 0.0016723999999999999 0 0.0016725 3.3 0.00167242 3.3 0.00167252 0 0.0016724399999999999 0 0.00167254 3.3 0.00167246 3.3 0.00167256 0 0.0016724799999999998 0 0.00167258 3.3 0.0016725 3.3 0.0016726 0 0.0016725199999999998 0 0.0016726199999999999 3.3 0.00167254 3.3 0.00167264 0 0.0016725599999999998 0 0.0016726599999999999 3.3 0.00167258 3.3 0.00167268 0 0.0016726 0 0.0016727 3.3 0.0016726199999999999 3.3 0.00167272 0 0.00167264 0 0.00167274 3.3 0.0016726599999999999 3.3 0.00167276 0 0.00167268 0 0.00167278 3.3 0.0016726999999999998 3.3 0.0016728 0 0.00167272 0 0.00167282 3.3 0.0016727399999999998 3.3 0.0016728399999999999 0 0.00167276 0 0.00167286 3.3 0.00167278 3.3 0.00167288 0 0.0016728 0 0.0016729 3.3 0.00167282 3.3 0.00167292 0 0.0016728399999999999 0 0.00167294 3.3 0.00167286 3.3 0.00167296 0 0.0016728799999999999 0 0.00167298 3.3 0.0016729 3.3 0.001673 0 0.0016729199999999998 0 0.0016730199999999999 3.3 0.00167294 3.3 0.00167304 0 0.0016729599999999998 0 0.0016730599999999999 3.3 0.00167298 3.3 0.00167308 0 0.001673 0 0.0016731 3.3 0.0016730199999999999 3.3 0.00167312 0 0.00167304 0 0.00167314 3.3 0.0016730599999999999 3.3 0.00167316 0 0.00167308 0 0.00167318 3.3 0.0016730999999999998 3.3 0.0016732 0 0.00167312 0 0.00167322 3.3 0.0016731399999999998 3.3 0.0016732399999999999 0 0.00167316 0 0.00167326 3.3 0.0016731799999999998 3.3 0.0016732799999999999 0 0.0016732 0 0.0016733 3.3 0.00167322 3.3 0.00167332 0 0.0016732399999999999 0 0.00167334 3.3 0.00167326 3.3 0.00167336 0 0.0016732799999999999 0 0.00167338 3.3 0.0016733 3.3 0.0016734 0 0.0016733199999999998 0 0.00167342 3.3 0.00167334 3.3 0.00167344 0 0.0016733599999999998 0 0.0016734599999999999 3.3 0.00167338 3.3 0.00167348 0 0.0016734 0 0.0016735 3.3 0.00167342 3.3 0.00167352 0 0.00167344 0 0.00167354 3.3 0.0016734599999999999 3.3 0.00167356 0 0.00167348 0 0.00167358 3.3 0.0016734999999999999 3.3 0.0016736 0 0.00167352 0 0.00167362 3.3 0.0016735399999999998 3.3 0.00167364 0 0.00167356 0 0.00167366 3.3 0.0016735799999999998 3.3 0.0016736799999999999 0 0.0016736 0 0.0016737 3.3 0.00167362 3.3 0.00167372 0 0.00167364 0 0.00167374 3.3 0.00167366 3.3 0.00167376 0 0.0016736799999999999 0 0.00167378 3.3 0.0016737 3.3 0.0016738 0 0.0016737199999999999 0 0.00167382 3.3 0.00167374 3.3 0.00167384 0 0.0016737599999999998 0 0.0016738599999999999 3.3 0.00167378 3.3 0.00167388 0 0.0016737999999999998 0 0.0016738999999999999 3.3 0.00167382 3.3 0.00167392 0 0.00167384 0 0.00167394 3.3 0.0016738599999999999 3.3 0.00167396 0 0.00167388 0 0.00167398 3.3 0.0016738999999999999 3.3 0.001674 0 0.00167392 0 0.00167402 3.3 0.0016739399999999998 3.3 0.00167404 0 0.00167396 0 0.00167406 3.3 0.0016739799999999998 3.3 0.0016740799999999999 0 0.001674 0 0.0016741 3.3 0.0016740199999999998 3.3 0.0016741199999999999 0 0.00167404 0 0.00167414 3.3 0.00167406 3.3 0.00167416 0 0.0016740799999999999 0 0.00167418 3.3 0.0016741 3.3 0.0016742 0 0.0016741199999999999 0 0.00167422 3.3 0.00167414 3.3 0.00167424 0 0.0016741599999999998 0 0.00167426 3.3 0.00167418 3.3 0.00167428 0 0.0016741999999999998 0 0.0016742999999999999 3.3 0.00167422 3.3 0.00167432 0 0.00167424 0 0.00167434 3.3 0.00167426 3.3 0.00167436 0 0.00167428 0 0.00167438 3.3 0.0016742999999999999 3.3 0.0016744 0 0.00167432 0 0.00167442 3.3 0.0016743399999999999 3.3 0.00167444 0 0.00167436 0 0.00167446 3.3 0.0016743799999999998 3.3 0.00167448 0 0.0016744 0 0.0016745 3.3 0.0016744199999999998 3.3 0.0016745199999999999 0 0.00167444 0 0.00167454 3.3 0.00167446 3.3 0.00167456 0 0.00167448 0 0.00167458 3.3 0.0016745 3.3 0.0016746 0 0.0016745199999999999 0 0.00167462 3.3 0.00167454 3.3 0.00167464 0 0.0016745599999999999 0 0.00167466 3.3 0.00167458 3.3 0.00167468 0 0.0016745999999999998 0 0.0016746999999999999 3.3 0.00167462 3.3 0.00167472 0 0.0016746399999999998 0 0.0016747399999999999 3.3 0.00167466 3.3 0.00167476 0 0.00167468 0 0.00167478 3.3 0.0016746999999999999 3.3 0.0016748 0 0.00167472 0 0.00167482 3.3 0.0016747399999999999 3.3 0.00167484 0 0.00167476 0 0.00167486 3.3 0.0016747799999999998 3.3 0.00167488 0 0.0016748 0 0.0016749 3.3 0.0016748199999999998 3.3 0.0016749199999999999 0 0.00167484 0 0.00167494 3.3 0.0016748599999999998 3.3 0.0016749599999999999 0 0.00167488 0 0.00167498 3.3 0.0016749 3.3 0.001675 0 0.0016749199999999999 0 0.00167502 3.3 0.00167494 3.3 0.00167504 0 0.0016749599999999999 0 0.00167506 3.3 0.00167498 3.3 0.00167508 0 0.0016749999999999998 0 0.0016751 3.3 0.00167502 3.3 0.00167512 0 0.0016750399999999998 0 0.0016751399999999999 3.3 0.00167506 3.3 0.00167516 0 0.00167508 0 0.00167518 3.3 0.0016751 3.3 0.0016752 0 0.00167512 0 0.00167522 3.3 0.0016751399999999999 3.3 0.00167524 0 0.00167516 0 0.00167526 3.3 0.0016751799999999999 3.3 0.00167528 0 0.0016752 0 0.0016753 3.3 0.0016752199999999998 3.3 0.0016753199999999999 0 0.00167524 0 0.00167534 3.3 0.0016752599999999998 3.3 0.0016753599999999999 0 0.00167528 0 0.00167538 3.3 0.0016753 3.3 0.0016754 0 0.0016753199999999999 0 0.00167542 3.3 0.00167534 3.3 0.00167544 0 0.0016753599999999999 0 0.00167546 3.3 0.00167538 3.3 0.00167548 0 0.0016753999999999998 0 0.0016755 3.3 0.00167542 3.3 0.00167552 0 0.0016754399999999998 0 0.0016755399999999999 3.3 0.00167546 3.3 0.00167556 0 0.0016754799999999998 0 0.0016755799999999999 3.3 0.0016755 3.3 0.0016756 0 0.00167552 0 0.00167562 3.3 0.0016755399999999999 3.3 0.00167564 0 0.00167556 0 0.00167566 3.3 0.0016755799999999999 3.3 0.00167568 0 0.0016756 0 0.0016757 3.3 0.0016756199999999998 3.3 0.00167572 0 0.00167564 0 0.00167574 3.3 0.0016756599999999998 3.3 0.0016757599999999999 0 0.00167568 0 0.00167578 3.3 0.0016756999999999998 3.3 0.0016757999999999999 0 0.00167572 0 0.00167582 3.3 0.00167574 3.3 0.00167584 0 0.0016757599999999999 0 0.00167586 3.3 0.00167578 3.3 0.00167588 0 0.0016757999999999999 0 0.0016759 3.3 0.00167582 3.3 0.00167592 0 0.0016758399999999998 0 0.00167594 3.3 0.00167586 3.3 0.00167596 0 0.0016758799999999998 0 0.0016759799999999999 3.3 0.0016759 3.3 0.001676 0 0.00167592 0 0.00167602 3.3 0.00167594 3.3 0.00167604 0 0.00167596 0 0.00167606 3.3 0.0016759799999999999 3.3 0.00167608 0 0.001676 0 0.0016761 3.3 0.0016760199999999999 3.3 0.00167612 0 0.00167604 0 0.00167614 3.3 0.0016760599999999998 3.3 0.0016761599999999999 0 0.00167608 0 0.00167618 3.3 0.0016760999999999998 3.3 0.0016761999999999999 0 0.00167612 0 0.00167622 3.3 0.00167614 3.3 0.00167624 0 0.0016761599999999999 0 0.00167626 3.3 0.00167618 3.3 0.00167628 0 0.0016761999999999999 0 0.0016763 3.3 0.00167622 3.3 0.00167632 0 0.0016762399999999998 0 0.00167634 3.3 0.00167626 3.3 0.00167636 0 0.0016762799999999998 0 0.0016763799999999999 3.3 0.0016763 3.3 0.0016764 0 0.0016763199999999998 0 0.0016764199999999999 3.3 0.00167634 3.3 0.00167644 0 0.00167636 0 0.00167646 3.3 0.0016763799999999999 3.3 0.00167648 0 0.0016764 0 0.0016765 3.3 0.0016764199999999999 3.3 0.00167652 0 0.00167644 0 0.00167654 3.3 0.0016764599999999998 3.3 0.00167656 0 0.00167648 0 0.00167658 3.3 0.0016764999999999998 3.3 0.0016765999999999999 0 0.00167652 0 0.00167662 3.3 0.0016765399999999998 3.3 0.0016766399999999999 0 0.00167656 0 0.00167666 3.3 0.00167658 3.3 0.00167668 0 0.0016765999999999999 0 0.0016767 3.3 0.00167662 3.3 0.00167672 0 0.0016766399999999999 0 0.00167674 3.3 0.00167666 3.3 0.00167676 0 0.0016766799999999998 0 0.00167678 3.3 0.0016767 3.3 0.0016768 0 0.0016767199999999998 0 0.0016768199999999999 3.3 0.00167674 3.3 0.00167684 0 0.00167676 0 0.00167686 3.3 0.00167678 3.3 0.00167688 0 0.0016768 0 0.0016769 3.3 0.0016768199999999999 3.3 0.00167692 0 0.00167684 0 0.00167694 3.3 0.0016768599999999999 3.3 0.00167696 0 0.00167688 0 0.00167698 3.3 0.0016768999999999998 3.3 0.0016769999999999999 0 0.00167692 0 0.00167702 3.3 0.0016769399999999998 3.3 0.0016770399999999999 0 0.00167696 0 0.00167706 3.3 0.00167698 3.3 0.00167708 0 0.0016769999999999999 0 0.0016771 3.3 0.00167702 3.3 0.00167712 0 0.0016770399999999999 0 0.00167714 3.3 0.00167706 3.3 0.00167716 0 0.0016770799999999998 0 0.00167718 3.3 0.0016771 3.3 0.0016772 0 0.0016771199999999998 0 0.0016772199999999999 3.3 0.00167714 3.3 0.00167724 0 0.0016771599999999998 0 0.0016772599999999999 3.3 0.00167718 3.3 0.00167728 0 0.0016772 0 0.0016773 3.3 0.0016772199999999999 3.3 0.00167732 0 0.00167724 0 0.00167734 3.3 0.0016772599999999999 3.3 0.00167736 0 0.00167728 0 0.00167738 3.3 0.0016772999999999998 3.3 0.0016774 0 0.00167732 0 0.00167742 3.3 0.0016773399999999998 3.3 0.0016774399999999999 0 0.00167736 0 0.00167746 3.3 0.00167738 3.3 0.00167748 0 0.0016774 0 0.0016775 3.3 0.00167742 3.3 0.00167752 0 0.0016774399999999999 0 0.00167754 3.3 0.00167746 3.3 0.00167756 0 0.0016774799999999999 0 0.00167758 3.3 0.0016775 3.3 0.0016776 0 0.0016775199999999998 0 0.00167762 3.3 0.00167754 3.3 0.00167764 0 0.0016775599999999998 0 0.0016776599999999999 3.3 0.00167758 3.3 0.00167768 0 0.0016776 0 0.0016777 3.3 0.00167762 3.3 0.00167772 0 0.00167764 0 0.00167774 3.3 0.0016776599999999999 3.3 0.00167776 0 0.00167768 0 0.00167778 3.3 0.0016776999999999999 3.3 0.0016778 0 0.00167772 0 0.00167782 3.3 0.0016777399999999998 3.3 0.0016778399999999999 0 0.00167776 0 0.00167786 3.3 0.0016777799999999998 3.3 0.0016778799999999999 0 0.0016778 0 0.0016779 3.3 0.00167782 3.3 0.00167792 0 0.0016778399999999999 0 0.00167794 3.3 0.00167786 3.3 0.00167796 0 0.0016778799999999999 0 0.00167798 3.3 0.0016779 3.3 0.001678 0 0.0016779199999999998 0 0.00167802 3.3 0.00167794 3.3 0.00167804 0 0.0016779599999999998 0 0.0016780599999999999 3.3 0.00167798 3.3 0.00167808 0 0.0016779999999999998 0 0.0016780999999999999 3.3 0.00167802 3.3 0.00167812 0 0.00167804 0 0.00167814 3.3 0.0016780599999999999 3.3 0.00167816 0 0.00167808 0 0.00167818 3.3 0.0016780999999999999 3.3 0.0016782 0 0.00167812 0 0.00167822 3.3 0.0016781399999999998 3.3 0.00167824 0 0.00167816 0 0.00167826 3.3 0.0016781799999999998 3.3 0.0016782799999999999 0 0.0016782 0 0.0016783 3.3 0.00167822 3.3 0.00167832 0 0.00167824 0 0.00167834 3.3 0.00167826 3.3 0.00167836 0 0.0016782799999999999 0 0.00167838 3.3 0.0016783 3.3 0.0016784 0 0.0016783199999999999 0 0.00167842 3.3 0.00167834 3.3 0.00167844 0 0.0016783599999999998 0 0.0016784599999999999 3.3 0.00167838 3.3 0.00167848 0 0.0016783999999999998 0 0.0016784999999999999 3.3 0.00167842 3.3 0.00167852 0 0.00167844 0 0.00167854 3.3 0.0016784599999999999 3.3 0.00167856 0 0.00167848 0 0.00167858 3.3 0.0016784999999999999 3.3 0.0016786 0 0.00167852 0 0.00167862 3.3 0.0016785399999999998 3.3 0.00167864 0 0.00167856 0 0.00167866 3.3 0.0016785799999999998 3.3 0.0016786799999999999 0 0.0016786 0 0.0016787 3.3 0.0016786199999999998 3.3 0.0016787199999999999 0 0.00167864 0 0.00167874 3.3 0.00167866 3.3 0.00167876 0 0.0016786799999999999 0 0.00167878 3.3 0.0016787 3.3 0.0016788 0 0.0016787199999999999 0 0.00167882 3.3 0.00167874 3.3 0.00167884 0 0.0016787599999999998 0 0.00167886 3.3 0.00167878 3.3 0.00167888 0 0.0016787999999999998 0 0.0016788999999999999 3.3 0.00167882 3.3 0.00167892 0 0.0016788399999999998 0 0.0016789399999999999 3.3 0.00167886 3.3 0.00167896 0 0.00167888 0 0.00167898 3.3 0.0016788999999999999 3.3 0.001679 0 0.00167892 0 0.00167902 3.3 0.0016789399999999999 3.3 0.00167904 0 0.00167896 0 0.00167906 3.3 0.0016789799999999998 3.3 0.00167908 0 0.001679 0 0.0016791 3.3 0.0016790199999999998 3.3 0.0016791199999999999 0 0.00167904 0 0.00167914 3.3 0.00167906 3.3 0.00167916 0 0.00167908 0 0.00167918 3.3 0.0016791 3.3 0.0016792 0 0.0016791199999999999 0 0.00167922 3.3 0.00167914 3.3 0.00167924 0 0.0016791599999999999 0 0.00167926 3.3 0.00167918 3.3 0.00167928 0 0.0016791999999999998 0 0.0016792999999999999 3.3 0.00167922 3.3 0.00167932 0 0.0016792399999999998 0 0.0016793399999999999 3.3 0.00167926 3.3 0.00167936 0 0.00167928 0 0.00167938 3.3 0.0016792999999999999 3.3 0.0016794 0 0.00167932 0 0.00167942 3.3 0.0016793399999999999 3.3 0.00167944 0 0.00167936 0 0.00167946 3.3 0.0016793799999999998 3.3 0.00167948 0 0.0016794 0 0.0016795 3.3 0.0016794199999999998 3.3 0.0016795199999999999 0 0.00167944 0 0.00167954 3.3 0.0016794599999999998 3.3 0.0016795599999999999 0 0.00167948 0 0.00167958 3.3 0.0016795 3.3 0.0016796 0 0.0016795199999999999 0 0.00167962 3.3 0.00167954 3.3 0.00167964 0 0.0016795599999999999 0 0.00167966 3.3 0.00167958 3.3 0.00167968 0 0.0016795999999999998 0 0.0016797 3.3 0.00167962 3.3 0.00167972 0 0.0016796399999999998 0 0.0016797399999999999 3.3 0.00167966 3.3 0.00167976 0 0.0016796799999999998 0 0.0016797799999999999 3.3 0.0016797 3.3 0.0016798 0 0.00167972 0 0.00167982 3.3 0.0016797399999999999 3.3 0.00167984 0 0.00167976 0 0.00167986 3.3 0.0016797799999999999 3.3 0.00167988 0 0.0016798 0 0.0016799 3.3 0.0016798199999999998 3.3 0.00167992 0 0.00167984 0 0.00167994 3.3 0.0016798599999999998 3.3 0.0016799599999999999 0 0.00167988 0 0.00167998 3.3 0.0016799 3.3 0.00168 0 0.00167992 0 0.00168002 3.3 0.00167994 3.3 0.00168004 0 0.0016799599999999999 0 0.00168006 3.3 0.00167998 3.3 0.00168008 0 0.0016799999999999999 0 0.0016801 3.3 0.00168002 3.3 0.00168012 0 0.0016800399999999998 0 0.0016801399999999999 3.3 0.00168006 3.3 0.00168016 0 0.0016800799999999998 0 0.0016801799999999999 3.3 0.0016801 3.3 0.0016802 0 0.00168012 0 0.00168022 3.3 0.0016801399999999999 3.3 0.00168024 0 0.00168016 0 0.00168026 3.3 0.0016801799999999999 3.3 0.00168028 0 0.0016802 0 0.0016803 3.3 0.0016802199999999998 3.3 0.00168032 0 0.00168024 0 0.00168034 3.3 0.0016802599999999998 3.3 0.0016803599999999999 0 0.00168028 0 0.00168038 3.3 0.0016802999999999998 3.3 0.0016803999999999999 0 0.00168032 0 0.00168042 3.3 0.00168034 3.3 0.00168044 0 0.0016803599999999999 0 0.00168046 3.3 0.00168038 3.3 0.00168048 0 0.0016803999999999999 0 0.0016805 3.3 0.00168042 3.3 0.00168052 0 0.0016804399999999998 0 0.00168054 3.3 0.00168046 3.3 0.00168056 0 0.0016804799999999998 0 0.0016805799999999999 3.3 0.0016805 3.3 0.0016806 0 0.00168052 0 0.00168062 3.3 0.00168054 3.3 0.00168064 0 0.00168056 0 0.00168066 3.3 0.0016805799999999999 3.3 0.00168068 0 0.0016806 0 0.0016807 3.3 0.0016806199999999999 3.3 0.00168072 0 0.00168064 0 0.00168074 3.3 0.0016806599999999998 3.3 0.00168076 0 0.00168068 0 0.00168078 3.3 0.0016806999999999998 3.3 0.0016807999999999999 0 0.00168072 0 0.00168082 3.3 0.00168074 3.3 0.00168084 0 0.00168076 0 0.00168086 3.3 0.00168078 3.3 0.00168088 0 0.0016807999999999999 0 0.0016809 3.3 0.00168082 3.3 0.00168092 0 0.0016808399999999999 0 0.00168094 3.3 0.00168086 3.3 0.00168096 0 0.0016808799999999998 0 0.0016809799999999999 3.3 0.0016809 3.3 0.001681 0 0.0016809199999999998 0 0.0016810199999999999 3.3 0.00168094 3.3 0.00168104 0 0.00168096 0 0.00168106 3.3 0.0016809799999999999 3.3 0.00168108 0 0.001681 0 0.0016811 3.3 0.0016810199999999999 3.3 0.00168112 0 0.00168104 0 0.00168114 3.3 0.0016810599999999998 3.3 0.00168116 0 0.00168108 0 0.00168118 3.3 0.0016810999999999998 3.3 0.0016811999999999999 0 0.00168112 0 0.00168122 3.3 0.0016811399999999998 3.3 0.0016812399999999999 0 0.00168116 0 0.00168126 3.3 0.00168118 3.3 0.00168128 0 0.0016811999999999999 0 0.0016813 3.3 0.00168122 3.3 0.00168132 0 0.0016812399999999999 0 0.00168134 3.3 0.00168126 3.3 0.00168136 0 0.0016812799999999998 0 0.00168138 3.3 0.0016813 3.3 0.0016814 0 0.0016813199999999998 0 0.0016814199999999999 3.3 0.00168134 3.3 0.00168144 0 0.00168136 0 0.00168146 3.3 0.00168138 3.3 0.00168148 0 0.0016814 0 0.0016815 3.3 0.0016814199999999999 3.3 0.00168152 0 0.00168144 0 0.00168154 3.3 0.0016814599999999999 3.3 0.00168156 0 0.00168148 0 0.00168158 3.3 0.0016814999999999998 3.3 0.0016816 0 0.00168152 0 0.00168162 3.3 0.0016815399999999998 3.3 0.0016816399999999999 0 0.00168156 0 0.00168166 3.3 0.00168158 3.3 0.00168168 0 0.0016816 0 0.0016817 3.3 0.00168162 3.3 0.00168172 0 0.0016816399999999999 0 0.00168174 3.3 0.00168166 3.3 0.00168176 0 0.0016816799999999999 0 0.00168178 3.3 0.0016817 3.3 0.0016818 0 0.0016817199999999998 0 0.0016818199999999999 3.3 0.00168174 3.3 0.00168184 0 0.0016817599999999998 0 0.0016818599999999999 3.3 0.00168178 3.3 0.00168188 0 0.0016818 0 0.0016819 3.3 0.0016818199999999999 3.3 0.00168192 0 0.00168184 0 0.00168194 3.3 0.0016818599999999999 3.3 0.00168196 0 0.00168188 0 0.00168198 3.3 0.0016818999999999998 3.3 0.001682 0 0.00168192 0 0.00168202 3.3 0.0016819399999999998 3.3 0.0016820399999999999 0 0.00168196 0 0.00168206 3.3 0.0016819799999999998 3.3 0.0016820799999999999 0 0.001682 0 0.0016821 3.3 0.00168202 3.3 0.00168212 0 0.0016820399999999999 0 0.00168214 3.3 0.00168206 3.3 0.00168216 0 0.0016820799999999999 0 0.00168218 3.3 0.0016821 3.3 0.0016822 0 0.0016821199999999998 0 0.00168222 3.3 0.00168214 3.3 0.00168224 0 0.0016821599999999998 0 0.0016822599999999999 3.3 0.00168218 3.3 0.00168228 0 0.0016822 0 0.0016823 3.3 0.00168222 3.3 0.00168232 0 0.00168224 0 0.00168234 3.3 0.0016822599999999999 3.3 0.00168236 0 0.00168228 0 0.00168238 3.3 0.0016822999999999999 3.3 0.0016824 0 0.00168232 0 0.00168242 3.3 0.0016823399999999998 3.3 0.0016824399999999999 0 0.00168236 0 0.00168246 3.3 0.0016823799999999998 3.3 0.0016824799999999999 0 0.0016824 0 0.0016825 3.3 0.00168242 3.3 0.00168252 0 0.0016824399999999999 0 0.00168254 3.3 0.00168246 3.3 0.00168256 0 0.0016824799999999999 0 0.00168258 3.3 0.0016825 3.3 0.0016826 0 0.0016825199999999998 0 0.00168262 3.3 0.00168254 3.3 0.00168264 0 0.0016825599999999998 0 0.0016826599999999999 3.3 0.00168258 3.3 0.00168268 0 0.0016825999999999998 0 0.0016826999999999999 3.3 0.00168262 3.3 0.00168272 0 0.00168264 0 0.00168274 3.3 0.0016826599999999999 3.3 0.00168276 0 0.00168268 0 0.00168278 3.3 0.0016826999999999999 3.3 0.0016828 0 0.00168272 0 0.00168282 3.3 0.0016827399999999998 3.3 0.00168284 0 0.00168276 0 0.00168286 3.3 0.0016827799999999998 3.3 0.0016828799999999999 0 0.0016828 0 0.0016829 3.3 0.0016828199999999998 3.3 0.0016829199999999999 0 0.00168284 0 0.00168294 3.3 0.00168286 3.3 0.00168296 0 0.0016828799999999999 0 0.00168298 3.3 0.0016829 3.3 0.001683 0 0.0016829199999999999 0 0.00168302 3.3 0.00168294 3.3 0.00168304 0 0.0016829599999999998 0 0.00168306 3.3 0.00168298 3.3 0.00168308 0 0.0016829999999999998 0 0.0016830999999999999 3.3 0.00168302 3.3 0.00168312 0 0.00168304 0 0.00168314 3.3 0.00168306 3.3 0.00168316 0 0.00168308 0 0.00168318 3.3 0.0016830999999999999 3.3 0.0016832 0 0.00168312 0 0.00168322 3.3 0.0016831399999999999 3.3 0.00168324 0 0.00168316 0 0.00168326 3.3 0.0016831799999999998 3.3 0.0016832799999999999 0 0.0016832 0 0.0016833 3.3 0.0016832199999999998 3.3 0.0016833199999999999 0 0.00168324 0 0.00168334 3.3 0.00168326 3.3 0.00168336 0 0.0016832799999999999 0 0.00168338 3.3 0.0016833 3.3 0.0016834 0 0.0016833199999999999 0 0.00168342 3.3 0.00168334 3.3 0.00168344 0 0.0016833599999999998 0 0.00168346 3.3 0.00168338 3.3 0.00168348 0 0.0016833999999999998 0 0.0016834999999999999 3.3 0.00168342 3.3 0.00168352 0 0.0016834399999999998 0 0.0016835399999999999 3.3 0.00168346 3.3 0.00168356 0 0.00168348 0 0.00168358 3.3 0.0016834999999999999 3.3 0.0016836 0 0.00168352 0 0.00168362 3.3 0.0016835399999999999 3.3 0.00168364 0 0.00168356 0 0.00168366 3.3 0.0016835799999999998 3.3 0.00168368 0 0.0016836 0 0.0016837 3.3 0.0016836199999999998 3.3 0.0016837199999999999 0 0.00168364 0 0.00168374 3.3 0.00168366 3.3 0.00168376 0 0.00168368 0 0.00168378 3.3 0.0016837 3.3 0.0016838 0 0.0016837199999999999 0 0.00168382 3.3 0.00168374 3.3 0.00168384 0 0.0016837599999999999 0 0.00168386 3.3 0.00168378 3.3 0.00168388 0 0.0016837999999999998 0 0.0016839 3.3 0.00168382 3.3 0.00168392 0 0.0016838399999999998 0 0.0016839399999999999 3.3 0.00168386 3.3 0.00168396 0 0.00168388 0 0.00168398 3.3 0.0016839 3.3 0.001684 0 0.00168392 0 0.00168402 3.3 0.0016839399999999999 3.3 0.00168404 0 0.00168396 0 0.00168406 3.3 0.0016839799999999999 3.3 0.00168408 0 0.001684 0 0.0016841 3.3 0.0016840199999999998 3.3 0.0016841199999999999 0 0.00168404 0 0.00168414 3.3 0.0016840599999999998 3.3 0.0016841599999999999 0 0.00168408 0 0.00168418 3.3 0.0016841 3.3 0.0016842 0 0.0016841199999999999 0 0.00168422 3.3 0.00168414 3.3 0.00168424 0 0.0016841599999999999 0 0.00168426 3.3 0.00168418 3.3 0.00168428 0 0.0016841999999999998 0 0.0016843 3.3 0.00168422 3.3 0.00168432 0 0.0016842399999999998 0 0.0016843399999999999 3.3 0.00168426 3.3 0.00168436 0 0.0016842799999999998 0 0.0016843799999999999 3.3 0.0016843 3.3 0.0016844 0 0.00168432 0 0.00168442 3.3 0.0016843399999999999 3.3 0.00168444 0 0.00168436 0 0.00168446 3.3 0.0016843799999999999 3.3 0.00168448 0 0.0016844 0 0.0016845 3.3 0.0016844199999999998 3.3 0.00168452 0 0.00168444 0 0.00168454 3.3 0.0016844599999999998 3.3 0.0016845599999999999 0 0.00168448 0 0.00168458 3.3 0.0016845 3.3 0.0016846 0 0.00168452 0 0.00168462 3.3 0.00168454 3.3 0.00168464 0 0.0016845599999999999 0 0.00168466 3.3 0.00168458 3.3 0.00168468 0 0.0016845999999999999 0 0.0016847 3.3 0.00168462 3.3 0.00168472 0 0.0016846399999999998 0 0.00168474 3.3 0.00168466 3.3 0.00168476 0 0.0016846799999999998 0 0.0016847799999999999 3.3 0.0016847 3.3 0.0016848 0 0.00168472 0 0.00168482 3.3 0.00168474 3.3 0.00168484 0 0.00168476 0 0.00168486 3.3 0.0016847799999999999 3.3 0.00168488 0 0.0016848 0 0.0016849 3.3 0.0016848199999999999 3.3 0.00168492 0 0.00168484 0 0.00168494 3.3 0.0016848599999999998 3.3 0.0016849599999999999 0 0.00168488 0 0.00168498 3.3 0.0016848999999999998 3.3 0.0016849999999999999 0 0.00168492 0 0.00168502 3.3 0.00168494 3.3 0.00168504 0 0.0016849599999999999 0 0.00168506 3.3 0.00168498 3.3 0.00168508 0 0.0016849999999999999 0 0.0016851 3.3 0.00168502 3.3 0.00168512 0 0.0016850399999999998 0 0.00168514 3.3 0.00168506 3.3 0.00168516 0 0.0016850799999999998 0 0.0016851799999999999 3.3 0.0016851 3.3 0.0016852 0 0.0016851199999999998 0 0.0016852199999999999 3.3 0.00168514 3.3 0.00168524 0 0.00168516 0 0.00168526 3.3 0.0016851799999999999 3.3 0.00168528 0 0.0016852 0 0.0016853 3.3 0.0016852199999999999 3.3 0.00168532 0 0.00168524 0 0.00168534 3.3 0.0016852599999999998 3.3 0.00168536 0 0.00168528 0 0.00168538 3.3 0.0016852999999999998 3.3 0.0016853999999999999 0 0.00168532 0 0.00168542 3.3 0.00168534 3.3 0.00168544 0 0.00168536 0 0.00168546 3.3 0.00168538 3.3 0.00168548 0 0.0016853999999999999 0 0.0016855 3.3 0.00168542 3.3 0.00168552 0 0.0016854399999999999 0 0.00168554 3.3 0.00168546 3.3 0.00168556 0 0.0016854799999999998 0 0.0016855799999999999 3.3 0.0016855 3.3 0.0016856 0 0.0016855199999999998 0 0.0016856199999999999 3.3 0.00168554 3.3 0.00168564 0 0.00168556 0 0.00168566 3.3 0.0016855799999999999 3.3 0.00168568 0 0.0016856 0 0.0016857 3.3 0.0016856199999999999 3.3 0.00168572 0 0.00168564 0 0.00168574 3.3 0.0016856599999999998 3.3 0.00168576 0 0.00168568 0 0.00168578 3.3 0.0016856999999999998 3.3 0.0016857999999999999 0 0.00168572 0 0.00168582 3.3 0.0016857399999999998 3.3 0.0016858399999999999 0 0.00168576 0 0.00168586 3.3 0.00168578 3.3 0.00168588 0 0.0016857999999999999 0 0.0016859 3.3 0.00168582 3.3 0.00168592 0 0.0016858399999999999 0 0.00168594 3.3 0.00168586 3.3 0.00168596 0 0.0016858799999999998 0 0.00168598 3.3 0.0016859 3.3 0.001686 0 0.0016859199999999998 0 0.0016860199999999999 3.3 0.00168594 3.3 0.00168604 0 0.0016859599999999998 0 0.0016860599999999999 3.3 0.00168598 3.3 0.00168608 0 0.001686 0 0.0016861 3.3 0.0016860199999999999 3.3 0.00168612 0 0.00168604 0 0.00168614 3.3 0.0016860599999999999 3.3 0.00168616 0 0.00168608 0 0.00168618 3.3 0.0016860999999999998 3.3 0.0016862 0 0.00168612 0 0.00168622 3.3 0.0016861399999999998 3.3 0.0016862399999999999 0 0.00168616 0 0.00168626 3.3 0.00168618 3.3 0.00168628 0 0.0016862 0 0.0016863 3.3 0.00168622 3.3 0.00168632 0 0.0016862399999999999 0 0.00168634 3.3 0.00168626 3.3 0.00168636 0 0.0016862799999999999 0 0.00168638 3.3 0.0016863 3.3 0.0016864 0 0.0016863199999999998 0 0.0016864199999999999 3.3 0.00168634 3.3 0.00168644 0 0.0016863599999999998 0 0.0016864599999999999 3.3 0.00168638 3.3 0.00168648 0 0.0016864 0 0.0016865 3.3 0.0016864199999999999 3.3 0.00168652 0 0.00168644 0 0.00168654 3.3 0.0016864599999999999 3.3 0.00168656 0 0.00168648 0 0.00168658 3.3 0.0016864999999999998 3.3 0.0016866 0 0.00168652 0 0.00168662 3.3 0.0016865399999999998 3.3 0.0016866399999999999 0 0.00168656 0 0.00168666 3.3 0.0016865799999999998 3.3 0.0016866799999999999 0 0.0016866 0 0.0016867 3.3 0.00168662 3.3 0.00168672 0 0.0016866399999999999 0 0.00168674 3.3 0.00168666 3.3 0.00168676 0 0.0016866799999999999 0 0.00168678 3.3 0.0016867 3.3 0.0016868 0 0.0016867199999999998 0 0.00168682 3.3 0.00168674 3.3 0.00168684 0 0.0016867599999999998 0 0.0016868599999999999 3.3 0.00168678 3.3 0.00168688 0 0.0016867999999999998 0 0.0016868999999999999 3.3 0.00168682 3.3 0.00168692 0 0.00168684 0 0.00168694 3.3 0.0016868599999999999 3.3 0.00168696 0 0.00168688 0 0.00168698 3.3 0.0016868999999999999 3.3 0.001687 0 0.00168692 0 0.00168702 3.3 0.0016869399999999998 3.3 0.00168704 0 0.00168696 0 0.00168706 3.3 0.0016869799999999998 3.3 0.0016870799999999999 0 0.001687 0 0.0016871 3.3 0.00168702 3.3 0.00168712 0 0.00168704 0 0.00168714 3.3 0.00168706 3.3 0.00168716 0 0.0016870799999999999 0 0.00168718 3.3 0.0016871 3.3 0.0016872 0 0.0016871199999999999 0 0.00168722 3.3 0.00168714 3.3 0.00168724 0 0.0016871599999999998 0 0.0016872599999999999 3.3 0.00168718 3.3 0.00168728 0 0.0016871999999999998 0 0.0016872999999999999 3.3 0.00168722 3.3 0.00168732 0 0.00168724 0 0.00168734 3.3 0.0016872599999999999 3.3 0.00168736 0 0.00168728 0 0.00168738 3.3 0.0016872999999999999 3.3 0.0016874 0 0.00168732 0 0.00168742 3.3 0.0016873399999999998 3.3 0.00168744 0 0.00168736 0 0.00168746 3.3 0.0016873799999999998 3.3 0.0016874799999999999 0 0.0016874 0 0.0016875 3.3 0.0016874199999999998 3.3 0.0016875199999999999 0 0.00168744 0 0.00168754 3.3 0.00168746 3.3 0.00168756 0 0.0016874799999999999 0 0.00168758 3.3 0.0016875 3.3 0.0016876 0 0.0016875199999999999 0 0.00168762 3.3 0.00168754 3.3 0.00168764 0 0.0016875599999999998 0 0.00168766 3.3 0.00168758 3.3 0.00168768 0 0.0016875999999999998 0 0.0016876999999999999 3.3 0.00168762 3.3 0.00168772 0 0.00168764 0 0.00168774 3.3 0.00168766 3.3 0.00168776 0 0.00168768 0 0.00168778 3.3 0.0016876999999999999 3.3 0.0016878 0 0.00168772 0 0.00168782 3.3 0.0016877399999999999 3.3 0.00168784 0 0.00168776 0 0.00168786 3.3 0.0016877799999999998 3.3 0.00168788 0 0.0016878 0 0.0016879 3.3 0.0016878199999999998 3.3 0.0016879199999999999 0 0.00168784 0 0.00168794 3.3 0.00168786 3.3 0.00168796 0 0.00168788 0 0.00168798 3.3 0.0016879 3.3 0.001688 0 0.0016879199999999999 0 0.00168802 3.3 0.00168794 3.3 0.00168804 0 0.0016879599999999999 0 0.00168806 3.3 0.00168798 3.3 0.00168808 0 0.0016879999999999998 0 0.0016880999999999999 3.3 0.00168802 3.3 0.00168812 0 0.0016880399999999998 0 0.0016881399999999999 3.3 0.00168806 3.3 0.00168816 0 0.00168808 0 0.00168818 3.3 0.0016880999999999999 3.3 0.0016882 0 0.00168812 0 0.00168822 3.3 0.0016881399999999999 3.3 0.00168824 0 0.00168816 0 0.00168826 3.3 0.0016881799999999998 3.3 0.00168828 0 0.0016882 0 0.0016883 3.3 0.0016882199999999998 3.3 0.0016883199999999999 0 0.00168824 0 0.00168834 3.3 0.0016882599999999998 3.3 0.0016883599999999999 0 0.00168828 0 0.00168838 3.3 0.0016883 3.3 0.0016884 0 0.0016883199999999999 0 0.00168842 3.3 0.00168834 3.3 0.00168844 0 0.0016883599999999999 0 0.00168846 3.3 0.00168838 3.3 0.00168848 0 0.0016883999999999998 0 0.0016885 3.3 0.00168842 3.3 0.00168852 0 0.0016884399999999998 0 0.0016885399999999999 3.3 0.00168846 3.3 0.00168856 0 0.00168848 0 0.00168858 3.3 0.0016885 3.3 0.0016886 0 0.00168852 0 0.00168862 3.3 0.0016885399999999999 3.3 0.00168864 0 0.00168856 0 0.00168866 3.3 0.0016885799999999999 3.3 0.00168868 0 0.0016886 0 0.0016887 3.3 0.0016886199999999998 3.3 0.0016887199999999999 0 0.00168864 0 0.00168874 3.3 0.0016886599999999998 3.3 0.0016887599999999999 0 0.00168868 0 0.00168878 3.3 0.0016887 3.3 0.0016888 0 0.0016887199999999999 0 0.00168882 3.3 0.00168874 3.3 0.00168884 0 0.0016887599999999999 0 0.00168886 3.3 0.00168878 3.3 0.00168888 0 0.0016887999999999998 0 0.0016889 3.3 0.00168882 3.3 0.00168892 0 0.0016888399999999998 0 0.0016889399999999999 3.3 0.00168886 3.3 0.00168896 0 0.0016888799999999998 0 0.0016889799999999999 3.3 0.0016889 3.3 0.001689 0 0.00168892 0 0.00168902 3.3 0.0016889399999999999 3.3 0.00168904 0 0.00168896 0 0.00168906 3.3 0.0016889799999999999 3.3 0.00168908 0 0.001689 0 0.0016891 3.3 0.0016890199999999998 3.3 0.00168912 0 0.00168904 0 0.00168914 3.3 0.0016890599999999998 3.3 0.0016891599999999999 0 0.00168908 0 0.00168918 3.3 0.0016890999999999998 3.3 0.0016891999999999999 0 0.00168912 0 0.00168922 3.3 0.00168914 3.3 0.00168924 0 0.0016891599999999999 0 0.00168926 3.3 0.00168918 3.3 0.00168928 0 0.0016891999999999999 0 0.0016893 3.3 0.00168922 3.3 0.00168932 0 0.0016892399999999998 0 0.00168934 3.3 0.00168926 3.3 0.00168936 0 0.0016892799999999998 0 0.0016893799999999999 3.3 0.0016893 3.3 0.0016894 0 0.00168932 0 0.00168942 3.3 0.00168934 3.3 0.00168944 0 0.00168936 0 0.00168946 3.3 0.0016893799999999999 3.3 0.00168948 0 0.0016894 0 0.0016895 3.3 0.0016894199999999999 3.3 0.00168952 0 0.00168944 0 0.00168954 3.3 0.0016894599999999998 3.3 0.0016895599999999999 0 0.00168948 0 0.00168958 3.3 0.0016894999999999998 3.3 0.0016895999999999999 0 0.00168952 0 0.00168962 3.3 0.00168954 3.3 0.00168964 0 0.0016895599999999999 0 0.00168966 3.3 0.00168958 3.3 0.00168968 0 0.0016895999999999999 0 0.0016897 3.3 0.00168962 3.3 0.00168972 0 0.0016896399999999998 0 0.00168974 3.3 0.00168966 3.3 0.00168976 0 0.0016896799999999998 0 0.0016897799999999999 3.3 0.0016897 3.3 0.0016898 0 0.0016897199999999998 0 0.0016898199999999999 3.3 0.00168974 3.3 0.00168984 0 0.00168976 0 0.00168986 3.3 0.0016897799999999999 3.3 0.00168988 0 0.0016898 0 0.0016899 3.3 0.0016898199999999999 3.3 0.00168992 0 0.00168984 0 0.00168994 3.3 0.0016898599999999998 3.3 0.00168996 0 0.00168988 0 0.00168998 3.3 0.0016898999999999998 3.3 0.0016899999999999999 0 0.00168992 0 0.00169002 3.3 0.0016899399999999998 3.3 0.0016900399999999999 0 0.00168996 0 0.00169006 3.3 0.00168998 3.3 0.00169008 0 0.0016899999999999999 0 0.0016901 3.3 0.00169002 3.3 0.00169012 0 0.0016900399999999999 0 0.00169014 3.3 0.00169006 3.3 0.00169016 0 0.0016900799999999998 0 0.00169018 3.3 0.0016901 3.3 0.0016902 0 0.0016901199999999998 0 0.0016902199999999999 3.3 0.00169014 3.3 0.00169024 0 0.00169016 0 0.00169026 3.3 0.00169018 3.3 0.00169028 0 0.0016902 0 0.0016903 3.3 0.0016902199999999999 3.3 0.00169032 0 0.00169024 0 0.00169034 3.3 0.0016902599999999999 3.3 0.00169036 0 0.00169028 0 0.00169038 3.3 0.0016902999999999998 3.3 0.0016903999999999999 0 0.00169032 0 0.00169042 3.3 0.0016903399999999998 3.3 0.0016904399999999999 0 0.00169036 0 0.00169046 3.3 0.00169038 3.3 0.00169048 0 0.0016903999999999999 0 0.0016905 3.3 0.00169042 3.3 0.00169052 0 0.0016904399999999999 0 0.00169054 3.3 0.00169046 3.3 0.00169056 0 0.0016904799999999998 0 0.00169058 3.3 0.0016905 3.3 0.0016906 0 0.0016905199999999998 0 0.0016906199999999999 3.3 0.00169054 3.3 0.00169064 0 0.0016905599999999998 0 0.0016906599999999999 3.3 0.00169058 3.3 0.00169068 0 0.0016906 0 0.0016907 3.3 0.0016906199999999999 3.3 0.00169072 0 0.00169064 0 0.00169074 3.3 0.0016906599999999999 3.3 0.00169076 0 0.00169068 0 0.00169078 3.3 0.0016906999999999998 3.3 0.0016908 0 0.00169072 0 0.00169082 3.3 0.0016907399999999998 3.3 0.0016908399999999999 0 0.00169076 0 0.00169086 3.3 0.00169078 3.3 0.00169088 0 0.0016908 0 0.0016909 3.3 0.00169082 3.3 0.00169092 0 0.0016908399999999999 0 0.00169094 3.3 0.00169086 3.3 0.00169096 0 0.0016908799999999999 0 0.00169098 3.3 0.0016909 3.3 0.001691 0 0.0016909199999999998 0 0.00169102 3.3 0.00169094 3.3 0.00169104 0 0.0016909599999999998 0 0.0016910599999999999 3.3 0.00169098 3.3 0.00169108 0 0.001691 0 0.0016911 3.3 0.00169102 3.3 0.00169112 0 0.00169104 0 0.00169114 3.3 0.0016910599999999999 3.3 0.00169116 0 0.00169108 0 0.00169118 3.3 0.0016910999999999999 3.3 0.0016912 0 0.00169112 0 0.00169122 3.3 0.0016911399999999998 3.3 0.0016912399999999999 0 0.00169116 0 0.00169126 3.3 0.0016911799999999998 3.3 0.0016912799999999999 0 0.0016912 0 0.0016913 3.3 0.00169122 3.3 0.00169132 0 0.0016912399999999999 0 0.00169134 3.3 0.00169126 3.3 0.00169136 0 0.0016912799999999999 0 0.00169138 3.3 0.0016913 3.3 0.0016914 0 0.0016913199999999998 0 0.00169142 3.3 0.00169134 3.3 0.00169144 0 0.0016913599999999998 0 0.0016914599999999999 3.3 0.00169138 3.3 0.00169148 0 0.0016913999999999998 0 0.0016914999999999999 3.3 0.00169142 3.3 0.00169152 0 0.00169144 0 0.00169154 3.3 0.0016914599999999999 3.3 0.00169156 0 0.00169148 0 0.00169158 3.3 0.0016914999999999999 3.3 0.0016916 0 0.00169152 0 0.00169162 3.3 0.0016915399999999998 3.3 0.00169164 0 0.00169156 0 0.00169166 3.3 0.0016915799999999998 3.3 0.0016916799999999999 0 0.0016916 0 0.0016917 3.3 0.00169162 3.3 0.00169172 0 0.00169164 0 0.00169174 3.3 0.00169166 3.3 0.00169176 0 0.0016916799999999999 0 0.00169178 3.3 0.0016917 3.3 0.0016918 0 0.0016917199999999999 0 0.00169182 3.3 0.00169174 3.3 0.00169184 0 0.0016917599999999998 0 0.00169186 3.3 0.00169178 3.3 0.00169188 0 0.0016917999999999998 0 0.0016918999999999999 3.3 0.00169182 3.3 0.00169192 0 0.00169184 0 0.00169194 3.3 0.00169186 3.3 0.00169196 0 0.00169188 0 0.00169198 3.3 0.0016918999999999999 3.3 0.001692 0 0.00169192 0 0.00169202 3.3 0.0016919399999999999 3.3 0.00169204 0 0.00169196 0 0.00169206 3.3 0.0016919799999999998 3.3 0.0016920799999999999 0 0.001692 0 0.0016921 3.3 0.0016920199999999998 3.3 0.0016921199999999999 0 0.00169204 0 0.00169214 3.3 0.00169206 3.3 0.00169216 0 0.0016920799999999999 0 0.00169218 3.3 0.0016921 3.3 0.0016922 0 0.0016921199999999999 0 0.00169222 3.3 0.00169214 3.3 0.00169224 0 0.0016921599999999998 0 0.00169226 3.3 0.00169218 3.3 0.00169228 0 0.0016921999999999998 0 0.0016922999999999999 3.3 0.00169222 3.3 0.00169232 0 0.0016922399999999998 0 0.0016923399999999999 3.3 0.00169226 3.3 0.00169236 0 0.00169228 0 0.00169238 3.3 0.0016922999999999999 3.3 0.0016924 0 0.00169232 0 0.00169242 3.3 0.0016923399999999999 3.3 0.00169244 0 0.00169236 0 0.00169246 3.3 0.0016923799999999998 3.3 0.00169248 0 0.0016924 0 0.0016925 3.3 0.0016924199999999998 3.3 0.0016925199999999999 0 0.00169244 0 0.00169254 3.3 0.00169246 3.3 0.00169256 0 0.00169248 0 0.00169258 3.3 0.0016925 3.3 0.0016926 0 0.0016925199999999999 0 0.00169262 3.3 0.00169254 3.3 0.00169264 0 0.0016925599999999999 0 0.00169266 3.3 0.00169258 3.3 0.00169268 0 0.0016925999999999998 0 0.0016926999999999999 3.3 0.00169262 3.3 0.00169272 0 0.0016926399999999998 0 0.0016927399999999999 3.3 0.00169266 3.3 0.00169276 0 0.00169268 0 0.00169278 3.3 0.0016926999999999999 3.3 0.0016928 0 0.00169272 0 0.00169282 3.3 0.0016927399999999999 3.3 0.00169284 0 0.00169276 0 0.00169286 3.3 0.0016927799999999998 3.3 0.00169288 0 0.0016928 0 0.0016929 3.3 0.0016928199999999998 3.3 0.0016929199999999999 0 0.00169284 0 0.00169294 3.3 0.0016928599999999998 3.3 0.0016929599999999999 0 0.00169288 0 0.00169298 3.3 0.0016929 3.3 0.001693 0 0.0016929199999999999 0 0.00169302 3.3 0.00169294 3.3 0.00169304 0 0.0016929599999999999 0 0.00169306 3.3 0.00169298 3.3 0.00169308 0 0.0016929999999999998 0 0.0016931 3.3 0.00169302 3.3 0.00169312 0 0.0016930399999999998 0 0.0016931399999999999 3.3 0.00169306 3.3 0.00169316 0 0.0016930799999999998 0 0.0016931799999999999 3.3 0.0016931 3.3 0.0016932 0 0.00169312 0 0.00169322 3.3 0.0016931399999999999 3.3 0.00169324 0 0.00169316 0 0.00169326 3.3 0.0016931799999999999 3.3 0.00169328 0 0.0016932 0 0.0016933 3.3 0.0016932199999999998 3.3 0.00169332 0 0.00169324 0 0.00169334 3.3 0.0016932599999999998 3.3 0.0016933599999999999 0 0.00169328 0 0.00169338 3.3 0.0016933 3.3 0.0016934 0 0.00169332 0 0.00169342 3.3 0.00169334 3.3 0.00169344 0 0.0016933599999999999 0 0.00169346 3.3 0.00169338 3.3 0.00169348 0 0.0016933999999999999 0 0.0016935 3.3 0.00169342 3.3 0.00169352 0 0.0016934399999999998 0 0.0016935399999999999 3.3 0.00169346 3.3 0.00169356 0 0.0016934799999999998 0 0.0016935799999999999 3.3 0.0016935 3.3 0.0016936 0 0.00169352 0 0.00169362 3.3 0.0016935399999999999 3.3 0.00169364 0 0.00169356 0 0.00169366 3.3 0.0016935799999999999 3.3 0.00169368 0 0.0016936 0 0.0016937 3.3 0.0016936199999999998 3.3 0.00169372 0 0.00169364 0 0.00169374 3.3 0.0016936599999999998 3.3 0.0016937599999999999 0 0.00169368 0 0.00169378 3.3 0.0016936999999999998 3.3 0.0016937999999999999 0 0.00169372 0 0.00169382 3.3 0.00169374 3.3 0.00169384 0 0.0016937599999999999 0 0.00169386 3.3 0.00169378 3.3 0.00169388 0 0.0016937999999999999 0 0.0016939 3.3 0.00169382 3.3 0.00169392 0 0.0016938399999999998 0 0.00169394 3.3 0.00169386 3.3 0.00169396 0 0.0016938799999999998 0 0.0016939799999999999 3.3 0.0016939 3.3 0.001694 0 0.00169392 0 0.00169402 3.3 0.00169394 3.3 0.00169404 0 0.00169396 0 0.00169406 3.3 0.0016939799999999999 3.3 0.00169408 0 0.001694 0 0.0016941 3.3 0.0016940199999999999 3.3 0.00169412 0 0.00169404 0 0.00169414 3.3 0.0016940599999999998 3.3 0.00169416 0 0.00169408 0 0.00169418 3.3 0.0016940999999999998 3.3 0.0016941999999999999 0 0.00169412 0 0.00169422 3.3 0.00169414 3.3 0.00169424 0 0.00169416 0 0.00169426 3.3 0.00169418 3.3 0.00169428 0 0.0016941999999999999 0 0.0016943 3.3 0.00169422 3.3 0.00169432 0 0.0016942399999999999 0 0.00169434 3.3 0.00169426 3.3 0.00169436 0 0.0016942799999999998 0 0.0016943799999999999 3.3 0.0016943 3.3 0.0016944 0 0.0016943199999999998 0 0.0016944199999999999 3.3 0.00169434 3.3 0.00169444 0 0.00169436 0 0.00169446 3.3 0.0016943799999999999 3.3 0.00169448 0 0.0016944 0 0.0016945 3.3 0.0016944199999999999 3.3 0.00169452 0 0.00169444 0 0.00169454 3.3 0.0016944599999999998 3.3 0.00169456 0 0.00169448 0 0.00169458 3.3 0.0016944999999999998 3.3 0.0016945999999999999 0 0.00169452 0 0.00169462 3.3 0.0016945399999999998 3.3 0.0016946399999999999 0 0.00169456 0 0.00169466 3.3 0.00169458 3.3 0.00169468 0 0.0016945999999999999 0 0.0016947 3.3 0.00169462 3.3 0.00169472 0 0.0016946399999999999 0 0.00169474 3.3 0.00169466 3.3 0.00169476 0 0.0016946799999999998 0 0.00169478 3.3 0.0016947 3.3 0.0016948 0 0.0016947199999999998 0 0.0016948199999999999 3.3 0.00169474 3.3 0.00169484 0 0.00169476 0 0.00169486 3.3 0.00169478 3.3 0.00169488 0 0.0016948 0 0.0016949 3.3 0.0016948199999999999 3.3 0.00169492 0 0.00169484 0 0.00169494 3.3 0.0016948599999999999 3.3 0.00169496 0 0.00169488 0 0.00169498 3.3 0.0016948999999999998 3.3 0.001695 0 0.00169492 0 0.00169502 3.3 0.0016949399999999998 3.3 0.0016950399999999999 0 0.00169496 0 0.00169506 3.3 0.00169498 3.3 0.00169508 0 0.001695 0 0.0016951 3.3 0.00169502 3.3 0.00169512 0 0.0016950399999999999 0 0.00169514 3.3 0.00169506 3.3 0.00169516 0 0.0016950799999999999 0 0.00169518 3.3 0.0016951 3.3 0.0016952 0 0.0016951199999999998 0 0.0016952199999999999 3.3 0.00169514 3.3 0.00169524 0 0.0016951599999999998 0 0.0016952599999999999 3.3 0.00169518 3.3 0.00169528 0 0.0016952 0 0.0016953 3.3 0.0016952199999999999 3.3 0.00169532 0 0.00169524 0 0.00169534 3.3 0.0016952599999999999 3.3 0.00169536 0 0.00169528 0 0.00169538 3.3 0.0016952999999999998 3.3 0.0016954 0 0.00169532 0 0.00169542 3.3 0.0016953399999999998 3.3 0.0016954399999999999 0 0.00169536 0 0.00169546 3.3 0.0016953799999999998 3.3 0.0016954799999999999 0 0.0016954 0 0.0016955 3.3 0.00169542 3.3 0.00169552 0 0.0016954399999999999 0 0.00169554 3.3 0.00169546 3.3 0.00169556 0 0.0016954799999999999 0 0.00169558 3.3 0.0016955 3.3 0.0016956 0 0.0016955199999999998 0 0.00169562 3.3 0.00169554 3.3 0.00169564 0 0.0016955599999999998 0 0.0016956599999999999 3.3 0.00169558 3.3 0.00169568 0 0.0016956 0 0.0016957 3.3 0.00169562 3.3 0.00169572 0 0.00169564 0 0.00169574 3.3 0.0016956599999999999 3.3 0.00169576 0 0.00169568 0 0.00169578 3.3 0.0016956999999999999 3.3 0.0016958 0 0.00169572 0 0.00169582 3.3 0.0016957399999999998 3.3 0.0016958399999999999 0 0.00169576 0 0.00169586 3.3 0.0016957799999999998 3.3 0.0016958799999999999 0 0.0016958 0 0.0016959 3.3 0.00169582 3.3 0.00169592 0 0.0016958399999999999 0 0.00169594 3.3 0.00169586 3.3 0.00169596 0 0.0016958799999999999 0 0.00169598 3.3 0.0016959 3.3 0.001696 0 0.0016959199999999998 0 0.00169602 3.3 0.00169594 3.3 0.00169604 0 0.0016959599999999998 0 0.0016960599999999999 3.3 0.00169598 3.3 0.00169608 0 0.0016959999999999998 0 0.0016960999999999999 3.3 0.00169602 3.3 0.00169612 0 0.00169604 0 0.00169614 3.3 0.0016960599999999999 3.3 0.00169616 0 0.00169608 0 0.00169618 3.3 0.0016960999999999999 3.3 0.0016962 0 0.00169612 0 0.00169622 3.3 0.0016961399999999998 3.3 0.00169624 0 0.00169616 0 0.00169626 3.3 0.0016961799999999998 3.3 0.0016962799999999999 0 0.0016962 0 0.0016963 3.3 0.0016962199999999998 3.3 0.0016963199999999999 0 0.00169624 0 0.00169634 3.3 0.00169626 3.3 0.00169636 0 0.0016962799999999999 0 0.00169638 3.3 0.0016963 3.3 0.0016964 0 0.0016963199999999999 0 0.00169642 3.3 0.00169634 3.3 0.00169644 0 0.0016963599999999998 0 0.00169646 3.3 0.00169638 3.3 0.00169648 0 0.0016963999999999998 0 0.0016964999999999999 3.3 0.00169642 3.3 0.00169652 0 0.00169644 0 0.00169654 3.3 0.00169646 3.3 0.00169656 0 0.00169648 0 0.00169658 3.3 0.0016964999999999999 3.3 0.0016966 0 0.00169652 0 0.00169662 3.3 0.0016965399999999999 3.3 0.00169664 0 0.00169656 0 0.00169666 3.3 0.0016965799999999998 3.3 0.0016966799999999999 0 0.0016966 0 0.0016967 3.3 0.0016966199999999998 3.3 0.0016967199999999999 0 0.00169664 0 0.00169674 3.3 0.00169666 3.3 0.00169676 0 0.0016966799999999999 0 0.00169678 3.3 0.0016967 3.3 0.0016968 0 0.0016967199999999999 0 0.00169682 3.3 0.00169674 3.3 0.00169684 0 0.0016967599999999998 0 0.00169686 3.3 0.00169678 3.3 0.00169688 0 0.0016967999999999998 0 0.0016968999999999999 3.3 0.00169682 3.3 0.00169692 0 0.0016968399999999998 0 0.0016969399999999999 3.3 0.00169686 3.3 0.00169696 0 0.00169688 0 0.00169698 3.3 0.0016968999999999999 3.3 0.001697 0 0.00169692 0 0.00169702 3.3 0.0016969399999999999 3.3 0.00169704 0 0.00169696 0 0.00169706 3.3 0.0016969799999999998 3.3 0.00169708 0 0.001697 0 0.0016971 3.3 0.0016970199999999998 3.3 0.0016971199999999999 0 0.00169704 0 0.00169714 3.3 0.0016970599999999998 3.3 0.0016971599999999999 0 0.00169708 0 0.00169718 3.3 0.0016971 3.3 0.0016972 0 0.0016971199999999999 0 0.00169722 3.3 0.00169714 3.3 0.00169724 0 0.0016971599999999999 0 0.00169726 3.3 0.00169718 3.3 0.00169728 0 0.0016971999999999998 0 0.0016973 3.3 0.00169722 3.3 0.00169732 0 0.0016972399999999998 0 0.0016973399999999999 3.3 0.00169726 3.3 0.00169736 0 0.00169728 0 0.00169738 3.3 0.0016973 3.3 0.0016974 0 0.00169732 0 0.00169742 3.3 0.0016973399999999999 3.3 0.00169744 0 0.00169736 0 0.00169746 3.3 0.0016973799999999999 3.3 0.00169748 0 0.0016974 0 0.0016975 3.3 0.0016974199999999998 3.3 0.0016975199999999999 0 0.00169744 0 0.00169754 3.3 0.0016974599999999998 3.3 0.0016975599999999999 0 0.00169748 0 0.00169758 3.3 0.0016975 3.3 0.0016976 0 0.0016975199999999999 0 0.00169762 3.3 0.00169754 3.3 0.00169764 0 0.0016975599999999999 0 0.00169766 3.3 0.00169758 3.3 0.00169768 0 0.0016975999999999998 0 0.0016977 3.3 0.00169762 3.3 0.00169772 0 0.0016976399999999998 0 0.0016977399999999999 3.3 0.00169766 3.3 0.00169776 0 0.0016976799999999998 0 0.0016977799999999999 3.3 0.0016977 3.3 0.0016978 0 0.00169772 0 0.00169782 3.3 0.0016977399999999999 3.3 0.00169784 0 0.00169776 0 0.00169786 3.3 0.0016977799999999999 3.3 0.00169788 0 0.0016978 0 0.0016979 3.3 0.0016978199999999998 3.3 0.00169792 0 0.00169784 0 0.00169794 3.3 0.0016978599999999998 3.3 0.0016979599999999999 0 0.00169788 0 0.00169798 3.3 0.0016979 3.3 0.001698 0 0.00169792 0 0.00169802 3.3 0.00169794 3.3 0.00169804 0 0.0016979599999999999 0 0.00169806 3.3 0.00169798 3.3 0.00169808 0 0.0016979999999999999 0 0.0016981 3.3 0.00169802 3.3 0.00169812 0 0.0016980399999999998 0 0.00169814 3.3 0.00169806 3.3 0.00169816 0 0.0016980799999999998 0 0.0016981799999999999 3.3 0.0016981 3.3 0.0016982 0 0.00169812 0 0.00169822 3.3 0.00169814 3.3 0.00169824 0 0.00169816 0 0.00169826 3.3 0.0016981799999999999 3.3 0.00169828 0 0.0016982 0 0.0016983 3.3 0.0016982199999999999 3.3 0.00169832 0 0.00169824 0 0.00169834 3.3 0.0016982599999999998 3.3 0.0016983599999999999 0 0.00169828 0 0.00169838 3.3 0.0016982999999999998 3.3 0.0016983999999999999 0 0.00169832 0 0.00169842 3.3 0.00169834 3.3 0.00169844 0 0.0016983599999999999 0 0.00169846 3.3 0.00169838 3.3 0.00169848 0 0.0016983999999999999 0 0.0016985 3.3 0.00169842 3.3 0.00169852 0 0.0016984399999999998 0 0.00169854 3.3 0.00169846 3.3 0.00169856 0 0.0016984799999999998 0 0.0016985799999999999 3.3 0.0016985 3.3 0.0016986 0 0.0016985199999999998 0 0.0016986199999999999 3.3 0.00169854 3.3 0.00169864 0 0.00169856 0 0.00169866 3.3 0.0016985799999999999 3.3 0.00169868 0 0.0016986 0 0.0016987 3.3 0.0016986199999999999 3.3 0.00169872 0 0.00169864 0 0.00169874 3.3 0.0016986599999999998 3.3 0.00169876 0 0.00169868 0 0.00169878 3.3 0.0016986999999999998 3.3 0.0016987999999999999 0 0.00169872 0 0.00169882 3.3 0.00169874 3.3 0.00169884 0 0.00169876 0 0.00169886 3.3 0.00169878 3.3 0.00169888 0 0.0016987999999999999 0 0.0016989 3.3 0.00169882 3.3 0.00169892 0 0.0016988399999999999 0 0.00169894 3.3 0.00169886 3.3 0.00169896 0 0.0016988799999999998 0 0.0016989799999999999 3.3 0.0016989 3.3 0.001699 0 0.0016989199999999998 0 0.0016990199999999999 3.3 0.00169894 3.3 0.00169904 0 0.00169896 0 0.00169906 3.3 0.0016989799999999999 3.3 0.00169908 0 0.001699 0 0.0016991 3.3 0.0016990199999999999 3.3 0.00169912 0 0.00169904 0 0.00169914 3.3 0.0016990599999999998 3.3 0.00169916 0 0.00169908 0 0.00169918 3.3 0.0016990999999999998 3.3 0.0016991999999999999 0 0.00169912 0 0.00169922 3.3 0.0016991399999999998 3.3 0.0016992399999999999 0 0.00169916 0 0.00169926 3.3 0.00169918 3.3 0.00169928 0 0.0016991999999999999 0 0.0016993 3.3 0.00169922 3.3 0.00169932 0 0.0016992399999999999 0 0.00169934 3.3 0.00169926 3.3 0.00169936 0 0.0016992799999999998 0 0.00169938 3.3 0.0016993 3.3 0.0016994 0 0.0016993199999999998 0 0.0016994199999999999 3.3 0.00169934 3.3 0.00169944 0 0.0016993599999999998 0 0.0016994599999999999 3.3 0.00169938 3.3 0.00169948 0 0.0016994 0 0.0016995 3.3 0.0016994199999999999 3.3 0.00169952 0 0.00169944 0 0.00169954 3.3 0.0016994599999999999 3.3 0.00169956 0 0.00169948 0 0.00169958 3.3 0.0016994999999999998 3.3 0.0016996 0 0.00169952 0 0.00169962 3.3 0.0016995399999999998 3.3 0.0016996399999999999 0 0.00169956 0 0.00169966 3.3 0.00169958 3.3 0.00169968 0 0.0016996 0 0.0016997 3.3 0.00169962 3.3 0.00169972 0 0.0016996399999999999 0 0.00169974 3.3 0.00169966 3.3 0.00169976 0 0.0016996799999999999 0 0.00169978 3.3 0.0016997 3.3 0.0016998 0 0.0016997199999999998 0 0.0016998199999999999 3.3 0.00169974 3.3 0.00169984 0 0.0016997599999999998 0 0.0016998599999999999 3.3 0.00169978 3.3 0.00169988 0 0.0016998 0 0.0016999 3.3 0.0016998199999999999 3.3 0.00169992 0 0.00169984 0 0.00169994 3.3 0.0016998599999999999 3.3 0.00169996 0 0.00169988 0 0.00169998 3.3 0.0016998999999999998 3.3 0.0017 0 0.00169992 0 0.00170002 3.3 0.0016999399999999998 3.3 0.0017000399999999999 0 0.00169996 0 0.00170006 3.3 0.0016999799999999998 3.3 0.0017000799999999999 0 0.0017 0 0.0017001 3.3 0.00170002 3.3 0.00170012 0 0.0017000399999999999 0 0.00170014 3.3 0.00170006 3.3 0.00170016 0 0.0017000799999999999 0 0.00170018 3.3 0.0017001 3.3 0.0017002 0 0.0017001199999999998 0 0.00170022 3.3 0.00170014 3.3 0.00170024 0 0.0017001599999999998 0 0.0017002599999999999 3.3 0.00170018 3.3 0.00170028 0 0.0017001999999999998 0 0.0017002999999999999 3.3 0.00170022 3.3 0.00170032 0 0.00170024 0 0.00170034 3.3 0.0017002599999999999 3.3 0.00170036 0 0.00170028 0 0.00170038 3.3 0.0017002999999999999 3.3 0.0017004 0 0.00170032 0 0.00170042 3.3 0.0017003399999999998 3.3 0.00170044 0 0.00170036 0 0.00170046 3.3 0.0017003799999999998 3.3 0.0017004799999999999 0 0.0017004 0 0.0017005 3.3 0.00170042 3.3 0.00170052 0 0.00170044 0 0.00170054 3.3 0.00170046 3.3 0.00170056 0 0.0017004799999999999 0 0.00170058 3.3 0.0017005 3.3 0.0017006 0 0.0017005199999999999 0 0.00170062 3.3 0.00170054 3.3 0.00170064 0 0.0017005599999999998 0 0.0017006599999999999 3.3 0.00170058 3.3 0.00170068 0 0.0017005999999999998 0 0.0017006999999999999 3.3 0.00170062 3.3 0.00170072 0 0.00170064 0 0.00170074 3.3 0.0017006599999999999 3.3 0.00170076 0 0.00170068 0 0.00170078 3.3 0.0017006999999999999 3.3 0.0017008 0 0.00170072 0 0.00170082 3.3 0.0017007399999999998 3.3 0.00170084 0 0.00170076 0 0.00170086 3.3 0.0017007799999999998 3.3 0.0017008799999999999 0 0.0017008 0 0.0017009 3.3 0.0017008199999999998 3.3 0.0017009199999999999 0 0.00170084 0 0.00170094 3.3 0.00170086 3.3 0.00170096 0 0.0017008799999999999 0 0.00170098 3.3 0.0017009 3.3 0.001701 0 0.0017009199999999999 0 0.00170102 3.3 0.00170094 3.3 0.00170104 0 0.0017009599999999998 0 0.00170106 3.3 0.00170098 3.3 0.00170108 0 0.0017009999999999998 0 0.0017010999999999999 3.3 0.00170102 3.3 0.00170112 0 0.00170104 0 0.00170114 3.3 0.00170106 3.3 0.00170116 0 0.00170108 0 0.00170118 3.3 0.0017010999999999999 3.3 0.0017012 0 0.00170112 0 0.00170122 3.3 0.0017011399999999999 3.3 0.00170124 0 0.00170116 0 0.00170126 3.3 0.0017011799999999998 3.3 0.00170128 0 0.0017012 0 0.0017013 3.3 0.0017012199999999998 3.3 0.0017013199999999999 0 0.00170124 0 0.00170134 3.3 0.00170126 3.3 0.00170136 0 0.00170128 0 0.00170138 3.3 0.0017013 3.3 0.0017014 0 0.0017013199999999999 0 0.00170142 3.3 0.00170134 3.3 0.00170144 0 0.0017013599999999999 0 0.00170146 3.3 0.00170138 3.3 0.00170148 0 0.0017013999999999998 0 0.0017014999999999999 3.3 0.00170142 3.3 0.00170152 0 0.0017014399999999998 0 0.0017015399999999999 3.3 0.00170146 3.3 0.00170156 0 0.00170148 0 0.00170158 3.3 0.0017014999999999999 3.3 0.0017016 0 0.00170152 0 0.00170162 3.3 0.0017015399999999999 3.3 0.00170164 0 0.00170156 0 0.00170166 3.3 0.0017015799999999998 3.3 0.00170168 0 0.0017016 0 0.0017017 3.3 0.0017016199999999998 3.3 0.0017017199999999999 0 0.00170164 0 0.00170174 3.3 0.0017016599999999998 3.3 0.0017017599999999999 0 0.00170168 0 0.00170178 3.3 0.0017017 3.3 0.0017018 0 0.0017017199999999999 0 0.00170182 3.3 0.00170174 3.3 0.00170184 0 0.0017017599999999999 0 0.00170186 3.3 0.00170178 3.3 0.00170188 0 0.0017017999999999998 0 0.0017019 3.3 0.00170182 3.3 0.00170192 0 0.0017018399999999998 0 0.0017019399999999999 3.3 0.00170186 3.3 0.00170196 0 0.00170188 0 0.00170198 3.3 0.0017019 3.3 0.001702 0 0.00170192 0 0.00170202 3.3 0.0017019399999999999 3.3 0.00170204 0 0.00170196 0 0.00170206 3.3 0.0017019799999999999 3.3 0.00170208 0 0.001702 0 0.0017021 3.3 0.0017020199999999998 3.3 0.00170212 0 0.00170204 0 0.00170214 3.3 0.0017020599999999998 3.3 0.0017021599999999999 0 0.00170208 0 0.00170218 3.3 0.0017021 3.3 0.0017022 0 0.00170212 0 0.00170222 3.3 0.00170214 3.3 0.00170224 0 0.0017021599999999999 0 0.00170226 3.3 0.00170218 3.3 0.00170228 0 0.0017021999999999999 0 0.0017023 3.3 0.00170222 3.3 0.00170232 0 0.0017022399999999998 0 0.0017023399999999999 3.3 0.00170226 3.3 0.00170236 0 0.0017022799999999998 0 0.0017023799999999999 3.3 0.0017023 3.3 0.0017024 0 0.00170232 0 0.00170242 3.3 0.0017023399999999999 3.3 0.00170244 0 0.00170236 0 0.00170246 3.3 0.0017023799999999999 3.3 0.00170248 0 0.0017024 0 0.0017025 3.3 0.0017024199999999998 3.3 0.00170252 0 0.00170244 0 0.00170254 3.3 0.0017024599999999998 3.3 0.0017025599999999999 0 0.00170248 0 0.00170258 3.3 0.0017024999999999998 3.3 0.0017025999999999999 0 0.00170252 0 0.00170262 3.3 0.00170254 3.3 0.00170264 0 0.0017025599999999999 0 0.00170266 3.3 0.00170258 3.3 0.00170268 0 0.0017025999999999999 0 0.0017027 3.3 0.00170262 3.3 0.00170272 0 0.0017026399999999998 0 0.00170274 3.3 0.00170266 3.3 0.00170276 0 0.0017026799999999998 0 0.0017027799999999999 3.3 0.0017027 3.3 0.0017028 0 0.00170272 0 0.00170282 3.3 0.00170274 3.3 0.00170284 0 0.00170276 0 0.00170286 3.3 0.0017027799999999999 3.3 0.00170288 0 0.0017028 0 0.0017029 3.3 0.0017028199999999999 3.3 0.00170292 0 0.00170284 0 0.00170294 3.3 0.0017028599999999998 3.3 0.0017029599999999999 0 0.00170288 0 0.00170298 3.3 0.0017028999999999998 3.3 0.0017029999999999999 0 0.00170292 0 0.00170302 3.3 0.00170294 3.3 0.00170304 0 0.0017029599999999999 0 0.00170306 3.3 0.00170298 3.3 0.00170308 0 0.0017029999999999999 0 0.0017031 3.3 0.00170302 3.3 0.00170312 0 0.0017030399999999998 0 0.00170314 3.3 0.00170306 3.3 0.00170316 0 0.0017030799999999998 0 0.0017031799999999999 3.3 0.0017031 3.3 0.0017032 0 0.0017031199999999998 0 0.0017032199999999999 3.3 0.00170314 3.3 0.00170324 0 0.00170316 0 0.00170326 3.3 0.0017031799999999999 3.3 0.00170328 0 0.0017032 0 0.0017033 3.3 0.0017032199999999999 3.3 0.00170332 0 0.00170324 0 0.00170334 3.3 0.0017032599999999998 3.3 0.00170336 0 0.00170328 0 0.00170338 3.3 0.0017032999999999998 3.3 0.0017033999999999999 0 0.00170332 0 0.00170342 3.3 0.0017033399999999998 3.3 0.0017034399999999999 0 0.00170336 0 0.00170346 3.3 0.00170338 3.3 0.00170348 0 0.0017033999999999999 0 0.0017035 3.3 0.00170342 3.3 0.00170352 0 0.0017034399999999999 0 0.00170354 3.3 0.00170346 3.3 0.00170356 0 0.0017034799999999998 0 0.00170358 3.3 0.0017035 3.3 0.0017036 0 0.0017035199999999998 0 0.0017036199999999999 3.3 0.00170354 3.3 0.00170364 0 0.00170356 0 0.00170366 3.3 0.00170358 3.3 0.00170368 0 0.0017036 0 0.0017037 3.3 0.0017036199999999999 3.3 0.00170372 0 0.00170364 0 0.00170374 3.3 0.0017036599999999999 3.3 0.00170376 0 0.00170368 0 0.00170378 3.3 0.0017036999999999998 3.3 0.0017037999999999999 0 0.00170372 0 0.00170382 3.3 0.0017037399999999998 3.3 0.0017038399999999999 0 0.00170376 0 0.00170386 3.3 0.00170378 3.3 0.00170388 0 0.0017037999999999999 0 0.0017039 3.3 0.00170382 3.3 0.00170392 0 0.0017038399999999999 0 0.00170394 3.3 0.00170386 3.3 0.00170396 0 0.0017038799999999998 0 0.00170398 3.3 0.0017039 3.3 0.001704 0 0.0017039199999999998 0 0.0017040199999999999 3.3 0.00170394 3.3 0.00170404 0 0.0017039599999999998 0 0.0017040599999999999 3.3 0.00170398 3.3 0.00170408 0 0.001704 0 0.0017041 3.3 0.0017040199999999999 3.3 0.00170412 0 0.00170404 0 0.00170414 3.3 0.0017040599999999999 3.3 0.00170416 0 0.00170408 0 0.00170418 3.3 0.0017040999999999998 3.3 0.0017042 0 0.00170412 0 0.00170422 3.3 0.0017041399999999998 3.3 0.0017042399999999999 0 0.00170416 0 0.00170426 3.3 0.0017041799999999998 3.3 0.0017042799999999999 0 0.0017042 0 0.0017043 3.3 0.00170422 3.3 0.00170432 0 0.0017042399999999999 0 0.00170434 3.3 0.00170426 3.3 0.00170436 0 0.0017042799999999999 0 0.00170438 3.3 0.0017043 3.3 0.0017044 0 0.0017043199999999998 0 0.00170442 3.3 0.00170434 3.3 0.00170444 0 0.0017043599999999998 0 0.0017044599999999999 3.3 0.00170438 3.3 0.00170448 0 0.0017044 0 0.0017045 3.3 0.00170442 3.3 0.00170452 0 0.00170444 0 0.00170454 3.3 0.0017044599999999999 3.3 0.00170456 0 0.00170448 0 0.00170458 3.3 0.0017044999999999999 3.3 0.0017046 0 0.00170452 0 0.00170462 3.3 0.0017045399999999998 3.3 0.0017046399999999999 0 0.00170456 0 0.00170466 3.3 0.0017045799999999998 3.3 0.0017046799999999999 0 0.0017046 0 0.0017047 3.3 0.00170462 3.3 0.00170472 0 0.0017046399999999999 0 0.00170474 3.3 0.00170466 3.3 0.00170476 0 0.0017046799999999999 0 0.00170478 3.3 0.0017047 3.3 0.0017048 0 0.0017047199999999998 0 0.00170482 3.3 0.00170474 3.3 0.00170484 0 0.0017047599999999998 0 0.0017048599999999999 3.3 0.00170478 3.3 0.00170488 0 0.0017047999999999998 0 0.0017048999999999999 3.3 0.00170482 3.3 0.00170492 0 0.00170484 0 0.00170494 3.3 0.0017048599999999999 3.3 0.00170496 0 0.00170488 0 0.00170498 3.3 0.0017048999999999999 3.3 0.001705 0 0.00170492 0 0.00170502 3.3 0.0017049399999999998 3.3 0.00170504 0 0.00170496 0 0.00170506 3.3 0.0017049799999999998 3.3 0.0017050799999999999 0 0.001705 0 0.0017051 3.3 0.00170502 3.3 0.00170512 0 0.00170504 0 0.00170514 3.3 0.00170506 3.3 0.00170516 0 0.0017050799999999999 0 0.00170518 3.3 0.0017051 3.3 0.0017052 0 0.0017051199999999999 0 0.00170522 3.3 0.00170514 3.3 0.00170524 0 0.0017051599999999998 0 0.00170526 3.3 0.00170518 3.3 0.00170528 0 0.0017051999999999998 0 0.0017052999999999999 3.3 0.00170522 3.3 0.00170532 0 0.00170524 0 0.00170534 3.3 0.00170526 3.3 0.00170536 0 0.00170528 0 0.00170538 3.3 0.0017052999999999999 3.3 0.0017054 0 0.00170532 0 0.00170542 3.3 0.0017053399999999999 3.3 0.00170544 0 0.00170536 0 0.00170546 3.3 0.0017053799999999998 3.3 0.0017054799999999999 0 0.0017054 0 0.0017055 3.3 0.0017054199999999998 3.3 0.0017055199999999999 0 0.00170544 0 0.00170554 3.3 0.00170546 3.3 0.00170556 0 0.0017054799999999999 0 0.00170558 3.3 0.0017055 3.3 0.0017056 0 0.0017055199999999999 0 0.00170562 3.3 0.00170554 3.3 0.00170564 0 0.0017055599999999998 0 0.00170566 3.3 0.00170558 3.3 0.00170568 0 0.0017055999999999998 0 0.0017056999999999999 3.3 0.00170562 3.3 0.00170572 0 0.0017056399999999998 0 0.0017057399999999999 3.3 0.00170566 3.3 0.00170576 0 0.00170568 0 0.00170578 3.3 0.0017056999999999999 3.3 0.0017058 0 0.00170572 0 0.00170582 3.3 0.0017057399999999999 3.3 0.00170584 0 0.00170576 0 0.00170586 3.3 0.0017057799999999998 3.3 0.00170588 0 0.0017058 0 0.0017059 3.3 0.0017058199999999998 3.3 0.0017059199999999999 0 0.00170584 0 0.00170594 3.3 0.00170586 3.3 0.00170596 0 0.00170588 0 0.00170598 3.3 0.0017059 3.3 0.001706 0 0.0017059199999999999 0 0.00170602 3.3 0.00170594 3.3 0.00170604 0 0.0017059599999999999 0 0.00170606 3.3 0.00170598 3.3 0.00170608 0 0.0017059999999999998 0 0.0017060999999999999 3.3 0.00170602 3.3 0.00170612 0 0.0017060399999999998 0 0.0017061399999999999 3.3 0.00170606 3.3 0.00170616 0 0.00170608 0 0.00170618 3.3 0.0017060999999999999 3.3 0.0017062 0 0.00170612 0 0.00170622 3.3 0.0017061399999999999 3.3 0.00170624 0 0.00170616 0 0.00170626 3.3 0.0017061799999999998 3.3 0.00170628 0 0.0017062 0 0.0017063 3.3 0.0017062199999999998 3.3 0.0017063199999999999 0 0.00170624 0 0.00170634 3.3 0.0017062599999999998 3.3 0.0017063599999999999 0 0.00170628 0 0.00170638 3.3 0.0017063 3.3 0.0017064 0 0.0017063199999999999 0 0.00170642 3.3 0.00170634 3.3 0.00170644 0 0.0017063599999999999 0 0.00170646 3.3 0.00170638 3.3 0.00170648 0 0.0017063999999999998 0 0.0017065 3.3 0.00170642 3.3 0.00170652 0 0.0017064399999999998 0 0.0017065399999999999 3.3 0.00170646 3.3 0.00170656 0 0.0017064799999999998 0 0.0017065799999999999 3.3 0.0017065 3.3 0.0017066 0 0.00170652 0 0.00170662 3.3 0.0017065399999999999 3.3 0.00170664 0 0.00170656 0 0.00170666 3.3 0.0017065799999999999 3.3 0.00170668 0 0.0017066 0 0.0017067 3.3 0.0017066199999999998 3.3 0.00170672 0 0.00170664 0 0.00170674 3.3 0.0017066599999999998 3.3 0.0017067599999999999 0 0.00170668 0 0.00170678 3.3 0.0017067 3.3 0.0017068 0 0.00170672 0 0.00170682 3.3 0.00170674 3.3 0.00170684 0 0.0017067599999999999 0 0.00170686 3.3 0.00170678 3.3 0.00170688 0 0.0017067999999999999 0 0.0017069 3.3 0.00170682 3.3 0.00170692 0 0.0017068399999999998 0 0.0017069399999999999 3.3 0.00170686 3.3 0.00170696 0 0.0017068799999999998 0 0.0017069799999999999 3.3 0.0017069 3.3 0.001707 0 0.00170692 0 0.00170702 3.3 0.0017069399999999999 3.3 0.00170704 0 0.00170696 0 0.00170706 3.3 0.0017069799999999999 3.3 0.00170708 0 0.001707 0 0.0017071 3.3 0.0017070199999999998 3.3 0.00170712 0 0.00170704 0 0.00170714 3.3 0.0017070599999999998 3.3 0.0017071599999999999 0 0.00170708 0 0.00170718 3.3 0.0017070999999999998 3.3 0.0017071999999999999 0 0.00170712 0 0.00170722 3.3 0.00170714 3.3 0.00170724 0 0.0017071599999999999 0 0.00170726 3.3 0.00170718 3.3 0.00170728 0 0.0017071999999999999 0 0.0017073 3.3 0.00170722 3.3 0.00170732 0 0.0017072399999999998 0 0.00170734 3.3 0.00170726 3.3 0.00170736 0 0.0017072799999999998 0 0.0017073799999999999 3.3 0.0017073 3.3 0.0017074 0 0.0017073199999999998 0 0.0017074199999999999 3.3 0.00170734 3.3 0.00170744 0 0.00170736 0 0.00170746 3.3 0.0017073799999999999 3.3 0.00170748 0 0.0017074 0 0.0017075 3.3 0.0017074199999999999 3.3 0.00170752 0 0.00170744 0 0.00170754 3.3 0.0017074599999999998 3.3 0.00170756 0 0.00170748 0 0.00170758 3.3 0.0017074999999999998 3.3 0.0017075999999999999 0 0.00170752 0 0.00170762 3.3 0.00170754 3.3 0.00170764 0 0.00170756 0 0.00170766 3.3 0.00170758 3.3 0.00170768 0 0.0017075999999999999 0 0.0017077 3.3 0.00170762 3.3 0.00170772 0 0.0017076399999999999 0 0.00170774 3.3 0.00170766 3.3 0.00170776 0 0.0017076799999999998 0 0.0017077799999999999 3.3 0.0017077 3.3 0.0017078 0 0.0017077199999999998 0 0.0017078199999999999 3.3 0.00170774 3.3 0.00170784 0 0.00170776 0 0.00170786 3.3 0.0017077799999999999 3.3 0.00170788 0 0.0017078 0 0.0017079 3.3 0.0017078199999999999 3.3 0.00170792 0 0.00170784 0 0.00170794 3.3 0.0017078599999999998 3.3 0.00170796 0 0.00170788 0 0.00170798 3.3 0.0017078999999999998 3.3 0.0017079999999999999 0 0.00170792 0 0.00170802 3.3 0.0017079399999999998 3.3 0.0017080399999999999 0 0.00170796 0 0.00170806 3.3 0.00170798 3.3 0.00170808 0 0.0017079999999999999 0 0.0017081 3.3 0.00170802 3.3 0.00170812 0 0.0017080399999999999 0 0.00170814 3.3 0.00170806 3.3 0.00170816 0 0.0017080799999999998 0 0.00170818 3.3 0.0017081 3.3 0.0017082 0 0.0017081199999999998 0 0.0017082199999999999 3.3 0.00170814 3.3 0.00170824 0 0.00170816 0 0.00170826 3.3 0.00170818 3.3 0.00170828 0 0.0017082 0 0.0017083 3.3 0.0017082199999999999 3.3 0.00170832 0 0.00170824 0 0.00170834 3.3 0.0017082599999999999 3.3 0.00170836 0 0.00170828 0 0.00170838 3.3 0.0017082999999999998 3.3 0.0017084 0 0.00170832 0 0.00170842 3.3 0.0017083399999999998 3.3 0.0017084399999999999 0 0.00170836 0 0.00170846 3.3 0.00170838 3.3 0.00170848 0 0.0017084 0 0.0017085 3.3 0.00170842 3.3 0.00170852 0 0.0017084399999999999 0 0.00170854 3.3 0.00170846 3.3 0.00170856 0 0.0017084799999999999 0 0.00170858 3.3 0.0017085 3.3 0.0017086 0 0.0017085199999999998 0 0.0017086199999999999 3.3 0.00170854 3.3 0.00170864 0 0.0017085599999999998 0 0.0017086599999999999 3.3 0.00170858 3.3 0.00170868 0 0.0017086 0 0.0017087 3.3 0.0017086199999999999 3.3 0.00170872 0 0.00170864 0 0.00170874 3.3 0.0017086599999999999 3.3 0.00170876 0 0.00170868 0 0.00170878 3.3 0.0017086999999999998 3.3 0.0017088 0 0.00170872 0 0.00170882 3.3 0.0017087399999999998 3.3 0.0017088399999999999 0 0.00170876 0 0.00170886 3.3 0.0017087799999999998 3.3 0.0017088799999999999 0 0.0017088 0 0.0017089 3.3 0.00170882 3.3 0.00170892 0 0.0017088399999999999 0 0.00170894 3.3 0.00170886 3.3 0.00170896 0 0.0017088799999999999 0 0.00170898 3.3 0.0017089 3.3 0.001709 0 0.0017089199999999998 0 0.00170902 3.3 0.00170894 3.3 0.00170904 0 0.0017089599999999998 0 0.0017090599999999999 3.3 0.00170898 3.3 0.00170908 0 0.001709 0 0.0017091 3.3 0.00170902 3.3 0.00170912 0 0.00170904 0 0.00170914 3.3 0.0017090599999999999 3.3 0.00170916 0 0.00170908 0 0.00170918 3.3 0.0017090999999999999 3.3 0.0017092 0 0.00170912 0 0.00170922 3.3 0.0017091399999999998 3.3 0.0017092399999999999 0 0.00170916 0 0.00170926 3.3 0.0017091799999999998 3.3 0.0017092799999999999 0 0.0017092 0 0.0017093 3.3 0.00170922 3.3 0.00170932 0 0.0017092399999999999 0 0.00170934 3.3 0.00170926 3.3 0.00170936 0 0.0017092799999999999 0 0.00170938 3.3 0.0017093 3.3 0.0017094 0 0.0017093199999999998 0 0.00170942 3.3 0.00170934 3.3 0.00170944 0 0.0017093599999999998 0 0.0017094599999999999 3.3 0.00170938 3.3 0.00170948 0 0.0017093999999999998 0 0.0017094999999999999 3.3 0.00170942 3.3 0.00170952 0 0.00170944 0 0.00170954 3.3 0.0017094599999999999 3.3 0.00170956 0 0.00170948 0 0.00170958 3.3 0.0017094999999999999 3.3 0.0017096 0 0.00170952 0 0.00170962 3.3 0.0017095399999999998 3.3 0.00170964 0 0.00170956 0 0.00170966 3.3 0.0017095799999999998 3.3 0.0017096799999999999 0 0.0017096 0 0.0017097 3.3 0.0017096199999999998 3.3 0.0017097199999999999 0 0.00170964 0 0.00170974 3.3 0.00170966 3.3 0.00170976 0 0.0017096799999999999 0 0.00170978 3.3 0.0017097 3.3 0.0017098 0 0.0017097199999999999 0 0.00170982 3.3 0.00170974 3.3 0.00170984 0 0.0017097599999999998 0 0.00170986 3.3 0.00170978 3.3 0.00170988 0 0.0017097999999999998 0 0.0017098999999999999 3.3 0.00170982 3.3 0.00170992 0 0.00170984 0 0.00170994 3.3 0.00170986 3.3 0.00170996 0 0.00170988 0 0.00170998 3.3 0.0017098999999999999 3.3 0.00171 0 0.00170992 0 0.00171002 3.3 0.0017099399999999999 3.3 0.00171004 0 0.00170996 0 0.00171006 3.3 0.0017099799999999998 3.3 0.0017100799999999999 0 0.00171 0 0.0017101 3.3 0.0017100199999999998 3.3 0.0017101199999999999 0 0.00171004 0 0.00171014 3.3 0.00171006 3.3 0.00171016 0 0.0017100799999999999 0 0.00171018 3.3 0.0017101 3.3 0.0017102 0 0.0017101199999999999 0 0.00171022 3.3 0.00171014 3.3 0.00171024 0 0.0017101599999999998 0 0.00171026 3.3 0.00171018 3.3 0.00171028 0 0.0017101999999999998 0 0.0017102999999999999 3.3 0.00171022 3.3 0.00171032 0 0.0017102399999999998 0 0.0017103399999999999 3.3 0.00171026 3.3 0.00171036 0 0.00171028 0 0.00171038 3.3 0.0017102999999999999 3.3 0.0017104 0 0.00171032 0 0.00171042 3.3 0.0017103399999999999 3.3 0.00171044 0 0.00171036 0 0.00171046 3.3 0.0017103799999999998 3.3 0.00171048 0 0.0017104 0 0.0017105 3.3 0.0017104199999999998 3.3 0.0017105199999999999 0 0.00171044 0 0.00171054 3.3 0.0017104599999999998 3.3 0.0017105599999999999 0 0.00171048 0 0.00171058 3.3 0.0017105 3.3 0.0017106 0 0.0017105199999999999 0 0.00171062 3.3 0.00171054 3.3 0.00171064 0 0.0017105599999999999 0 0.00171066 3.3 0.00171058 3.3 0.00171068 0 0.0017105999999999998 0 0.0017107 3.3 0.00171062 3.3 0.00171072 0 0.0017106399999999998 0 0.0017107399999999999 3.3 0.00171066 3.3 0.00171076 0 0.00171068 0 0.00171078 3.3 0.0017107 3.3 0.0017108 0 0.00171072 0 0.00171082 3.3 0.0017107399999999999 3.3 0.00171084 0 0.00171076 0 0.00171086 3.3 0.0017107799999999999 3.3 0.00171088 0 0.0017108 0 0.0017109 3.3 0.0017108199999999998 3.3 0.0017109199999999999 0 0.00171084 0 0.00171094 3.3 0.0017108599999999998 3.3 0.0017109599999999999 0 0.00171088 0 0.00171098 3.3 0.0017109 3.3 0.001711 0 0.0017109199999999999 0 0.00171102 3.3 0.00171094 3.3 0.00171104 0 0.0017109599999999999 0 0.00171106 3.3 0.00171098 3.3 0.00171108 0 0.0017109999999999998 0 0.0017111 3.3 0.00171102 3.3 0.00171112 0 0.0017110399999999998 0 0.0017111399999999999 3.3 0.00171106 3.3 0.00171116 0 0.0017110799999999998 0 0.0017111799999999999 3.3 0.0017111 3.3 0.0017112 0 0.00171112 0 0.00171122 3.3 0.0017111399999999999 3.3 0.00171124 0 0.00171116 0 0.00171126 3.3 0.0017111799999999999 3.3 0.00171128 0 0.0017112 0 0.0017113 3.3 0.0017112199999999998 3.3 0.00171132 0 0.00171124 0 0.00171134 3.3 0.0017112599999999998 3.3 0.0017113599999999999 0 0.00171128 0 0.00171138 3.3 0.0017113 3.3 0.0017114 0 0.00171132 0 0.00171142 3.3 0.00171134 3.3 0.00171144 0 0.0017113599999999999 0 0.00171146 3.3 0.00171138 3.3 0.00171148 0 0.0017113999999999999 0 0.0017115 3.3 0.00171142 3.3 0.00171152 0 0.0017114399999999998 0 0.00171154 3.3 0.00171146 3.3 0.00171156 0 0.0017114799999999998 0 0.0017115799999999999 3.3 0.0017115 3.3 0.0017116 0 0.00171152 0 0.00171162 3.3 0.00171154 3.3 0.00171164 0 0.00171156 0 0.00171166 3.3 0.0017115799999999999 3.3 0.00171168 0 0.0017116 0 0.0017117 3.3 0.0017116199999999999 3.3 0.00171172 0 0.00171164 0 0.00171174 3.3 0.0017116599999999998 3.3 0.0017117599999999999 0 0.00171168 0 0.00171178 3.3 0.0017116999999999998 3.3 0.0017117999999999999 0 0.00171172 0 0.00171182 3.3 0.00171174 3.3 0.00171184 0 0.0017117599999999999 0 0.00171186 3.3 0.00171178 3.3 0.00171188 0 0.0017117999999999999 0 0.0017119 3.3 0.00171182 3.3 0.00171192 0 0.0017118399999999998 0 0.00171194 3.3 0.00171186 3.3 0.00171196 0 0.0017118799999999998 0 0.0017119799999999999 3.3 0.0017119 3.3 0.001712 0 0.0017119199999999998 0 0.0017120199999999999 3.3 0.00171194 3.3 0.00171204 0 0.00171196 0 0.00171206 3.3 0.0017119799999999999 3.3 0.00171208 0 0.001712 0 0.0017121 3.3 0.0017120199999999999 3.3 0.00171212 0 0.00171204 0 0.00171214 3.3 0.0017120599999999998 3.3 0.00171216 0 0.00171208 0 0.00171218 3.3 0.0017120999999999998 3.3 0.0017121999999999999 0 0.00171212 0 0.00171222 3.3 0.00171214 3.3 0.00171224 0 0.00171216 0 0.00171226 3.3 0.00171218 3.3 0.00171228 0 0.0017121999999999999 0 0.0017123 3.3 0.00171222 3.3 0.00171232 0 0.0017122399999999999 0 0.00171234 3.3 0.00171226 3.3 0.00171236 0 0.0017122799999999998 0 0.00171238 3.3 0.0017123 3.3 0.0017124 0 0.0017123199999999998 0 0.0017124199999999999 3.3 0.00171234 3.3 0.00171244 0 0.00171236 0 0.00171246 3.3 0.00171238 3.3 0.00171248 0 0.0017124 0 0.0017125 3.3 0.0017124199999999999 3.3 0.00171252 0 0.00171244 0 0.00171254 3.3 0.0017124599999999999 3.3 0.00171256 0 0.00171248 0 0.00171258 3.3 0.0017124999999999998 3.3 0.0017125999999999999 0 0.00171252 0 0.00171262 3.3 0.0017125399999999998 3.3 0.0017126399999999999 0 0.00171256 0 0.00171266 3.3 0.00171258 3.3 0.00171268 0 0.0017125999999999999 0 0.0017127 3.3 0.00171262 3.3 0.00171272 0 0.0017126399999999999 0 0.00171274 3.3 0.00171266 3.3 0.00171276 0 0.0017126799999999998 0 0.00171278 3.3 0.0017127 3.3 0.0017128 0 0.0017127199999999998 0 0.0017128199999999999 3.3 0.00171274 3.3 0.00171284 0 0.0017127599999999998 0 0.0017128599999999999 3.3 0.00171278 3.3 0.00171288 0 0.0017128 0 0.0017129 3.3 0.0017128199999999999 3.3 0.00171292 0 0.00171284 0 0.00171294 3.3 0.0017128599999999999 3.3 0.00171296 0 0.00171288 0 0.00171298 3.3 0.0017128999999999998 3.3 0.001713 0 0.00171292 0 0.00171302 3.3 0.0017129399999999998 3.3 0.0017130399999999999 0 0.00171296 0 0.00171306 3.3 0.00171298 3.3 0.00171308 0 0.001713 0 0.0017131 3.3 0.00171302 3.3 0.00171312 0 0.0017130399999999999 0 0.00171314 3.3 0.00171306 3.3 0.00171316 0 0.0017130799999999999 0 0.00171318 3.3 0.0017131 3.3 0.0017132 0 0.0017131199999999998 0 0.0017132199999999999 3.3 0.00171314 3.3 0.00171324 0 0.0017131599999999998 0 0.0017132599999999999 3.3 0.00171318 3.3 0.00171328 0 0.0017132 0 0.0017133 3.3 0.0017132199999999999 3.3 0.00171332 0 0.00171324 0 0.00171334 3.3 0.0017132599999999999 3.3 0.00171336 0 0.00171328 0 0.00171338 3.3 0.0017132999999999998 3.3 0.0017134 0 0.00171332 0 0.00171342 3.3 0.0017133399999999998 3.3 0.0017134399999999999 0 0.00171336 0 0.00171346 3.3 0.0017133799999999998 3.3 0.0017134799999999999 0 0.0017134 0 0.0017135 3.3 0.00171342 3.3 0.00171352 0 0.0017134399999999999 0 0.00171354 3.3 0.00171346 3.3 0.00171356 0 0.0017134799999999999 0 0.00171358 3.3 0.0017135 3.3 0.0017136 0 0.0017135199999999998 0 0.00171362 3.3 0.00171354 3.3 0.00171364 0 0.0017135599999999998 0 0.0017136599999999999 3.3 0.00171358 3.3 0.00171368 0 0.0017135999999999998 0 0.0017136999999999999 3.3 0.00171362 3.3 0.00171372 0 0.00171364 0 0.00171374 3.3 0.0017136599999999999 3.3 0.00171376 0 0.00171368 0 0.00171378 3.3 0.0017136999999999999 3.3 0.0017138 0 0.00171372 0 0.00171382 3.3 0.0017137399999999998 3.3 0.00171384 0 0.00171376 0 0.00171386 3.3 0.0017137799999999998 3.3 0.0017138799999999999 0 0.0017138 0 0.0017139 3.3 0.00171382 3.3 0.00171392 0 0.00171384 0 0.00171394 3.3 0.00171386 3.3 0.00171396 0 0.0017138799999999999 0 0.00171398 3.3 0.0017139 3.3 0.001714 0 0.0017139199999999999 0 0.00171402 3.3 0.00171394 3.3 0.00171404 0 0.0017139599999999998 0 0.0017140599999999999 3.3 0.00171398 3.3 0.00171408 0 0.0017139999999999998 0 0.0017140999999999999 3.3 0.00171402 3.3 0.00171412 0 0.00171404 0 0.00171414 3.3 0.0017140599999999999 3.3 0.00171416 0 0.00171408 0 0.00171418 3.3 0.0017140999999999999 3.3 0.0017142 0 0.00171412 0 0.00171422 3.3 0.0017141399999999998 3.3 0.00171424 0 0.00171416 0 0.00171426 3.3 0.0017141799999999998 3.3 0.0017142799999999999 0 0.0017142 0 0.0017143 3.3 0.0017142199999999998 3.3 0.0017143199999999999 0 0.00171424 0 0.00171434 3.3 0.00171426 3.3 0.00171436 0 0.0017142799999999999 0 0.00171438 3.3 0.0017143 3.3 0.0017144 0 0.0017143199999999999 0 0.00171442 3.3 0.00171434 3.3 0.00171444 0 0.0017143599999999998 0 0.00171446 3.3 0.00171438 3.3 0.00171448 0 0.0017143999999999998 0 0.0017144999999999999 3.3 0.00171442 3.3 0.00171452 0 0.0017144399999999998 0 0.0017145399999999999 3.3 0.00171446 3.3 0.00171456 0 0.00171448 0 0.00171458 3.3 0.0017144999999999999 3.3 0.0017146 0 0.00171452 0 0.00171462 3.3 0.0017145399999999999 3.3 0.00171464 0 0.00171456 0 0.00171466 3.3 0.0017145799999999998 3.3 0.00171468 0 0.0017146 0 0.0017147 3.3 0.0017146199999999998 3.3 0.0017147199999999999 0 0.00171464 0 0.00171474 3.3 0.00171466 3.3 0.00171476 0 0.00171468 0 0.00171478 3.3 0.0017147 3.3 0.0017148 0 0.0017147199999999999 0 0.00171482 3.3 0.00171474 3.3 0.00171484 0 0.0017147599999999999 0 0.00171486 3.3 0.00171478 3.3 0.00171488 0 0.0017147999999999998 0 0.0017148999999999999 3.3 0.00171482 3.3 0.00171492 0 0.0017148399999999998 0 0.0017149399999999999 3.3 0.00171486 3.3 0.00171496 0 0.00171488 0 0.00171498 3.3 0.0017148999999999999 3.3 0.001715 0 0.00171492 0 0.00171502 3.3 0.0017149399999999999 3.3 0.00171504 0 0.00171496 0 0.00171506 3.3 0.0017149799999999998 3.3 0.00171508 0 0.001715 0 0.0017151 3.3 0.0017150199999999998 3.3 0.0017151199999999999 0 0.00171504 0 0.00171514 3.3 0.0017150599999999998 3.3 0.0017151599999999999 0 0.00171508 0 0.00171518 3.3 0.0017151 3.3 0.0017152 0 0.0017151199999999999 0 0.00171522 3.3 0.00171514 3.3 0.00171524 0 0.0017151599999999999 0 0.00171526 3.3 0.00171518 3.3 0.00171528 0 0.0017151999999999998 0 0.0017153 3.3 0.00171522 3.3 0.00171532 0 0.0017152399999999998 0 0.0017153399999999999 3.3 0.00171526 3.3 0.00171536 0 0.00171528 0 0.00171538 3.3 0.0017153 3.3 0.0017154 0 0.00171532 0 0.00171542 3.3 0.0017153399999999999 3.3 0.00171544 0 0.00171536 0 0.00171546 3.3 0.0017153799999999999 3.3 0.00171548 0 0.0017154 0 0.0017155 3.3 0.0017154199999999998 3.3 0.00171552 0 0.00171544 0 0.00171554 3.3 0.0017154599999999998 3.3 0.0017155599999999999 0 0.00171548 0 0.00171558 3.3 0.0017155 3.3 0.0017156 0 0.00171552 0 0.00171562 3.3 0.00171554 3.3 0.00171564 0 0.0017155599999999999 0 0.00171566 3.3 0.00171558 3.3 0.00171568 0 0.0017155999999999999 0 0.0017157 3.3 0.00171562 3.3 0.00171572 0 0.0017156399999999998 0 0.0017157399999999999 3.3 0.00171566 3.3 0.00171576 0 0.0017156799999999998 0 0.0017157799999999999 3.3 0.0017157 3.3 0.0017158 0 0.00171572 0 0.00171582 3.3 0.0017157399999999999 3.3 0.00171584 0 0.00171576 0 0.00171586 3.3 0.0017157799999999999 3.3 0.00171588 0 0.0017158 0 0.0017159 3.3 0.0017158199999999998 3.3 0.00171592 0 0.00171584 0 0.00171594 3.3 0.0017158599999999998 3.3 0.0017159599999999999 0 0.00171588 0 0.00171598 3.3 0.0017158999999999998 3.3 0.0017159999999999999 0 0.00171592 0 0.00171602 3.3 0.00171594 3.3 0.00171604 0 0.0017159599999999999 0 0.00171606 3.3 0.00171598 3.3 0.00171608 0 0.0017159999999999999 0 0.0017161 3.3 0.00171602 3.3 0.00171612 0 0.0017160399999999998 0 0.00171614 3.3 0.00171606 3.3 0.00171616 0 0.0017160799999999998 0 0.0017161799999999999 3.3 0.0017161 3.3 0.0017162 0 0.00171612 0 0.00171622 3.3 0.00171614 3.3 0.00171624 0 0.00171616 0 0.00171626 3.3 0.0017161799999999999 3.3 0.00171628 0 0.0017162 0 0.0017163 3.3 0.0017162199999999999 3.3 0.00171632 0 0.00171624 0 0.00171634 3.3 0.0017162599999999998 3.3 0.0017163599999999999 0 0.00171628 0 0.00171638 3.3 0.0017162999999999998 3.3 0.0017163999999999999 0 0.00171632 0 0.00171642 3.3 0.00171634 3.3 0.00171644 0 0.0017163599999999999 0 0.00171646 3.3 0.00171638 3.3 0.00171648 0 0.0017163999999999999 0 0.0017165 3.3 0.00171642 3.3 0.00171652 0 0.0017164399999999998 0 0.00171654 3.3 0.00171646 3.3 0.00171656 0 0.0017164799999999998 0 0.0017165799999999999 3.3 0.0017165 3.3 0.0017166 0 0.0017165199999999998 0 0.0017166199999999999 3.3 0.00171654 3.3 0.00171664 0 0.00171656 0 0.00171666 3.3 0.0017165799999999999 3.3 0.00171668 0 0.0017166 0 0.0017167 3.3 0.0017166199999999999 3.3 0.00171672 0 0.00171664 0 0.00171674 3.3 0.0017166599999999998 3.3 0.00171676 0 0.00171668 0 0.00171678 3.3 0.0017166999999999998 3.3 0.0017167999999999999 0 0.00171672 0 0.00171682 3.3 0.0017167399999999998 3.3 0.0017168399999999999 0 0.00171676 0 0.00171686 3.3 0.00171678 3.3 0.00171688 0 0.0017167999999999999 0 0.0017169 3.3 0.00171682 3.3 0.00171692 0 0.0017168399999999999 0 0.00171694 3.3 0.00171686 3.3 0.00171696 0 0.0017168799999999998 0 0.00171698 3.3 0.0017169 3.3 0.001717 0 0.0017169199999999998 0 0.0017170199999999999 3.3 0.00171694 3.3 0.00171704 0 0.00171696 0 0.00171706 3.3 0.00171698 3.3 0.00171708 0 0.001717 0 0.0017171 3.3 0.0017170199999999999 3.3 0.00171712 0 0.00171704 0 0.00171714 3.3 0.0017170599999999999 3.3 0.00171716 0 0.00171708 0 0.00171718 3.3 0.0017170999999999998 3.3 0.0017171999999999999 0 0.00171712 0 0.00171722 3.3 0.0017171399999999998 3.3 0.0017172399999999999 0 0.00171716 0 0.00171726 3.3 0.00171718 3.3 0.00171728 0 0.0017171999999999999 0 0.0017173 3.3 0.00171722 3.3 0.00171732 0 0.0017172399999999999 0 0.00171734 3.3 0.00171726 3.3 0.00171736 0 0.0017172799999999998 0 0.00171738 3.3 0.0017173 3.3 0.0017174 0 0.0017173199999999998 0 0.0017174199999999999 3.3 0.00171734 3.3 0.00171744 0 0.0017173599999999998 0 0.0017174599999999999 3.3 0.00171738 3.3 0.00171748 0 0.0017174 0 0.0017175 3.3 0.0017174199999999999 3.3 0.00171752 0 0.00171744 0 0.00171754 3.3 0.0017174599999999999 3.3 0.00171756 0 0.00171748 0 0.00171758 3.3 0.0017174999999999998 3.3 0.0017176 0 0.00171752 0 0.00171762 3.3 0.0017175399999999998 3.3 0.0017176399999999999 0 0.00171756 0 0.00171766 3.3 0.0017175799999999998 3.3 0.0017176799999999999 0 0.0017176 0 0.0017177 3.3 0.00171762 3.3 0.00171772 0 0.0017176399999999999 0 0.00171774 3.3 0.00171766 3.3 0.00171776 0 0.0017176799999999999 0 0.00171778 3.3 0.0017177 3.3 0.0017178 0 0.0017177199999999998 0 0.00171782 3.3 0.00171774 3.3 0.00171784 0 0.0017177599999999998 0 0.0017178599999999999 3.3 0.00171778 3.3 0.00171788 0 0.0017178 0 0.0017179 3.3 0.00171782 3.3 0.00171792 0 0.00171784 0 0.00171794 3.3 0.0017178599999999999 3.3 0.00171796 0 0.00171788 0 0.00171798 3.3 0.0017178999999999999 3.3 0.001718 0 0.00171792 0 0.00171802 3.3 0.0017179399999999998 3.3 0.0017180399999999999 0 0.00171796 0 0.00171806 3.3 0.0017179799999999998 3.3 0.0017180799999999999 0 0.001718 0 0.0017181 3.3 0.00171802 3.3 0.00171812 0 0.0017180399999999999 0 0.00171814 3.3 0.00171806 3.3 0.00171816 0 0.0017180799999999999 0 0.00171818 3.3 0.0017181 3.3 0.0017182 0 0.0017181199999999998 0 0.00171822 3.3 0.00171814 3.3 0.00171824 0 0.0017181599999999998 0 0.0017182599999999999 3.3 0.00171818 3.3 0.00171828 0 0.0017181999999999998 0 0.0017182999999999999 3.3 0.00171822 3.3 0.00171832 0 0.00171824 0 0.00171834 3.3 0.0017182599999999999 3.3 0.00171836 0 0.00171828 0 0.00171838 3.3 0.0017182999999999999 3.3 0.0017184 0 0.00171832 0 0.00171842 3.3 0.0017183399999999998 3.3 0.00171844 0 0.00171836 0 0.00171846 3.3 0.0017183799999999998 3.3 0.0017184799999999999 0 0.0017184 0 0.0017185 3.3 0.00171842 3.3 0.00171852 0 0.00171844 0 0.00171854 3.3 0.00171846 3.3 0.00171856 0 0.0017184799999999999 0 0.00171858 3.3 0.0017185 3.3 0.0017186 0 0.0017185199999999999 0 0.00171862 3.3 0.00171854 3.3 0.00171864 0 0.0017185599999999998 0 0.00171866 3.3 0.00171858 3.3 0.00171868 0 0.0017185999999999998 0 0.0017186999999999999 3.3 0.00171862 3.3 0.00171872 0 0.00171864 0 0.00171874 3.3 0.00171866 3.3 0.00171876 0 0.00171868 0 0.00171878 3.3 0.0017186999999999999 3.3 0.0017188 0 0.00171872 0 0.00171882 3.3 0.0017187399999999999 3.3 0.00171884 0 0.00171876 0 0.00171886 3.3 0.0017187799999999998 3.3 0.0017188799999999999 0 0.0017188 0 0.0017189 3.3 0.0017188199999999998 3.3 0.0017189199999999999 0 0.00171884 0 0.00171894 3.3 0.00171886 3.3 0.00171896 0 0.0017188799999999999 0 0.00171898 3.3 0.0017189 3.3 0.001719 0 0.0017189199999999999 0 0.00171902 3.3 0.00171894 3.3 0.00171904 0 0.0017189599999999998 0 0.00171906 3.3 0.00171898 3.3 0.00171908 0 0.0017189999999999998 0 0.0017190999999999999 3.3 0.00171902 3.3 0.00171912 0 0.0017190399999999998 0 0.0017191399999999999 3.3 0.00171906 3.3 0.00171916 0 0.00171908 0 0.00171918 3.3 0.0017190999999999999 3.3 0.0017192 0 0.00171912 0 0.00171922 3.3 0.0017191399999999999 3.3 0.00171924 0 0.00171916 0 0.00171926 3.3 0.0017191799999999998 3.3 0.00171928 0 0.0017192 0 0.0017193 3.3 0.0017192199999999998 3.3 0.0017193199999999999 0 0.00171924 0 0.00171934 3.3 0.00171926 3.3 0.00171936 0 0.00171928 0 0.00171938 3.3 0.0017193 3.3 0.0017194 0 0.0017193199999999999 0 0.00171942 3.3 0.00171934 3.3 0.00171944 0 0.0017193599999999999 0 0.00171946 3.3 0.00171938 3.3 0.00171948 0 0.0017193999999999998 0 0.0017194999999999999 3.3 0.00171942 3.3 0.00171952 0 0.0017194399999999998 0 0.0017195399999999999 3.3 0.00171946 3.3 0.00171956 0 0.00171948 0 0.00171958 3.3 0.0017194999999999999 3.3 0.0017196 0 0.00171952 0 0.00171962 3.3 0.0017195399999999999 3.3 0.00171964 0 0.00171956 0 0.00171966 3.3 0.0017195799999999998 3.3 0.00171968 0 0.0017196 0 0.0017197 3.3 0.0017196199999999998 3.3 0.0017197199999999999 0 0.00171964 0 0.00171974 3.3 0.0017196599999999998 3.3 0.0017197599999999999 0 0.00171968 0 0.00171978 3.3 0.0017197 3.3 0.0017198 0 0.0017197199999999999 0 0.00171982 3.3 0.00171974 3.3 0.00171984 0 0.0017197599999999999 0 0.00171986 3.3 0.00171978 3.3 0.00171988 0 0.0017197999999999998 0 0.0017199 3.3 0.00171982 3.3 0.00171992 0 0.0017198399999999998 0 0.0017199399999999999 3.3 0.00171986 3.3 0.00171996 0 0.0017198799999999998 0 0.0017199799999999999 3.3 0.0017199 3.3 0.00172 0 0.00171992 0 0.00172002 3.3 0.0017199399999999999 3.3 0.00172004 0 0.00171996 0 0.00172006 3.3 0.0017199799999999999 3.3 0.00172008 0 0.00172 0 0.0017201 3.3 0.0017200199999999998 3.3 0.00172012 0 0.00172004 0 0.00172014 3.3 0.0017200599999999998 3.3 0.0017201599999999999 0 0.00172008 0 0.00172018 3.3 0.0017201 3.3 0.0017202 0 0.00172012 0 0.00172022 3.3 0.00172014 3.3 0.00172024 0 0.0017201599999999999 0 0.00172026 3.3 0.00172018 3.3 0.00172028 0 0.0017201999999999999 0 0.0017203 3.3 0.00172022 3.3 0.00172032 0 0.0017202399999999998 0 0.0017203399999999999 3.3 0.00172026 3.3 0.00172036 0 0.0017202799999999998 0 0.0017203799999999999 3.3 0.0017203 3.3 0.0017204 0 0.00172032 0 0.00172042 3.3 0.0017203399999999999 3.3 0.00172044 0 0.00172036 0 0.00172046 3.3 0.0017203799999999999 3.3 0.00172048 0 0.0017204 0 0.0017205 3.3 0.0017204199999999998 3.3 0.00172052 0 0.00172044 0 0.00172054 3.3 0.0017204599999999998 3.3 0.0017205599999999999 0 0.00172048 0 0.00172058 3.3 0.0017204999999999998 3.3 0.0017205999999999999 0 0.00172052 0 0.00172062 3.3 0.00172054 3.3 0.00172064 0 0.0017205599999999999 0 0.00172066 3.3 0.00172058 3.3 0.00172068 0 0.0017205999999999999 0 0.0017207 3.3 0.00172062 3.3 0.00172072 0 0.0017206399999999998 0 0.00172074 3.3 0.00172066 3.3 0.00172076 0 0.0017206799999999998 0 0.0017207799999999999 3.3 0.0017207 3.3 0.0017208 0 0.0017207199999999998 0 0.0017208199999999999 3.3 0.00172074 3.3 0.00172084 0 0.00172076 0 0.00172086 3.3 0.0017207799999999999 3.3 0.00172088 0 0.0017208 0 0.0017209 3.3 0.0017208199999999999 3.3 0.00172092 0 0.00172084 0 0.00172094 3.3 0.0017208599999999998 3.3 0.00172096 0 0.00172088 0 0.00172098 3.3 0.0017208999999999998 3.3 0.0017209999999999999 0 0.00172092 0 0.00172102 3.3 0.00172094 3.3 0.00172104 0 0.00172096 0 0.00172106 3.3 0.00172098 3.3 0.00172108 0 0.0017209999999999999 0 0.0017211 3.3 0.00172102 3.3 0.00172112 0 0.0017210399999999999 0 0.00172114 3.3 0.00172106 3.3 0.00172116 0 0.0017210799999999998 0 0.0017211799999999999 3.3 0.0017211 3.3 0.0017212 0 0.0017211199999999998 0 0.0017212199999999999 3.3 0.00172114 3.3 0.00172124 0 0.00172116 0 0.00172126 3.3 0.0017211799999999999 3.3 0.00172128 0 0.0017212 0 0.0017213 3.3 0.0017212199999999999 3.3 0.00172132 0 0.00172124 0 0.00172134 3.3 0.0017212599999999998 3.3 0.00172136 0 0.00172128 0 0.00172138 3.3 0.0017212999999999998 3.3 0.0017213999999999999 0 0.00172132 0 0.00172142 3.3 0.0017213399999999998 3.3 0.0017214399999999999 0 0.00172136 0 0.00172146 3.3 0.00172138 3.3 0.00172148 0 0.0017213999999999999 0 0.0017215 3.3 0.00172142 3.3 0.00172152 0 0.0017214399999999999 0 0.00172154 3.3 0.00172146 3.3 0.00172156 0 0.0017214799999999998 0 0.00172158 3.3 0.0017215 3.3 0.0017216 0 0.0017215199999999998 0 0.0017216199999999999 3.3 0.00172154 3.3 0.00172164 0 0.0017215599999999998 0 0.0017216599999999999 3.3 0.00172158 3.3 0.00172168 0 0.0017216 0 0.0017217 3.3 0.0017216199999999999 3.3 0.00172172 0 0.00172164 0 0.00172174 3.3 0.0017216599999999999 3.3 0.00172176 0 0.00172168 0 0.00172178 3.3 0.0017216999999999998 3.3 0.0017218 0 0.00172172 0 0.00172182 3.3 0.0017217399999999998 3.3 0.0017218399999999999 0 0.00172176 0 0.00172186 3.3 0.00172178 3.3 0.00172188 0 0.0017218 0 0.0017219 3.3 0.00172182 3.3 0.00172192 0 0.0017218399999999999 0 0.00172194 3.3 0.00172186 3.3 0.00172196 0 0.0017218799999999999 0 0.00172198 3.3 0.0017219 3.3 0.001722 0 0.0017219199999999998 0 0.0017220199999999999 3.3 0.00172194 3.3 0.00172204 0 0.0017219599999999998 0 0.0017220599999999999 3.3 0.00172198 3.3 0.00172208 0 0.001722 0 0.0017221 3.3 0.0017220199999999999 3.3 0.00172212 0 0.00172204 0 0.00172214 3.3 0.0017220599999999999 3.3 0.00172216 0 0.00172208 0 0.00172218 3.3 0.0017220999999999998 3.3 0.0017222 0 0.00172212 0 0.00172222 3.3 0.0017221399999999998 3.3 0.0017222399999999999 0 0.00172216 0 0.00172226 3.3 0.0017221799999999998 3.3 0.0017222799999999999 0 0.0017222 0 0.0017223 3.3 0.00172222 3.3 0.00172232 0 0.0017222399999999999 0 0.00172234 3.3 0.00172226 3.3 0.00172236 0 0.0017222799999999999 0 0.00172238 3.3 0.0017223 3.3 0.0017224 0 0.0017223199999999998 0 0.00172242 3.3 0.00172234 3.3 0.00172244 0 0.0017223599999999998 0 0.0017224599999999999 3.3 0.00172238 3.3 0.00172248 0 0.0017224 0 0.0017225 3.3 0.00172242 3.3 0.00172252 0 0.00172244 0 0.00172254 3.3 0.0017224599999999999 3.3 0.00172256 0 0.00172248 0 0.00172258 3.3 0.0017224999999999999 3.3 0.0017226 0 0.00172252 0 0.00172262 3.3 0.0017225399999999998 3.3 0.00172264 0 0.00172256 0 0.00172266 3.3 0.0017225799999999998 3.3 0.0017226799999999999 0 0.0017226 0 0.0017227 3.3 0.00172262 3.3 0.00172272 0 0.00172264 0 0.00172274 3.3 0.00172266 3.3 0.00172276 0 0.0017226799999999999 0 0.00172278 3.3 0.0017227 3.3 0.0017228 0 0.0017227199999999999 0 0.00172282 3.3 0.00172274 3.3 0.00172284 0 0.0017227599999999998 0 0.0017228599999999999 3.3 0.00172278 3.3 0.00172288 0 0.0017227999999999998 0 0.0017228999999999999 3.3 0.00172282 3.3 0.00172292 0 0.00172284 0 0.00172294 3.3 0.0017228599999999999 3.3 0.00172296 0 0.00172288 0 0.00172298 3.3 0.0017228999999999999 3.3 0.001723 0 0.00172292 0 0.00172302 3.3 0.0017229399999999998 3.3 0.00172304 0 0.00172296 0 0.00172306 3.3 0.0017229799999999998 3.3 0.0017230799999999999 0 0.001723 0 0.0017231 3.3 0.0017230199999999998 3.3 0.0017231199999999999 0 0.00172304 0 0.00172314 3.3 0.00172306 3.3 0.00172316 0 0.0017230799999999999 0 0.00172318 3.3 0.0017231 3.3 0.0017232 0 0.0017231199999999999 0 0.00172322 3.3 0.00172314 3.3 0.00172324 0 0.0017231599999999998 0 0.00172326 3.3 0.00172318 3.3 0.00172328 0 0.0017231999999999998 0 0.0017232999999999999 3.3 0.00172322 3.3 0.00172332 0 0.00172324 0 0.00172334 3.3 0.00172326 3.3 0.00172336 0 0.00172328 0 0.00172338 3.3 0.0017232999999999999 3.3 0.0017234 0 0.00172332 0 0.00172342 3.3 0.0017233399999999999 3.3 0.00172344 0 0.00172336 0 0.00172346 3.3 0.0017233799999999998 3.3 0.0017234799999999999 0 0.0017234 0 0.0017235 3.3 0.0017234199999999998 3.3 0.0017235199999999999 0 0.00172344 0 0.00172354 3.3 0.00172346 3.3 0.00172356 0 0.0017234799999999999 0 0.00172358 3.3 0.0017235 3.3 0.0017236 0 0.0017235199999999999 0 0.00172362 3.3 0.00172354 3.3 0.00172364 0 0.0017235599999999998 0 0.00172366 3.3 0.00172358 3.3 0.00172368 0 0.0017235999999999998 0 0.0017236999999999999 3.3 0.00172362 3.3 0.00172372 0 0.0017236399999999998 0 0.0017237399999999999 3.3 0.00172366 3.3 0.00172376 0 0.00172368 0 0.00172378 3.3 0.0017236999999999999 3.3 0.0017238 0 0.00172372 0 0.00172382 3.3 0.0017237399999999999 3.3 0.00172384 0 0.00172376 0 0.00172386 3.3 0.0017237799999999998 3.3 0.00172388 0 0.0017238 0 0.0017239 3.3 0.0017238199999999998 3.3 0.0017239199999999999 0 0.00172384 0 0.00172394 3.3 0.0017238599999999998 3.3 0.0017239599999999999 0 0.00172388 0 0.00172398 3.3 0.0017239 3.3 0.001724 0 0.0017239199999999999 0 0.00172402 3.3 0.00172394 3.3 0.00172404 0 0.0017239599999999999 0 0.00172406 3.3 0.00172398 3.3 0.00172408 0 0.0017239999999999998 0 0.0017241 3.3 0.00172402 3.3 0.00172412 0 0.0017240399999999998 0 0.0017241399999999999 3.3 0.00172406 3.3 0.00172416 0 0.00172408 0 0.00172418 3.3 0.0017241 3.3 0.0017242 0 0.00172412 0 0.00172422 3.3 0.0017241399999999999 3.3 0.00172424 0 0.00172416 0 0.00172426 3.3 0.0017241799999999999 3.3 0.00172428 0 0.0017242 0 0.0017243 3.3 0.0017242199999999998 3.3 0.0017243199999999999 0 0.00172424 0 0.00172434 3.3 0.0017242599999999998 3.3 0.0017243599999999999 0 0.00172428 0 0.00172438 3.3 0.0017243 3.3 0.0017244 0 0.0017243199999999999 0 0.00172442 3.3 0.00172434 3.3 0.00172444 0 0.0017243599999999999 0 0.00172446 3.3 0.00172438 3.3 0.00172448 0 0.0017243999999999998 0 0.0017245 3.3 0.00172442 3.3 0.00172452 0 0.0017244399999999998 0 0.0017245399999999999 3.3 0.00172446 3.3 0.00172456 0 0.0017244799999999998 0 0.0017245799999999999 3.3 0.0017245 3.3 0.0017246 0 0.00172452 0 0.00172462 3.3 0.0017245399999999999 3.3 0.00172464 0 0.00172456 0 0.00172466 3.3 0.0017245799999999999 3.3 0.00172468 0 0.0017246 0 0.0017247 3.3 0.0017246199999999998 3.3 0.00172472 0 0.00172464 0 0.00172474 3.3 0.0017246599999999998 3.3 0.0017247599999999999 0 0.00172468 0 0.00172478 3.3 0.0017246999999999998 3.3 0.0017247999999999999 0 0.00172472 0 0.00172482 3.3 0.00172474 3.3 0.00172484 0 0.0017247599999999999 0 0.00172486 3.3 0.00172478 3.3 0.00172488 0 0.0017247999999999999 0 0.0017249 3.3 0.00172482 3.3 0.00172492 0 0.0017248399999999998 0 0.00172494 3.3 0.00172486 3.3 0.00172496 0 0.0017248799999999998 0 0.0017249799999999999 3.3 0.0017249 3.3 0.001725 0 0.00172492 0 0.00172502 3.3 0.00172494 3.3 0.00172504 0 0.00172496 0 0.00172506 3.3 0.0017249799999999999 3.3 0.00172508 0 0.001725 0 0.0017251 3.3 0.0017250199999999999 3.3 0.00172512 0 0.00172504 0 0.00172514 3.3 0.0017250599999999998 3.3 0.0017251599999999999 0 0.00172508 0 0.00172518 3.3 0.0017250999999999998 3.3 0.0017251999999999999 0 0.00172512 0 0.00172522 3.3 0.00172514 3.3 0.00172524 0 0.0017251599999999999 0 0.00172526 3.3 0.00172518 3.3 0.00172528 0 0.0017251999999999999 0 0.0017253 3.3 0.00172522 3.3 0.00172532 0 0.0017252399999999998 0 0.00172534 3.3 0.00172526 3.3 0.00172536 0 0.0017252799999999998 0 0.0017253799999999999 3.3 0.0017253 3.3 0.0017254 0 0.0017253199999999998 0 0.0017254199999999999 3.3 0.00172534 3.3 0.00172544 0 0.00172536 0 0.00172546 3.3 0.0017253799999999999 3.3 0.00172548 0 0.0017254 0 0.0017255 3.3 0.0017254199999999999 3.3 0.00172552 0 0.00172544 0 0.00172554 3.3 0.0017254599999999998 3.3 0.00172556 0 0.00172548 0 0.00172558 3.3 0.0017254999999999998 3.3 0.0017255999999999999 0 0.00172552 0 0.00172562 3.3 0.00172554 3.3 0.00172564 0 0.00172556 0 0.00172566 3.3 0.00172558 3.3 0.00172568 0 0.0017255999999999999 0 0.0017257 3.3 0.00172562 3.3 0.00172572 0 0.0017256399999999999 0 0.00172574 3.3 0.00172566 3.3 0.00172576 0 0.0017256799999999998 0 0.00172578 3.3 0.0017257 3.3 0.0017258 0 0.0017257199999999998 0 0.0017258199999999999 3.3 0.00172574 3.3 0.00172584 0 0.00172576 0 0.00172586 3.3 0.00172578 3.3 0.00172588 0 0.0017258 0 0.0017259 3.3 0.0017258199999999999 3.3 0.00172592 0 0.00172584 0 0.00172594 3.3 0.0017258599999999999 3.3 0.00172596 0 0.00172588 0 0.00172598 3.3 0.0017258999999999998 3.3 0.0017259999999999999 0 0.00172592 0 0.00172602 3.3 0.0017259399999999998 3.3 0.0017260399999999999 0 0.00172596 0 0.00172606 3.3 0.00172598 3.3 0.00172608 0 0.0017259999999999999 0 0.0017261 3.3 0.00172602 3.3 0.00172612 0 0.0017260399999999999 0 0.00172614 3.3 0.00172606 3.3 0.00172616 0 0.0017260799999999998 0 0.00172618 3.3 0.0017261 3.3 0.0017262 0 0.0017261199999999998 0 0.0017262199999999999 3.3 0.00172614 3.3 0.00172624 0 0.0017261599999999998 0 0.0017262599999999999 3.3 0.00172618 3.3 0.00172628 0 0.0017262 0 0.0017263 3.3 0.0017262199999999999 3.3 0.00172632 0 0.00172624 0 0.00172634 3.3 0.0017262599999999999 3.3 0.00172636 0 0.00172628 0 0.00172638 3.3 0.0017262999999999998 3.3 0.0017264 0 0.00172632 0 0.00172642 3.3 0.0017263399999999998 3.3 0.0017264399999999999 0 0.00172636 0 0.00172646 3.3 0.00172638 3.3 0.00172648 0 0.0017264 0 0.0017265 3.3 0.00172642 3.3 0.00172652 0 0.0017264399999999999 0 0.00172654 3.3 0.00172646 3.3 0.00172656 0 0.0017264799999999999 0 0.00172658 3.3 0.0017265 3.3 0.0017266 0 0.0017265199999999998 0 0.0017266199999999999 3.3 0.00172654 3.3 0.00172664 0 0.0017265599999999998 0 0.0017266599999999999 3.3 0.00172658 3.3 0.00172668 0 0.0017266 0 0.0017267 3.3 0.0017266199999999999 3.3 0.00172672 0 0.00172664 0 0.00172674 3.3 0.0017266599999999999 3.3 0.00172676 0 0.00172668 0 0.00172678 3.3 0.0017266999999999998 3.3 0.0017268 0 0.00172672 0 0.00172682 3.3 0.0017267399999999998 3.3 0.0017268399999999999 0 0.00172676 0 0.00172686 3.3 0.0017267799999999998 3.3 0.0017268799999999999 0 0.0017268 0 0.0017269 3.3 0.00172682 3.3 0.00172692 0 0.0017268399999999999 0 0.00172694 3.3 0.00172686 3.3 0.00172696 0 0.0017268799999999999 0 0.00172698 3.3 0.0017269 3.3 0.001727 0 0.0017269199999999998 0 0.00172702 3.3 0.00172694 3.3 0.00172704 0 0.0017269599999999998 0 0.0017270599999999999 3.3 0.00172698 3.3 0.00172708 0 0.0017269999999999998 0 0.0017270999999999999 3.3 0.00172702 3.3 0.00172712 0 0.00172704 0 0.00172714 3.3 0.0017270599999999999 3.3 0.00172716 0 0.00172708 0 0.00172718 3.3 0.0017270999999999999 3.3 0.0017272 0 0.00172712 0 0.00172722 3.3 0.0017271399999999998 3.3 0.00172724 0 0.00172716 0 0.00172726 3.3 0.0017271799999999998 3.3 0.0017272799999999999 0 0.0017272 0 0.0017273 3.3 0.00172722 3.3 0.00172732 0 0.00172724 0 0.00172734 3.3 0.00172726 3.3 0.00172736 0 0.0017272799999999999 0 0.00172738 3.3 0.0017273 3.3 0.0017274 0 0.0017273199999999999 0 0.00172742 3.3 0.00172734 3.3 0.00172744 0 0.0017273599999999998 0 0.0017274599999999999 3.3 0.00172738 3.3 0.00172748 0 0.0017273999999999998 0 0.0017274999999999999 3.3 0.00172742 3.3 0.00172752 0 0.00172744 0 0.00172754 3.3 0.0017274599999999999 3.3 0.00172756 0 0.00172748 0 0.00172758 3.3 0.0017274999999999999 3.3 0.0017276 0 0.00172752 0 0.00172762 3.3 0.0017275399999999998 3.3 0.00172764 0 0.00172756 0 0.00172766 3.3 0.0017275799999999998 3.3 0.0017276799999999999 0 0.0017276 0 0.0017277 3.3 0.0017276199999999998 3.3 0.0017277199999999999 0 0.00172764 0 0.00172774 3.3 0.00172766 3.3 0.00172776 0 0.0017276799999999999 0 0.00172778 3.3 0.0017277 3.3 0.0017278 0 0.0017277199999999999 0 0.00172782 3.3 0.00172774 3.3 0.00172784 0 0.0017277599999999998 0 0.00172786 3.3 0.00172778 3.3 0.00172788 0 0.0017277999999999998 0 0.0017278999999999999 3.3 0.00172782 3.3 0.00172792 0 0.0017278399999999998 0 0.0017279399999999999 3.3 0.00172786 3.3 0.00172796 0 0.00172788 0 0.00172798 3.3 0.0017278999999999999 3.3 0.001728 0 0.00172792 0 0.00172802 3.3 0.0017279399999999999 3.3 0.00172804 0 0.00172796 0 0.00172806 3.3 0.0017279799999999998 3.3 0.00172808 0 0.001728 0 0.0017281 3.3 0.0017280199999999998 3.3 0.0017281199999999999 0 0.00172804 0 0.00172814 3.3 0.00172806 3.3 0.00172816 0 0.00172808 0 0.00172818 3.3 0.0017281 3.3 0.0017282 0 0.0017281199999999999 0 0.00172822 3.3 0.00172814 3.3 0.00172824 0 0.0017281599999999999 0 0.00172826 3.3 0.00172818 3.3 0.00172828 0 0.0017281999999999998 0 0.0017282999999999999 3.3 0.00172822 3.3 0.00172832 0 0.0017282399999999998 0 0.0017283399999999999 3.3 0.00172826 3.3 0.00172836 0 0.00172828 0 0.00172838 3.3 0.0017282999999999999 3.3 0.0017284 0 0.00172832 0 0.00172842 3.3 0.0017283399999999999 3.3 0.00172844 0 0.00172836 0 0.00172846 3.3 0.0017283799999999998 3.3 0.00172848 0 0.0017284 0 0.0017285 3.3 0.0017284199999999998 3.3 0.0017285199999999999 0 0.00172844 0 0.00172854 3.3 0.0017284599999999998 3.3 0.0017285599999999999 0 0.00172848 0 0.00172858 3.3 0.0017285 3.3 0.0017286 0 0.0017285199999999999 0 0.00172862 3.3 0.00172854 3.3 0.00172864 0 0.0017285599999999999 0 0.00172866 3.3 0.00172858 3.3 0.00172868 0 0.0017285999999999998 0 0.0017287 3.3 0.00172862 3.3 0.00172872 0 0.0017286399999999998 0 0.0017287399999999999 3.3 0.00172866 3.3 0.00172876 0 0.00172868 0 0.00172878 3.3 0.0017287 3.3 0.0017288 0 0.00172872 0 0.00172882 3.3 0.0017287399999999999 3.3 0.00172884 0 0.00172876 0 0.00172886 3.3 0.0017287799999999999 3.3 0.00172888 0 0.0017288 0 0.0017289 3.3 0.0017288199999999998 3.3 0.00172892 0 0.00172884 0 0.00172894 3.3 0.0017288599999999998 3.3 0.0017289599999999999 0 0.00172888 0 0.00172898 3.3 0.0017289 3.3 0.001729 0 0.00172892 0 0.00172902 3.3 0.00172894 3.3 0.00172904 0 0.0017289599999999999 0 0.00172906 3.3 0.00172898 3.3 0.00172908 0 0.0017289999999999999 0 0.0017291 3.3 0.00172902 3.3 0.00172912 0 0.0017290399999999998 0 0.0017291399999999999 3.3 0.00172906 3.3 0.00172916 0 0.0017290799999999998 0 0.0017291799999999999 3.3 0.0017291 3.3 0.0017292 0 0.00172912 0 0.00172922 3.3 0.0017291399999999999 3.3 0.00172924 0 0.00172916 0 0.00172926 3.3 0.0017291799999999999 3.3 0.00172928 0 0.0017292 0 0.0017293 3.3 0.0017292199999999998 3.3 0.00172932 0 0.00172924 0 0.00172934 3.3 0.0017292599999999998 3.3 0.0017293599999999999 0 0.00172928 0 0.00172938 3.3 0.0017292999999999998 3.3 0.0017293999999999999 0 0.00172932 0 0.00172942 3.3 0.00172934 3.3 0.00172944 0 0.0017293599999999999 0 0.00172946 3.3 0.00172938 3.3 0.00172948 0 0.0017293999999999999 0 0.0017295 3.3 0.00172942 3.3 0.00172952 0 0.0017294399999999998 0 0.00172954 3.3 0.00172946 3.3 0.00172956 0 0.0017294799999999998 0 0.0017295799999999999 3.3 0.0017295 3.3 0.0017296 0 0.00172952 0 0.00172962 3.3 0.00172954 3.3 0.00172964 0 0.00172956 0 0.00172966 3.3 0.0017295799999999999 3.3 0.00172968 0 0.0017296 0 0.0017297 3.3 0.0017296199999999999 3.3 0.00172972 0 0.00172964 0 0.00172974 3.3 0.0017296599999999998 3.3 0.0017297599999999999 0 0.00172968 0 0.00172978 3.3 0.0017296999999999998 3.3 0.0017297999999999999 0 0.00172972 0 0.00172982 3.3 0.00172974 3.3 0.00172984 0 0.0017297599999999999 0 0.00172986 3.3 0.00172978 3.3 0.00172988 0 0.0017297999999999999 0 0.0017299 3.3 0.00172982 3.3 0.00172992 0 0.0017298399999999998 0 0.00172994 3.3 0.00172986 3.3 0.00172996 0 0.0017298799999999998 0 0.0017299799999999999 3.3 0.0017299 3.3 0.00173 0 0.0017299199999999998 0 0.0017300199999999999 3.3 0.00172994 3.3 0.00173004 0 0.00172996 0 0.00173006 3.3 0.0017299799999999999 3.3 0.00173008 0 0.00173 0 0.0017301 3.3 0.0017300199999999999 3.3 0.00173012 0 0.00173004 0 0.00173014 3.3 0.0017300599999999998 3.3 0.00173016 0 0.00173008 0 0.00173018 3.3 0.0017300999999999998 3.3 0.0017301999999999999 0 0.00173012 0 0.00173022 3.3 0.0017301399999999998 3.3 0.0017302399999999999 0 0.00173016 0 0.00173026 3.3 0.00173018 3.3 0.00173028 0 0.0017301999999999999 0 0.0017303 3.3 0.00173022 3.3 0.00173032 0 0.0017302399999999999 0 0.00173034 3.3 0.00173026 3.3 0.00173036 0 0.0017302799999999998 0 0.00173038 3.3 0.0017303 3.3 0.0017304 0 0.0017303199999999998 0 0.0017304199999999999 3.3 0.00173034 3.3 0.00173044 0 0.00173036 0 0.00173046 3.3 0.00173038 3.3 0.00173048 0 0.0017304 0 0.0017305 3.3 0.0017304199999999999 3.3 0.00173052 0 0.00173044 0 0.00173054 3.3 0.0017304599999999999 3.3 0.00173056 0 0.00173048 0 0.00173058 3.3 0.0017304999999999998 3.3 0.0017305999999999999 0 0.00173052 0 0.00173062 3.3 0.0017305399999999998 3.3 0.0017306399999999999 0 0.00173056 0 0.00173066 3.3 0.00173058 3.3 0.00173068 0 0.0017305999999999999 0 0.0017307 3.3 0.00173062 3.3 0.00173072 0 0.0017306399999999999 0 0.00173074 3.3 0.00173066 3.3 0.00173076 0 0.0017306799999999998 0 0.00173078 3.3 0.0017307 3.3 0.0017308 0 0.0017307199999999998 0 0.0017308199999999999 3.3 0.00173074 3.3 0.00173084 0 0.0017307599999999998 0 0.0017308599999999999 3.3 0.00173078 3.3 0.00173088 0 0.0017308 0 0.0017309 3.3 0.0017308199999999999 3.3 0.00173092 0 0.00173084 0 0.00173094 3.3 0.0017308599999999999 3.3 0.00173096 0 0.00173088 0 0.00173098 3.3 0.0017308999999999998 3.3 0.001731 0 0.00173092 0 0.00173102 3.3 0.0017309399999999998 3.3 0.0017310399999999999 0 0.00173096 0 0.00173106 3.3 0.0017309799999999998 3.3 0.0017310799999999999 0 0.001731 0 0.0017311 3.3 0.00173102 3.3 0.00173112 0 0.0017310399999999999 0 0.00173114 3.3 0.00173106 3.3 0.00173116 0 0.0017310799999999999 0 0.00173118 3.3 0.0017311 3.3 0.0017312 0 0.0017311199999999998 0 0.00173122 3.3 0.00173114 3.3 0.00173124 0 0.0017311599999999998 0 0.0017312599999999999 3.3 0.00173118 3.3 0.00173128 0 0.0017312 0 0.0017313 3.3 0.00173122 3.3 0.00173132 0 0.00173124 0 0.00173134 3.3 0.0017312599999999999 3.3 0.00173136 0 0.00173128 0 0.00173138 3.3 0.0017312999999999999 3.3 0.0017314 0 0.00173132 0 0.00173142 3.3 0.0017313399999999998 3.3 0.0017314399999999999 0 0.00173136 0 0.00173146 3.3 0.0017313799999999998 3.3 0.0017314799999999999 0 0.0017314 0 0.0017315 3.3 0.00173142 3.3 0.00173152 0 0.0017314399999999999 0 0.00173154 3.3 0.00173146 3.3 0.00173156 0 0.0017314799999999999 0 0.00173158 3.3 0.0017315 3.3 0.0017316 0 0.0017315199999999998 0 0.00173162 3.3 0.00173154 3.3 0.00173164 0 0.0017315599999999998 0 0.0017316599999999999 3.3 0.00173158 3.3 0.00173168 0 0.0017315999999999998 0 0.0017316999999999999 3.3 0.00173162 3.3 0.00173172 0 0.00173164 0 0.00173174 3.3 0.0017316599999999999 3.3 0.00173176 0 0.00173168 0 0.00173178 3.3 0.0017316999999999999 3.3 0.0017318 0 0.00173172 0 0.00173182 3.3 0.0017317399999999998 3.3 0.00173184 0 0.00173176 0 0.00173186 3.3 0.0017317799999999998 3.3 0.0017318799999999999 0 0.0017318 0 0.0017319 3.3 0.0017318199999999998 3.3 0.0017319199999999999 0 0.00173184 0 0.00173194 3.3 0.00173186 3.3 0.00173196 0 0.0017318799999999999 0 0.00173198 3.3 0.0017319 3.3 0.001732 0 0.0017319199999999999 0 0.00173202 3.3 0.00173194 3.3 0.00173204 0 0.0017319599999999998 0 0.00173206 3.3 0.00173198 3.3 0.00173208 0 0.0017319999999999998 0 0.0017320999999999999 3.3 0.00173202 3.3 0.00173212 0 0.00173204 0 0.00173214 3.3 0.00173206 3.3 0.00173216 0 0.00173208 0 0.00173218 3.3 0.0017320999999999999 3.3 0.0017322 0 0.00173212 0 0.00173222 3.3 0.0017321399999999999 3.3 0.00173224 0 0.00173216 0 0.00173226 3.3 0.0017321799999999998 3.3 0.0017322799999999999 0 0.0017322 0 0.0017323 3.3 0.0017322199999999998 3.3 0.0017323199999999999 0 0.00173224 0 0.00173234 3.3 0.00173226 3.3 0.00173236 0 0.0017322799999999999 0 0.00173238 3.3 0.0017323 3.3 0.0017324 0 0.0017323199999999999 0 0.00173242 3.3 0.00173234 3.3 0.00173244 0 0.0017323599999999998 0 0.00173246 3.3 0.00173238 3.3 0.00173248 0 0.0017323999999999998 0 0.0017324999999999999 3.3 0.00173242 3.3 0.00173252 0 0.0017324399999999998 0 0.0017325399999999999 3.3 0.00173246 3.3 0.00173256 0 0.00173248 0 0.00173258 3.3 0.0017324999999999999 3.3 0.0017326 0 0.00173252 0 0.00173262 3.3 0.0017325399999999999 3.3 0.00173264 0 0.00173256 0 0.00173266 3.3 0.0017325799999999998 3.3 0.00173268 0 0.0017326 0 0.0017327 3.3 0.0017326199999999998 3.3 0.0017327199999999999 0 0.00173264 0 0.00173274 3.3 0.00173266 3.3 0.00173276 0 0.00173268 0 0.00173278 3.3 0.0017327 3.3 0.0017328 0 0.0017327199999999999 0 0.00173282 3.3 0.00173274 3.3 0.00173284 0 0.0017327599999999999 0 0.00173286 3.3 0.00173278 3.3 0.00173288 0 0.0017327999999999998 0 0.0017329 3.3 0.00173282 3.3 0.00173292 0 0.0017328399999999998 0 0.0017329399999999999 3.3 0.00173286 3.3 0.00173296 0 0.00173288 0 0.00173298 3.3 0.0017329 3.3 0.001733 0 0.00173292 0 0.00173302 3.3 0.0017329399999999999 3.3 0.00173304 0 0.00173296 0 0.00173306 3.3 0.0017329799999999999 3.3 0.00173308 0 0.001733 0 0.0017331 3.3 0.0017330199999999998 3.3 0.0017331199999999999 0 0.00173304 0 0.00173314 3.3 0.0017330599999999998 3.3 0.0017331599999999999 0 0.00173308 0 0.00173318 3.3 0.0017331 3.3 0.0017332 0 0.0017331199999999999 0 0.00173322 3.3 0.00173314 3.3 0.00173324 0 0.0017331599999999999 0 0.00173326 3.3 0.00173318 3.3 0.00173328 0 0.0017331999999999998 0 0.0017333 3.3 0.00173322 3.3 0.00173332 0 0.0017332399999999998 0 0.0017333399999999999 3.3 0.00173326 3.3 0.00173336 0 0.0017332799999999998 0 0.0017333799999999999 3.3 0.0017333 3.3 0.0017334 0 0.00173332 0 0.00173342 3.3 0.0017333399999999999 3.3 0.00173344 0 0.00173336 0 0.00173346 3.3 0.0017333799999999999 3.3 0.00173348 0 0.0017334 0 0.0017335 3.3 0.0017334199999999998 3.3 0.00173352 0 0.00173344 0 0.00173354 3.3 0.0017334599999999998 3.3 0.0017335599999999999 0 0.00173348 0 0.00173358 3.3 0.0017335 3.3 0.0017336 0 0.00173352 0 0.00173362 3.3 0.00173354 3.3 0.00173364 0 0.0017335599999999999 0 0.00173366 3.3 0.00173358 3.3 0.00173368 0 0.0017335999999999999 0 0.0017337 3.3 0.00173362 3.3 0.00173372 0 0.0017336399999999998 0 0.0017337399999999999 3.3 0.00173366 3.3 0.00173376 0 0.0017336799999999998 0 0.0017337799999999999 3.3 0.0017337 3.3 0.0017338 0 0.00173372 0 0.00173382 3.3 0.0017337399999999999 3.3 0.00173384 0 0.00173376 0 0.00173386 3.3 0.0017337799999999999 3.3 0.00173388 0 0.0017338 0 0.0017339 3.3 0.0017338199999999998 3.3 0.00173392 0 0.00173384 0 0.00173394 3.3 0.0017338599999999998 3.3 0.0017339599999999999 0 0.00173388 0 0.00173398 3.3 0.0017338999999999998 3.3 0.0017339999999999999 0 0.00173392 0 0.00173402 3.3 0.00173394 3.3 0.00173404 0 0.0017339599999999999 0 0.00173406 3.3 0.00173398 3.3 0.00173408 0 0.0017339999999999999 0 0.0017341 3.3 0.00173402 3.3 0.00173412 0 0.0017340399999999998 0 0.00173414 3.3 0.00173406 3.3 0.00173416 0 0.0017340799999999998 0 0.0017341799999999999 3.3 0.0017341 3.3 0.0017342 0 0.0017341199999999998 0 0.0017342199999999999 3.3 0.00173414 3.3 0.00173424 0 0.00173416 0 0.00173426 3.3 0.0017341799999999999 3.3 0.00173428 0 0.0017342 0 0.0017343 3.3 0.0017342199999999999 3.3 0.00173432 0 0.00173424 0 0.00173434 3.3 0.0017342599999999998 3.3 0.00173436 0 0.00173428 0 0.00173438 3.3 0.0017342999999999998 3.3 0.0017343999999999999 0 0.00173432 0 0.00173442 3.3 0.00173434 3.3 0.00173444 0 0.00173436 0 0.00173446 3.3 0.00173438 3.3 0.00173448 0 0.0017343999999999999 0 0.0017345 3.3 0.00173442 3.3 0.00173452 0 0.0017344399999999999 0 0.00173454 3.3 0.00173446 3.3 0.00173456 0 0.0017344799999999998 0 0.0017345799999999999 3.3 0.0017345 3.3 0.0017346 0 0.0017345199999999998 0 0.0017346199999999999 3.3 0.00173454 3.3 0.00173464 0 0.00173456 0 0.00173466 3.3 0.0017345799999999999 3.3 0.00173468 0 0.0017346 0 0.0017347 3.3 0.0017346199999999999 3.3 0.00173472 0 0.00173464 0 0.00173474 3.3 0.0017346599999999998 3.3 0.00173476 0 0.00173468 0 0.00173478 3.3 0.0017346999999999998 3.3 0.0017347999999999999 0 0.00173472 0 0.00173482 3.3 0.0017347399999999998 3.3 0.0017348399999999999 0 0.00173476 0 0.00173486 3.3 0.00173478 3.3 0.00173488 0 0.0017347999999999999 0 0.0017349 3.3 0.00173482 3.3 0.00173492 0 0.0017348399999999999 0 0.00173494 3.3 0.00173486 3.3 0.00173496 0 0.0017348799999999998 0 0.00173498 3.3 0.0017349 3.3 0.001735 0 0.0017349199999999998 0 0.0017350199999999999 3.3 0.00173494 3.3 0.00173504 0 0.0017349599999999998 0 0.0017350599999999999 3.3 0.00173498 3.3 0.00173508 0 0.001735 0 0.0017351 3.3 0.0017350199999999999 3.3 0.00173512 0 0.00173504 0 0.00173514 3.3 0.0017350599999999999 3.3 0.00173516 0 0.00173508 0 0.00173518 3.3 0.0017350999999999998 3.3 0.0017352 0 0.00173512 0 0.00173522 3.3 0.0017351399999999998 3.3 0.0017352399999999999 0 0.00173516 0 0.00173526 3.3 0.00173518 3.3 0.00173528 0 0.0017352 0 0.0017353 3.3 0.00173522 3.3 0.00173532 0 0.0017352399999999999 0 0.00173534 3.3 0.00173526 3.3 0.00173536 0 0.0017352799999999999 0 0.00173538 3.3 0.0017353 3.3 0.0017354 0 0.0017353199999999998 0 0.0017354199999999999 3.3 0.00173534 3.3 0.00173544 0 0.0017353599999999998 0 0.0017354599999999999 3.3 0.00173538 3.3 0.00173548 0 0.0017354 0 0.0017355 3.3 0.0017354199999999999 3.3 0.00173552 0 0.00173544 0 0.00173554 3.3 0.0017354599999999999 3.3 0.00173556 0 0.00173548 0 0.00173558 3.3 0.0017354999999999998 3.3 0.0017356 0 0.00173552 0 0.00173562 3.3 0.0017355399999999998 3.3 0.0017356399999999999 0 0.00173556 0 0.00173566 3.3 0.0017355799999999998 3.3 0.0017356799999999999 0 0.0017356 0 0.0017357 3.3 0.00173562 3.3 0.00173572 0 0.0017356399999999999 0 0.00173574 3.3 0.00173566 3.3 0.00173576 0 0.0017356799999999999 0 0.00173578 3.3 0.0017357 3.3 0.0017358 0 0.0017357199999999998 0 0.00173582 3.3 0.00173574 3.3 0.00173584 0 0.0017357599999999998 0 0.0017358599999999999 3.3 0.00173578 3.3 0.00173588 0 0.0017358 0 0.0017359 3.3 0.00173582 3.3 0.00173592 0 0.00173584 0 0.00173594 3.3 0.0017358599999999999 3.3 0.00173596 0 0.00173588 0 0.00173598 3.3 0.0017358999999999999 3.3 0.001736 0 0.00173592 0 0.00173602 3.3 0.0017359399999999998 3.3 0.00173604 0 0.00173596 0 0.00173606 3.3 0.0017359799999999998 3.3 0.0017360799999999999 0 0.001736 0 0.0017361 3.3 0.00173602 3.3 0.00173612 0 0.00173604 0 0.00173614 3.3 0.00173606 3.3 0.00173616 0 0.0017360799999999999 0 0.00173618 3.3 0.0017361 3.3 0.0017362 0 0.0017361199999999999 0 0.00173622 3.3 0.00173614 3.3 0.00173624 0 0.0017361599999999998 0 0.0017362599999999999 3.3 0.00173618 3.3 0.00173628 0 0.0017361999999999998 0 0.0017362999999999999 3.3 0.00173622 3.3 0.00173632 0 0.00173624 0 0.00173634 3.3 0.0017362599999999999 3.3 0.00173636 0 0.00173628 0 0.00173638 3.3 0.0017362999999999999 3.3 0.0017364 0 0.00173632 0 0.00173642 3.3 0.0017363399999999998 3.3 0.00173644 0 0.00173636 0 0.00173646 3.3 0.0017363799999999998 3.3 0.0017364799999999999 0 0.0017364 0 0.0017365 3.3 0.0017364199999999998 3.3 0.0017365199999999999 0 0.00173644 0 0.00173654 3.3 0.00173646 3.3 0.00173656 0 0.0017364799999999999 0 0.00173658 3.3 0.0017365 3.3 0.0017366 0 0.0017365199999999999 0 0.00173662 3.3 0.00173654 3.3 0.00173664 0 0.0017365599999999998 0 0.00173666 3.3 0.00173658 3.3 0.00173668 0 0.0017365999999999998 0 0.0017366999999999999 3.3 0.00173662 3.3 0.00173672 0 0.00173664 0 0.00173674 3.3 0.00173666 3.3 0.00173676 0 0.00173668 0 0.00173678 3.3 0.0017366999999999999 3.3 0.0017368 0 0.00173672 0 0.00173682 3.3 0.0017367399999999999 3.3 0.00173684 0 0.00173676 0 0.00173686 3.3 0.0017367799999999998 3.3 0.0017368799999999999 0 0.0017368 0 0.0017369 3.3 0.0017368199999999998 3.3 0.0017369199999999999 0 0.00173684 0 0.00173694 3.3 0.00173686 3.3 0.00173696 0 0.0017368799999999999 0 0.00173698 3.3 0.0017369 3.3 0.001737 0 0.0017369199999999999 0 0.00173702 3.3 0.00173694 3.3 0.00173704 0 0.0017369599999999998 0 0.00173706 3.3 0.00173698 3.3 0.00173708 0 0.0017369999999999998 0 0.0017370999999999999 3.3 0.00173702 3.3 0.00173712 0 0.0017370399999999998 0 0.0017371399999999999 3.3 0.00173706 3.3 0.00173716 0 0.00173708 0 0.00173718 3.3 0.0017370999999999999 3.3 0.0017372 0 0.00173712 0 0.00173722 3.3 0.0017371399999999999 3.3 0.00173724 0 0.00173716 0 0.00173726 3.3 0.0017371799999999998 3.3 0.00173728 0 0.0017372 0 0.0017373 3.3 0.0017372199999999998 3.3 0.0017373199999999999 0 0.00173724 0 0.00173734 3.3 0.0017372599999999998 3.3 0.0017373599999999999 0 0.00173728 0 0.00173738 3.3 0.0017373 3.3 0.0017374 0 0.0017373199999999999 0 0.00173742 3.3 0.00173734 3.3 0.00173744 0 0.0017373599999999999 0 0.00173746 3.3 0.00173738 3.3 0.00173748 0 0.0017373999999999998 0 0.0017375 3.3 0.00173742 3.3 0.00173752 0 0.0017374399999999998 0 0.0017375399999999999 3.3 0.00173746 3.3 0.00173756 0 0.00173748 0 0.00173758 3.3 0.0017375 3.3 0.0017376 0 0.00173752 0 0.00173762 3.3 0.0017375399999999999 3.3 0.00173764 0 0.00173756 0 0.00173766 3.3 0.0017375799999999999 3.3 0.00173768 0 0.0017376 0 0.0017377 3.3 0.0017376199999999998 3.3 0.0017377199999999999 0 0.00173764 0 0.00173774 3.3 0.0017376599999999998 3.3 0.0017377599999999999 0 0.00173768 0 0.00173778 3.3 0.0017377 3.3 0.0017378 0 0.0017377199999999999 0 0.00173782 3.3 0.00173774 3.3 0.00173784 0 0.0017377599999999999 0 0.00173786 3.3 0.00173778 3.3 0.00173788 0 0.0017377999999999998 0 0.0017379 3.3 0.00173782 3.3 0.00173792 0 0.0017378399999999998 0 0.0017379399999999999 3.3 0.00173786 3.3 0.00173796 0 0.0017378799999999998 0 0.0017379799999999999 3.3 0.0017379 3.3 0.001738 0 0.00173792 0 0.00173802 3.3 0.0017379399999999999 3.3 0.00173804 0 0.00173796 0 0.00173806 3.3 0.0017379799999999999 3.3 0.00173808 0 0.001738 0 0.0017381 3.3 0.0017380199999999998 3.3 0.00173812 0 0.00173804 0 0.00173814 3.3 0.0017380599999999998 3.3 0.0017381599999999999 0 0.00173808 0 0.00173818 3.3 0.0017380999999999998 3.3 0.0017381999999999999 0 0.00173812 0 0.00173822 3.3 0.00173814 3.3 0.00173824 0 0.0017381599999999999 0 0.00173826 3.3 0.00173818 3.3 0.00173828 0 0.0017381999999999999 0 0.0017383 3.3 0.00173822 3.3 0.00173832 0 0.0017382399999999998 0 0.00173834 3.3 0.00173826 3.3 0.00173836 0 0.0017382799999999998 0 0.0017383799999999999 3.3 0.0017383 3.3 0.0017384 0 0.00173832 0 0.00173842 3.3 0.00173834 3.3 0.00173844 0 0.00173836 0 0.00173846 3.3 0.0017383799999999999 3.3 0.00173848 0 0.0017384 0 0.0017385 3.3 0.0017384199999999999 3.3 0.00173852 0 0.00173844 0 0.00173854 3.3 0.0017384599999999998 3.3 0.0017385599999999999 0 0.00173848 0 0.00173858 3.3 0.0017384999999999998 3.3 0.0017385999999999999 0 0.00173852 0 0.00173862 3.3 0.00173854 3.3 0.00173864 0 0.0017385599999999999 0 0.00173866 3.3 0.00173858 3.3 0.00173868 0 0.0017385999999999999 0 0.0017387 3.3 0.00173862 3.3 0.00173872 0 0.0017386399999999998 0 0.00173874 3.3 0.00173866 3.3 0.00173876 0 0.0017386799999999998 0 0.0017387799999999999 3.3 0.0017387 3.3 0.0017388 0 0.0017387199999999998 0 0.0017388199999999999 3.3 0.00173874 3.3 0.00173884 0 0.00173876 0 0.00173886 3.3 0.0017387799999999999 3.3 0.00173888 0 0.0017388 0 0.0017389 3.3 0.0017388199999999999 3.3 0.00173892 0 0.00173884 0 0.00173894 3.3 0.0017388599999999998 3.3 0.00173896 0 0.00173888 0 0.00173898 3.3 0.0017388999999999998 3.3 0.0017389999999999999 0 0.00173892 0 0.00173902 3.3 0.0017389399999999998 3.3 0.0017390399999999999 0 0.00173896 0 0.00173906 3.3 0.00173898 3.3 0.00173908 0 0.0017389999999999999 0 0.0017391 3.3 0.00173902 3.3 0.00173912 0 0.0017390399999999999 0 0.00173914 3.3 0.00173906 3.3 0.00173916 0 0.0017390799999999998 0 0.00173918 3.3 0.0017391 3.3 0.0017392 0 0.0017391199999999998 0 0.0017392199999999999 3.3 0.00173914 3.3 0.00173924 0 0.00173916 0 0.00173926 3.3 0.00173918 3.3 0.00173928 0 0.0017392 0 0.0017393 3.3 0.0017392199999999999 3.3 0.00173932 0 0.00173924 0 0.00173934 3.3 0.0017392599999999999 3.3 0.00173936 0 0.00173928 0 0.00173938 3.3 0.0017392999999999998 3.3 0.0017393999999999999 0 0.00173932 0 0.00173942 3.3 0.0017393399999999998 3.3 0.0017394399999999999 0 0.00173936 0 0.00173946 3.3 0.00173938 3.3 0.00173948 0 0.0017393999999999999 0 0.0017395 3.3 0.00173942 3.3 0.00173952 0 0.0017394399999999999 0 0.00173954 3.3 0.00173946 3.3 0.00173956 0 0.0017394799999999998 0 0.00173958 3.3 0.0017395 3.3 0.0017396 0 0.0017395199999999998 0 0.0017396199999999999 3.3 0.00173954 3.3 0.00173964 0 0.0017395599999999998 0 0.0017396599999999999 3.3 0.00173958 3.3 0.00173968 0 0.0017396 0 0.0017397 3.3 0.0017396199999999999 3.3 0.00173972 0 0.00173964 0 0.00173974 3.3 0.0017396599999999999 3.3 0.00173976 0 0.00173968 0 0.00173978 3.3 0.0017396999999999998 3.3 0.0017398 0 0.00173972 0 0.00173982 3.3 0.0017397399999999998 3.3 0.0017398399999999999 0 0.00173976 0 0.00173986 3.3 0.00173978 3.3 0.00173988 0 0.0017398 0 0.0017399 3.3 0.00173982 3.3 0.00173992 0 0.0017398399999999999 0 0.00173994 3.3 0.00173986 3.3 0.00173996 0 0.0017398799999999999 0 0.00173998 3.3 0.0017399 3.3 0.00174 0 0.0017399199999999998 0 0.0017400199999999999 3.3 0.00173994 3.3 0.00174004 0 0.0017399599999999998 0 0.0017400599999999999 3.3 0.00173998 3.3 0.00174008 0 0.00174 0 0.0017401 3.3 0.0017400199999999999 3.3 0.00174012 0 0.00174004 0 0.00174014 3.3 0.0017400599999999999 3.3 0.00174016 0 0.00174008 0 0.00174018 3.3 0.0017400999999999999 3.3 0.0017402 0 0.00174012 0 0.00174022 3.3 0.0017401399999999998 3.3 0.0017402399999999999 0 0.00174016 0 0.00174026 3.3 0.0017401799999999998 3.3 0.0017402799999999999 0 0.0017402 0 0.0017403 3.3 0.00174022 3.3 0.00174032 0 0.0017402399999999999 0 0.00174034 3.3 0.00174026 3.3 0.00174036 0 0.0017402799999999999 0 0.00174038 3.3 0.0017403 3.3 0.0017404 0 0.0017403199999999998 0 0.00174042 3.3 0.00174034 3.3 0.00174044 0 0.0017403599999999998 0 0.0017404599999999999 3.3 0.00174038 3.3 0.00174048 0 0.0017403999999999998 0 0.0017404999999999999 3.3 0.00174042 3.3 0.00174052 0 0.00174044 0 0.00174054 3.3 0.0017404599999999999 3.3 0.00174056 0 0.00174048 0 0.00174058 3.3 0.0017404999999999999 3.3 0.0017406 0 0.00174052 0 0.00174062 3.3 0.0017405399999999998 3.3 0.00174064 0 0.00174056 0 0.00174066 3.3 0.0017405799999999998 3.3 0.0017406799999999999 0 0.0017406 0 0.0017407 3.3 0.00174062 3.3 0.00174072 0 0.00174064 0 0.00174074 3.3 0.00174066 3.3 0.00174076 0 0.0017406799999999999 0 0.00174078 3.3 0.0017407 3.3 0.0017408 0 0.0017407199999999999 0 0.00174082 3.3 0.00174074 3.3 0.00174084 0 0.0017407599999999998 0 0.0017408599999999999 3.3 0.00174078 3.3 0.00174088 0 0.0017407999999999998 0 0.0017408999999999999 3.3 0.00174082 3.3 0.00174092 0 0.00174084 0 0.00174094 3.3 0.0017408599999999999 3.3 0.00174096 0 0.00174088 0 0.00174098 3.3 0.0017408999999999999 3.3 0.001741 0 0.00174092 0 0.00174102 3.3 0.0017409399999999998 3.3 0.00174104 0 0.00174096 0 0.00174106 3.3 0.0017409799999999998 3.3 0.0017410799999999999 0 0.001741 0 0.0017411 3.3 0.0017410199999999998 3.3 0.0017411199999999999 0 0.00174104 0 0.00174114 3.3 0.00174106 3.3 0.00174116 0 0.0017410799999999999 0 0.00174118 3.3 0.0017411 3.3 0.0017412 0 0.0017411199999999999 0 0.00174122 3.3 0.00174114 3.3 0.00174124 0 0.0017411599999999998 0 0.00174126 3.3 0.00174118 3.3 0.00174128 0 0.0017411999999999998 0 0.0017412999999999999 3.3 0.00174122 3.3 0.00174132 0 0.0017412399999999998 0 0.0017413399999999999 3.3 0.00174126 3.3 0.00174136 0 0.00174128 0 0.00174138 3.3 0.0017412999999999999 3.3 0.0017414 0 0.00174132 0 0.00174142 3.3 0.0017413399999999999 3.3 0.00174144 0 0.00174136 0 0.00174146 3.3 0.0017413799999999998 3.3 0.00174148 0 0.0017414 0 0.0017415 3.3 0.0017414199999999998 3.3 0.0017415199999999999 0 0.00174144 0 0.00174154 3.3 0.00174146 3.3 0.00174156 0 0.00174148 0 0.00174158 3.3 0.0017415 3.3 0.0017416 0 0.0017415199999999999 0 0.00174162 3.3 0.00174154 3.3 0.00174164 0 0.0017415599999999999 0 0.00174166 3.3 0.00174158 3.3 0.00174168 0 0.0017415999999999998 0 0.0017416999999999999 3.3 0.00174162 3.3 0.00174172 0 0.0017416399999999998 0 0.0017417399999999999 3.3 0.00174166 3.3 0.00174176 0 0.00174168 0 0.00174178 3.3 0.0017416999999999999 3.3 0.0017418 0 0.00174172 0 0.00174182 3.3 0.0017417399999999999 3.3 0.00174184 0 0.00174176 0 0.00174186 3.3 0.0017417799999999998 3.3 0.00174188 0 0.0017418 0 0.0017419 3.3 0.0017418199999999998 3.3 0.0017419199999999999 0 0.00174184 0 0.00174194 3.3 0.0017418599999999998 3.3 0.0017419599999999999 0 0.00174188 0 0.00174198 3.3 0.0017419 3.3 0.001742 0 0.0017419199999999999 0 0.00174202 3.3 0.00174194 3.3 0.00174204 0 0.0017419599999999999 0 0.00174206 3.3 0.00174198 3.3 0.00174208 0 0.0017419999999999998 0 0.0017421 3.3 0.00174202 3.3 0.00174212 0 0.0017420399999999998 0 0.0017421399999999999 3.3 0.00174206 3.3 0.00174216 0 0.0017420799999999998 0 0.0017421799999999999 3.3 0.0017421 3.3 0.0017422 0 0.00174212 0 0.00174222 3.3 0.0017421399999999999 3.3 0.00174224 0 0.00174216 0 0.00174226 3.3 0.0017421799999999999 3.3 0.00174228 0 0.0017422 0 0.0017423 3.3 0.0017422199999999998 3.3 0.00174232 0 0.00174224 0 0.00174234 3.3 0.0017422599999999998 3.3 0.0017423599999999999 0 0.00174228 0 0.00174238 3.3 0.0017423 3.3 0.0017424 0 0.00174232 0 0.00174242 3.3 0.00174234 3.3 0.00174244 0 0.0017423599999999999 0 0.00174246 3.3 0.00174238 3.3 0.00174248 0 0.0017423999999999999 0 0.0017425 3.3 0.00174242 3.3 0.00174252 0 0.0017424399999999998 0 0.0017425399999999999 3.3 0.00174246 3.3 0.00174256 0 0.0017424799999999998 0 0.0017425799999999999 3.3 0.0017425 3.3 0.0017426 0 0.00174252 0 0.00174262 3.3 0.0017425399999999999 3.3 0.00174264 0 0.00174256 0 0.00174266 3.3 0.0017425799999999999 3.3 0.00174268 0 0.0017426 0 0.0017427 3.3 0.0017426199999999998 3.3 0.00174272 0 0.00174264 0 0.00174274 3.3 0.0017426599999999998 3.3 0.0017427599999999999 0 0.00174268 0 0.00174278 3.3 0.0017426999999999998 3.3 0.0017427999999999999 0 0.00174272 0 0.00174282 3.3 0.00174274 3.3 0.00174284 0 0.0017427599999999999 0 0.00174286 3.3 0.00174278 3.3 0.00174288 0 0.0017427999999999999 0 0.0017429 3.3 0.00174282 3.3 0.00174292 0 0.0017428399999999998 0 0.00174294 3.3 0.00174286 3.3 0.00174296 0 0.0017428799999999998 0 0.0017429799999999999 3.3 0.0017429 3.3 0.001743 0 0.00174292 0 0.00174302 3.3 0.00174294 3.3 0.00174304 0 0.00174296 0 0.00174306 3.3 0.0017429799999999999 3.3 0.00174308 0 0.001743 0 0.0017431 3.3 0.0017430199999999999 3.3 0.00174312 0 0.00174304 0 0.00174314 3.3 0.0017430599999999998 3.3 0.00174316 0 0.00174308 0 0.00174318 3.3 0.0017430999999999998 3.3 0.0017431999999999999 0 0.00174312 0 0.00174322 3.3 0.00174314 3.3 0.00174324 0 0.00174316 0 0.00174326 3.3 0.00174318 3.3 0.00174328 0 0.0017431999999999999 0 0.0017433 3.3 0.00174322 3.3 0.00174332 0 0.0017432399999999999 0 0.00174334 3.3 0.00174326 3.3 0.00174336 0 0.0017432799999999998 0 0.0017433799999999999 3.3 0.0017433 3.3 0.0017434 0 0.0017433199999999998 0 0.0017434199999999999 3.3 0.00174334 3.3 0.00174344 0 0.00174336 0 0.00174346 3.3 0.0017433799999999999 3.3 0.00174348 0 0.0017434 0 0.0017435 3.3 0.0017434199999999999 3.3 0.00174352 0 0.00174344 0 0.00174354 3.3 0.0017434599999999998 3.3 0.00174356 0 0.00174348 0 0.00174358 3.3 0.0017434999999999998 3.3 0.0017435999999999999 0 0.00174352 0 0.00174362 3.3 0.0017435399999999998 3.3 0.0017436399999999999 0 0.00174356 0 0.00174366 3.3 0.00174358 3.3 0.00174368 0 0.0017435999999999999 0 0.0017437 3.3 0.00174362 3.3 0.00174372 0 0.0017436399999999999 0 0.00174374 3.3 0.00174366 3.3 0.00174376 0 0.0017436799999999998 0 0.00174378 3.3 0.0017437 3.3 0.0017438 0 0.0017437199999999998 0 0.0017438199999999999 3.3 0.00174374 3.3 0.00174384 0 0.00174376 0 0.00174386 3.3 0.00174378 3.3 0.00174388 0 0.0017438 0 0.0017439 3.3 0.0017438199999999999 3.3 0.00174392 0 0.00174384 0 0.00174394 3.3 0.0017438599999999999 3.3 0.00174396 0 0.00174388 0 0.00174398 3.3 0.0017438999999999998 3.3 0.0017439999999999999 0 0.00174392 0 0.00174402 3.3 0.0017439399999999998 3.3 0.0017440399999999999 0 0.00174396 0 0.00174406 3.3 0.00174398 3.3 0.00174408 0 0.0017439999999999999 0 0.0017441 3.3 0.00174402 3.3 0.00174412 0 0.0017440399999999999 0 0.00174414 3.3 0.00174406 3.3 0.00174416 0 0.0017440799999999998 0 0.00174418 3.3 0.0017441 3.3 0.0017442 0 0.0017441199999999998 0 0.0017442199999999999 3.3 0.00174414 3.3 0.00174424 0 0.0017441599999999998 0 0.0017442599999999999 3.3 0.00174418 3.3 0.00174428 0 0.0017442 0 0.0017443 3.3 0.0017442199999999999 3.3 0.00174432 0 0.00174424 0 0.00174434 3.3 0.0017442599999999999 3.3 0.00174436 0 0.00174428 0 0.00174438 3.3 0.0017442999999999998 3.3 0.0017444 0 0.00174432 0 0.00174442 3.3 0.0017443399999999998 3.3 0.0017444399999999999 0 0.00174436 0 0.00174446 3.3 0.0017443799999999998 3.3 0.0017444799999999999 0 0.0017444 0 0.0017445 3.3 0.00174442 3.3 0.00174452 0 0.0017444399999999999 0 0.00174454 3.3 0.00174446 3.3 0.00174456 0 0.0017444799999999999 0 0.00174458 3.3 0.0017445 3.3 0.0017446 0 0.0017445199999999998 0 0.00174462 3.3 0.00174454 3.3 0.00174464 0 0.0017445599999999998 0 0.0017446599999999999 3.3 0.00174458 3.3 0.00174468 0 0.0017446 0 0.0017447 3.3 0.00174462 3.3 0.00174472 0 0.00174464 0 0.00174474 3.3 0.0017446599999999999 3.3 0.00174476 0 0.00174468 0 0.00174478 3.3 0.0017446999999999999 3.3 0.0017448 0 0.00174472 0 0.00174482 3.3 0.0017447399999999998 3.3 0.0017448399999999999 0 0.00174476 0 0.00174486 3.3 0.0017447799999999998 3.3 0.0017448799999999999 0 0.0017448 0 0.0017449 3.3 0.00174482 3.3 0.00174492 0 0.0017448399999999999 0 0.00174494 3.3 0.00174486 3.3 0.00174496 0 0.0017448799999999999 0 0.00174498 3.3 0.0017449 3.3 0.001745 0 0.0017449199999999998 0 0.00174502 3.3 0.00174494 3.3 0.00174504 0 0.0017449599999999998 0 0.0017450599999999999 3.3 0.00174498 3.3 0.00174508 0 0.0017449999999999998 0 0.0017450999999999999 3.3 0.00174502 3.3 0.00174512 0 0.00174504 0 0.00174514 3.3 0.0017450599999999999 3.3 0.00174516 0 0.00174508 0 0.00174518 3.3 0.0017450999999999999 3.3 0.0017452 0 0.00174512 0 0.00174522 3.3 0.0017451399999999998 3.3 0.00174524 0 0.00174516 0 0.00174526 3.3 0.0017451799999999998 3.3 0.0017452799999999999 0 0.0017452 0 0.0017453 3.3 0.0017452199999999998 3.3 0.0017453199999999999 0 0.00174524 0 0.00174534 3.3 0.00174526 3.3 0.00174536 0 0.0017452799999999999 0 0.00174538 3.3 0.0017453 3.3 0.0017454 0 0.0017453199999999999 0 0.00174542 3.3 0.00174534 3.3 0.00174544 0 0.0017453599999999998 0 0.00174546 3.3 0.00174538 3.3 0.00174548 0 0.0017453999999999998 0 0.0017454999999999999 3.3 0.00174542 3.3 0.00174552 0 0.00174544 0 0.00174554 3.3 0.00174546 3.3 0.00174556 0 0.00174548 0 0.00174558 3.3 0.0017454999999999999 3.3 0.0017456 0 0.00174552 0 0.00174562 3.3 0.0017455399999999999 3.3 0.00174564 0 0.00174556 0 0.00174566 3.3 0.0017455799999999998 3.3 0.0017456799999999999 0 0.0017456 0 0.0017457 3.3 0.0017456199999999998 3.3 0.0017457199999999999 0 0.00174564 0 0.00174574 3.3 0.00174566 3.3 0.00174576 0 0.0017456799999999999 0 0.00174578 3.3 0.0017457 3.3 0.0017458 0 0.0017457199999999999 0 0.00174582 3.3 0.00174574 3.3 0.00174584 0 0.0017457599999999998 0 0.00174586 3.3 0.00174578 3.3 0.00174588 0 0.0017457999999999998 0 0.0017458999999999999 3.3 0.00174582 3.3 0.00174592 0 0.0017458399999999998 0 0.0017459399999999999 3.3 0.00174586 3.3 0.00174596 0 0.00174588 0 0.00174598 3.3 0.0017458999999999999 3.3 0.001746 0 0.00174592 0 0.00174602 3.3 0.0017459399999999999 3.3 0.00174604 0 0.00174596 0 0.00174606 3.3 0.0017459799999999998 3.3 0.00174608 0 0.001746 0 0.0017461 3.3 0.0017460199999999998 3.3 0.0017461199999999999 0 0.00174604 0 0.00174614 3.3 0.00174606 3.3 0.00174616 0 0.00174608 0 0.00174618 3.3 0.0017461 3.3 0.0017462 0 0.0017461199999999999 0 0.00174622 3.3 0.00174614 3.3 0.00174624 0 0.0017461599999999999 0 0.00174626 3.3 0.00174618 3.3 0.00174628 0 0.0017461999999999998 0 0.0017463 3.3 0.00174622 3.3 0.00174632 0 0.0017462399999999998 0 0.0017463399999999999 3.3 0.00174626 3.3 0.00174636 0 0.00174628 0 0.00174638 3.3 0.0017463 3.3 0.0017464 0 0.00174632 0 0.00174642 3.3 0.0017463399999999999 3.3 0.00174644 0 0.00174636 0 0.00174646 3.3 0.0017463799999999999 3.3 0.00174648 0 0.0017464 0 0.0017465 3.3 0.0017464199999999998 3.3 0.0017465199999999999 0 0.00174644 0 0.00174654 3.3 0.0017464599999999998 3.3 0.0017465599999999999 0 0.00174648 0 0.00174658 3.3 0.0017465 3.3 0.0017466 0 0.0017465199999999999 0 0.00174662 3.3 0.00174654 3.3 0.00174664 0 0.0017465599999999999 0 0.00174666 3.3 0.00174658 3.3 0.00174668 0 0.0017465999999999998 0 0.0017467 3.3 0.00174662 3.3 0.00174672 0 0.0017466399999999998 0 0.0017467399999999999 3.3 0.00174666 3.3 0.00174676 0 0.0017466799999999998 0 0.0017467799999999999 3.3 0.0017467 3.3 0.0017468 0 0.00174672 0 0.00174682 3.3 0.0017467399999999999 3.3 0.00174684 0 0.00174676 0 0.00174686 3.3 0.0017467799999999999 3.3 0.00174688 0 0.0017468 0 0.0017469 3.3 0.0017468199999999998 3.3 0.00174692 0 0.00174684 0 0.00174694 3.3 0.0017468599999999998 3.3 0.0017469599999999999 0 0.00174688 0 0.00174698 3.3 0.0017469 3.3 0.001747 0 0.00174692 0 0.00174702 3.3 0.00174694 3.3 0.00174704 0 0.0017469599999999999 0 0.00174706 3.3 0.00174698 3.3 0.00174708 0 0.0017469999999999999 0 0.0017471 3.3 0.00174702 3.3 0.00174712 0 0.0017470399999999998 0 0.0017471399999999999 3.3 0.00174706 3.3 0.00174716 0 0.0017470799999999998 0 0.0017471799999999999 3.3 0.0017471 3.3 0.0017472 0 0.00174712 0 0.00174722 3.3 0.0017471399999999999 3.3 0.00174724 0 0.00174716 0 0.00174726 3.3 0.0017471799999999999 3.3 0.00174728 0 0.0017472 0 0.0017473 3.3 0.0017472199999999998 3.3 0.00174732 0 0.00174724 0 0.00174734 3.3 0.0017472599999999998 3.3 0.0017473599999999999 0 0.00174728 0 0.00174738 3.3 0.0017472999999999998 3.3 0.0017473999999999999 0 0.00174732 0 0.00174742 3.3 0.00174734 3.3 0.00174744 0 0.0017473599999999999 0 0.00174746 3.3 0.00174738 3.3 0.00174748 0 0.0017473999999999999 0 0.0017475 3.3 0.00174742 3.3 0.00174752 0 0.0017474399999999998 0 0.00174754 3.3 0.00174746 3.3 0.00174756 0 0.0017474799999999998 0 0.0017475799999999999 3.3 0.0017475 3.3 0.0017476 0 0.0017475199999999998 0 0.0017476199999999999 3.3 0.00174754 3.3 0.00174764 0 0.00174756 0 0.00174766 3.3 0.0017475799999999999 3.3 0.00174768 0 0.0017476 0 0.0017477 3.3 0.0017476199999999999 3.3 0.00174772 0 0.00174764 0 0.00174774 3.3 0.0017476599999999998 3.3 0.00174776 0 0.00174768 0 0.00174778 3.3 0.0017476999999999998 3.3 0.0017477999999999999 0 0.00174772 0 0.00174782 3.3 0.00174774 3.3 0.00174784 0 0.00174776 0 0.00174786 3.3 0.00174778 3.3 0.00174788 0 0.0017477999999999999 0 0.0017479 3.3 0.00174782 3.3 0.00174792 0 0.0017478399999999999 0 0.00174794 3.3 0.00174786 3.3 0.00174796 0 0.0017478799999999998 0 0.0017479799999999999 3.3 0.0017479 3.3 0.001748 0 0.0017479199999999998 0 0.0017480199999999999 3.3 0.00174794 3.3 0.00174804 0 0.00174796 0 0.00174806 3.3 0.0017479799999999999 3.3 0.00174808 0 0.001748 0 0.0017481 3.3 0.0017480199999999999 3.3 0.00174812 0 0.00174804 0 0.00174814 3.3 0.0017480599999999998 3.3 0.00174816 0 0.00174808 0 0.00174818 3.3 0.0017480999999999998 3.3 0.0017481999999999999 0 0.00174812 0 0.00174822 3.3 0.0017481399999999998 3.3 0.0017482399999999999 0 0.00174816 0 0.00174826 3.3 0.00174818 3.3 0.00174828 0 0.0017481999999999999 0 0.0017483 3.3 0.00174822 3.3 0.00174832 0 0.0017482399999999999 0 0.00174834 3.3 0.00174826 3.3 0.00174836 0 0.0017482799999999998 0 0.00174838 3.3 0.0017483 3.3 0.0017484 0 0.0017483199999999998 0 0.0017484199999999999 3.3 0.00174834 3.3 0.00174844 0 0.0017483599999999998 0 0.0017484599999999999 3.3 0.00174838 3.3 0.00174848 0 0.0017484 0 0.0017485 3.3 0.0017484199999999999 3.3 0.00174852 0 0.00174844 0 0.00174854 3.3 0.0017484599999999999 3.3 0.00174856 0 0.00174848 0 0.00174858 3.3 0.0017484999999999998 3.3 0.0017486 0 0.00174852 0 0.00174862 3.3 0.0017485399999999998 3.3 0.0017486399999999999 0 0.00174856 0 0.00174866 3.3 0.00174858 3.3 0.00174868 0 0.0017486 0 0.0017487 3.3 0.00174862 3.3 0.00174872 0 0.0017486399999999999 0 0.00174874 3.3 0.00174866 3.3 0.00174876 0 0.0017486799999999999 0 0.00174878 3.3 0.0017487 3.3 0.0017488 0 0.0017487199999999998 0 0.0017488199999999999 3.3 0.00174874 3.3 0.00174884 0 0.0017487599999999998 0 0.0017488599999999999 3.3 0.00174878 3.3 0.00174888 0 0.0017488 0 0.0017489 3.3 0.0017488199999999999 3.3 0.00174892 0 0.00174884 0 0.00174894 3.3 0.0017488599999999999 3.3 0.00174896 0 0.00174888 0 0.00174898 3.3 0.0017488999999999998 3.3 0.001749 0 0.00174892 0 0.00174902 3.3 0.0017489399999999998 3.3 0.0017490399999999999 0 0.00174896 0 0.00174906 3.3 0.0017489799999999998 3.3 0.0017490799999999999 0 0.001749 0 0.0017491 3.3 0.00174902 3.3 0.00174912 0 0.0017490399999999999 0 0.00174914 3.3 0.00174906 3.3 0.00174916 0 0.0017490799999999999 0 0.00174918 3.3 0.0017491 3.3 0.0017492 0 0.0017491199999999998 0 0.00174922 3.3 0.00174914 3.3 0.00174924 0 0.0017491599999999998 0 0.0017492599999999999 3.3 0.00174918 3.3 0.00174928 0 0.0017491999999999998 0 0.0017492999999999999 3.3 0.00174922 3.3 0.00174932 0 0.00174924 0 0.00174934 3.3 0.0017492599999999999 3.3 0.00174936 0 0.00174928 0 0.00174938 3.3 0.0017492999999999999 3.3 0.0017494 0 0.00174932 0 0.00174942 3.3 0.0017493399999999998 3.3 0.00174944 0 0.00174936 0 0.00174946 3.3 0.0017493799999999998 3.3 0.0017494799999999999 0 0.0017494 0 0.0017495 3.3 0.00174942 3.3 0.00174952 0 0.00174944 0 0.00174954 3.3 0.00174946 3.3 0.00174956 0 0.0017494799999999999 0 0.00174958 3.3 0.0017495 3.3 0.0017496 0 0.0017495199999999999 0 0.00174962 3.3 0.00174954 3.3 0.00174964 0 0.0017495599999999998 0 0.0017496599999999999 3.3 0.00174958 3.3 0.00174968 0 0.0017495999999999998 0 0.0017496999999999999 3.3 0.00174962 3.3 0.00174972 0 0.00174964 0 0.00174974 3.3 0.0017496599999999999 3.3 0.00174976 0 0.00174968 0 0.00174978 3.3 0.0017496999999999999 3.3 0.0017498 0 0.00174972 0 0.00174982 3.3 0.0017497399999999998 3.3 0.00174984 0 0.00174976 0 0.00174986 3.3 0.0017497799999999998 3.3 0.0017498799999999999 0 0.0017498 0 0.0017499 3.3 0.0017498199999999998 3.3 0.0017499199999999999 0 0.00174984 0 0.00174994 3.3 0.00174986 3.3 0.00174996 0 0.0017498799999999999 0 0.00174998 3.3 0.0017499 3.3 0.00175 0 0.0017499199999999999 0 0.00175002 3.3 0.00174994 3.3 0.00175004 0 0.0017499599999999998 0 0.00175006 3.3 0.00174998 3.3 0.00175008 0 0.0017499999999999998 0 0.0017500999999999999 3.3 0.00175002 3.3 0.00175012 0 0.00175004 0 0.00175014 3.3 0.00175006 3.3 0.00175016 0 0.00175008 0 0.00175018 3.3 0.0017500999999999999 3.3 0.0017502 0 0.00175012 0 0.00175022 3.3 0.0017501399999999999 3.3 0.00175024 0 0.00175016 0 0.00175026 3.3 0.0017501799999999998 3.3 0.0017502799999999999 0 0.0017502 0 0.0017503 3.3 0.0017502199999999998 3.3 0.0017503199999999999 0 0.00175024 0 0.00175034 3.3 0.00175026 3.3 0.00175036 0 0.0017502799999999999 0 0.00175038 3.3 0.0017503 3.3 0.0017504 0 0.0017503199999999999 0 0.00175042 3.3 0.00175034 3.3 0.00175044 0 0.0017503599999999999 0 0.00175046 3.3 0.00175038 3.3 0.00175048 0 0.0017503999999999998 0 0.0017504999999999999 3.3 0.00175042 3.3 0.00175052 0 0.0017504399999999998 0 0.0017505399999999999 3.3 0.00175046 3.3 0.00175056 0 0.00175048 0 0.00175058 3.3 0.0017504999999999999 3.3 0.0017506 0 0.00175052 0 0.00175062 3.3 0.0017505399999999999 3.3 0.00175064 0 0.00175056 0 0.00175066 3.3 0.0017505799999999998 3.3 0.00175068 0 0.0017506 0 0.0017507 3.3 0.0017506199999999998 3.3 0.0017507199999999999 0 0.00175064 0 0.00175074 3.3 0.0017506599999999998 3.3 0.0017507599999999999 0 0.00175068 0 0.00175078 3.3 0.0017507 3.3 0.0017508 0 0.0017507199999999999 0 0.00175082 3.3 0.00175074 3.3 0.00175084 0 0.0017507599999999999 0 0.00175086 3.3 0.00175078 3.3 0.00175088 0 0.0017507999999999998 0 0.0017509 3.3 0.00175082 3.3 0.00175092 0 0.0017508399999999998 0 0.0017509399999999999 3.3 0.00175086 3.3 0.00175096 0 0.00175088 0 0.00175098 3.3 0.0017509 3.3 0.001751 0 0.00175092 0 0.00175102 3.3 0.0017509399999999999 3.3 0.00175104 0 0.00175096 0 0.00175106 3.3 0.0017509799999999999 3.3 0.00175108 0 0.001751 0 0.0017511 3.3 0.0017510199999999998 3.3 0.0017511199999999999 0 0.00175104 0 0.00175114 3.3 0.0017510599999999998 3.3 0.0017511599999999999 0 0.00175108 0 0.00175118 3.3 0.0017511 3.3 0.0017512 0 0.0017511199999999999 0 0.00175122 3.3 0.00175114 3.3 0.00175124 0 0.0017511599999999999 0 0.00175126 3.3 0.00175118 3.3 0.00175128 0 0.0017511999999999998 0 0.0017513 3.3 0.00175122 3.3 0.00175132 0 0.0017512399999999998 0 0.0017513399999999999 3.3 0.00175126 3.3 0.00175136 0 0.0017512799999999998 0 0.0017513799999999999 3.3 0.0017513 3.3 0.0017514 0 0.00175132 0 0.00175142 3.3 0.0017513399999999999 3.3 0.00175144 0 0.00175136 0 0.00175146 3.3 0.0017513799999999999 3.3 0.00175148 0 0.0017514 0 0.0017515 3.3 0.0017514199999999998 3.3 0.00175152 0 0.00175144 0 0.00175154 3.3 0.0017514599999999998 3.3 0.0017515599999999999 0 0.00175148 0 0.00175158 3.3 0.0017514999999999998 3.3 0.0017515999999999999 0 0.00175152 0 0.00175162 3.3 0.00175154 3.3 0.00175164 0 0.0017515599999999999 0 0.00175166 3.3 0.00175158 3.3 0.00175168 0 0.0017515999999999999 0 0.0017517 3.3 0.00175162 3.3 0.00175172 0 0.0017516399999999998 0 0.00175174 3.3 0.00175166 3.3 0.00175176 0 0.0017516799999999998 0 0.0017517799999999999 3.3 0.0017517 3.3 0.0017518 0 0.00175172 0 0.00175182 3.3 0.00175174 3.3 0.00175184 0 0.00175176 0 0.00175186 3.3 0.0017517799999999999 3.3 0.00175188 0 0.0017518 0 0.0017519 3.3 0.0017518199999999999 3.3 0.00175192 0 0.00175184 0 0.00175194 3.3 0.0017518599999999998 3.3 0.0017519599999999999 0 0.00175188 0 0.00175198 3.3 0.0017518999999999998 3.3 0.0017519999999999999 0 0.00175192 0 0.00175202 3.3 0.00175194 3.3 0.00175204 0 0.0017519599999999999 0 0.00175206 3.3 0.00175198 3.3 0.00175208 0 0.0017519999999999999 0 0.0017521 3.3 0.00175202 3.3 0.00175212 0 0.0017520399999999998 0 0.00175214 3.3 0.00175206 3.3 0.00175216 0 0.0017520799999999998 0 0.0017521799999999999 3.3 0.0017521 3.3 0.0017522 0 0.0017521199999999998 0 0.0017522199999999999 3.3 0.00175214 3.3 0.00175224 0 0.00175216 0 0.00175226 3.3 0.0017521799999999999 3.3 0.00175228 0 0.0017522 0 0.0017523 3.3 0.0017522199999999999 3.3 0.00175232 0 0.00175224 0 0.00175234 3.3 0.0017522599999999998 3.3 0.00175236 0 0.00175228 0 0.00175238 3.3 0.0017522999999999998 3.3 0.0017523999999999999 0 0.00175232 0 0.00175242 3.3 0.0017523399999999998 3.3 0.0017524399999999999 0 0.00175236 0 0.00175246 3.3 0.00175238 3.3 0.00175248 0 0.0017523999999999999 0 0.0017525 3.3 0.00175242 3.3 0.00175252 0 0.0017524399999999999 0 0.00175254 3.3 0.00175246 3.3 0.00175256 0 0.0017524799999999998 0 0.00175258 3.3 0.0017525 3.3 0.0017526 0 0.0017525199999999998 0 0.0017526199999999999 3.3 0.00175254 3.3 0.00175264 0 0.00175256 0 0.00175266 3.3 0.00175258 3.3 0.00175268 0 0.0017526 0 0.0017527 3.3 0.0017526199999999999 3.3 0.00175272 0 0.00175264 0 0.00175274 3.3 0.0017526599999999999 3.3 0.00175276 0 0.00175268 0 0.00175278 3.3 0.0017526999999999998 3.3 0.0017527999999999999 0 0.00175272 0 0.00175282 3.3 0.0017527399999999998 3.3 0.0017528399999999999 0 0.00175276 0 0.00175286 3.3 0.00175278 3.3 0.00175288 0 0.0017527999999999999 0 0.0017529 3.3 0.00175282 3.3 0.00175292 0 0.0017528399999999999 0 0.00175294 3.3 0.00175286 3.3 0.00175296 0 0.0017528799999999998 0 0.00175298 3.3 0.0017529 3.3 0.001753 0 0.0017529199999999998 0 0.0017530199999999999 3.3 0.00175294 3.3 0.00175304 0 0.0017529599999999998 0 0.0017530599999999999 3.3 0.00175298 3.3 0.00175308 0 0.001753 0 0.0017531 3.3 0.0017530199999999999 3.3 0.00175312 0 0.00175304 0 0.00175314 3.3 0.0017530599999999999 3.3 0.00175316 0 0.00175308 0 0.00175318 3.3 0.0017530999999999998 3.3 0.0017532 0 0.00175312 0 0.00175322 3.3 0.0017531399999999998 3.3 0.0017532399999999999 0 0.00175316 0 0.00175326 3.3 0.00175318 3.3 0.00175328 0 0.0017532 0 0.0017533 3.3 0.00175322 3.3 0.00175332 0 0.0017532399999999999 0 0.00175334 3.3 0.00175326 3.3 0.00175336 0 0.0017532799999999999 0 0.00175338 3.3 0.0017533 3.3 0.0017534 0 0.0017533199999999998 0 0.00175342 3.3 0.00175334 3.3 0.00175344 0 0.0017533599999999998 0 0.0017534599999999999 3.3 0.00175338 3.3 0.00175348 0 0.0017534 0 0.0017535 3.3 0.00175342 3.3 0.00175352 0 0.00175344 0 0.00175354 3.3 0.0017534599999999999 3.3 0.00175356 0 0.00175348 0 0.00175358 3.3 0.0017534999999999999 3.3 0.0017536 0 0.00175352 0 0.00175362 3.3 0.0017535399999999998 3.3 0.0017536399999999999 0 0.00175356 0 0.00175366 3.3 0.0017535799999999998 3.3 0.0017536799999999999 0 0.0017536 0 0.0017537 3.3 0.00175362 3.3 0.00175372 0 0.0017536399999999999 0 0.00175374 3.3 0.00175366 3.3 0.00175376 0 0.0017536799999999999 0 0.00175378 3.3 0.0017537 3.3 0.0017538 0 0.0017537199999999998 0 0.00175382 3.3 0.00175374 3.3 0.00175384 0 0.0017537599999999998 0 0.0017538599999999999 3.3 0.00175378 3.3 0.00175388 0 0.0017537999999999998 0 0.0017538999999999999 3.3 0.00175382 3.3 0.00175392 0 0.00175384 0 0.00175394 3.3 0.0017538599999999999 3.3 0.00175396 0 0.00175388 0 0.00175398 3.3 0.0017538999999999999 3.3 0.001754 0 0.00175392 0 0.00175402 3.3 0.0017539399999999998 3.3 0.00175404 0 0.00175396 0 0.00175406 3.3 0.0017539799999999998 3.3 0.0017540799999999999 0 0.001754 0 0.0017541 3.3 0.00175402 3.3 0.00175412 0 0.00175404 0 0.00175414 3.3 0.00175406 3.3 0.00175416 0 0.0017540799999999999 0 0.00175418 3.3 0.0017541 3.3 0.0017542 0 0.0017541199999999999 0 0.00175422 3.3 0.00175414 3.3 0.00175424 0 0.0017541599999999998 0 0.0017542599999999999 3.3 0.00175418 3.3 0.00175428 0 0.0017541999999999998 0 0.0017542999999999999 3.3 0.00175422 3.3 0.00175432 0 0.00175424 0 0.00175434 3.3 0.0017542599999999999 3.3 0.00175436 0 0.00175428 0 0.00175438 3.3 0.0017542999999999999 3.3 0.0017544 0 0.00175432 0 0.00175442 3.3 0.0017543399999999998 3.3 0.00175444 0 0.00175436 0 0.00175446 3.3 0.0017543799999999998 3.3 0.0017544799999999999 0 0.0017544 0 0.0017545 3.3 0.0017544199999999998 3.3 0.0017545199999999999 0 0.00175444 0 0.00175454 3.3 0.00175446 3.3 0.00175456 0 0.0017544799999999999 0 0.00175458 3.3 0.0017545 3.3 0.0017546 0 0.0017545199999999999 0 0.00175462 3.3 0.00175454 3.3 0.00175464 0 0.0017545599999999998 0 0.00175466 3.3 0.00175458 3.3 0.00175468 0 0.0017545999999999998 0 0.0017546999999999999 3.3 0.00175462 3.3 0.00175472 0 0.0017546399999999998 0 0.0017547399999999999 3.3 0.00175466 3.3 0.00175476 0 0.00175468 0 0.00175478 3.3 0.0017546999999999999 3.3 0.0017548 0 0.00175472 0 0.00175482 3.3 0.0017547399999999999 3.3 0.00175484 0 0.00175476 0 0.00175486 3.3 0.0017547799999999998 3.3 0.00175488 0 0.0017548 0 0.0017549 3.3 0.0017548199999999998 3.3 0.0017549199999999999 0 0.00175484 0 0.00175494 3.3 0.00175486 3.3 0.00175496 0 0.00175488 0 0.00175498 3.3 0.0017549 3.3 0.001755 0 0.0017549199999999999 0 0.00175502 3.3 0.00175494 3.3 0.00175504 0 0.0017549599999999999 0 0.00175506 3.3 0.00175498 3.3 0.00175508 0 0.0017549999999999998 0 0.0017550999999999999 3.3 0.00175502 3.3 0.00175512 0 0.0017550399999999998 0 0.0017551399999999999 3.3 0.00175506 3.3 0.00175516 0 0.00175508 0 0.00175518 3.3 0.0017550999999999999 3.3 0.0017552 0 0.00175512 0 0.00175522 3.3 0.0017551399999999999 3.3 0.00175524 0 0.00175516 0 0.00175526 3.3 0.0017551799999999998 3.3 0.00175528 0 0.0017552 0 0.0017553 3.3 0.0017552199999999998 3.3 0.0017553199999999999 0 0.00175524 0 0.00175534 3.3 0.0017552599999999998 3.3 0.0017553599999999999 0 0.00175528 0 0.00175538 3.3 0.0017553 3.3 0.0017554 0 0.0017553199999999999 0 0.00175542 3.3 0.00175534 3.3 0.00175544 0 0.0017553599999999999 0 0.00175546 3.3 0.00175538 3.3 0.00175548 0 0.0017553999999999998 0 0.0017555 3.3 0.00175542 3.3 0.00175552 0 0.0017554399999999998 0 0.0017555399999999999 3.3 0.00175546 3.3 0.00175556 0 0.0017554799999999998 0 0.0017555799999999999 3.3 0.0017555 3.3 0.0017556 0 0.00175552 0 0.00175562 3.3 0.0017555399999999999 3.3 0.00175564 0 0.00175556 0 0.00175566 3.3 0.0017555799999999999 3.3 0.00175568 0 0.0017556 0 0.0017557 3.3 0.0017556199999999998 3.3 0.00175572 0 0.00175564 0 0.00175574 3.3 0.0017556599999999998 3.3 0.0017557599999999999 0 0.00175568 0 0.00175578 3.3 0.0017557 3.3 0.0017558 0 0.00175572 0 0.00175582 3.3 0.00175574 3.3 0.00175584 0 0.0017557599999999999 0 0.00175586 3.3 0.00175578 3.3 0.00175588 0 0.0017557999999999999 0 0.0017559 3.3 0.00175582 3.3 0.00175592 0 0.0017558399999999998 0 0.0017559399999999999 3.3 0.00175586 3.3 0.00175596 0 0.0017558799999999998 0 0.0017559799999999999 3.3 0.0017559 3.3 0.001756 0 0.00175592 0 0.00175602 3.3 0.0017559399999999999 3.3 0.00175604 0 0.00175596 0 0.00175606 3.3 0.0017559799999999999 3.3 0.00175608 0 0.001756 0 0.0017561 3.3 0.0017560199999999998 3.3 0.00175612 0 0.00175604 0 0.00175614 3.3 0.0017560599999999998 3.3 0.0017561599999999999 0 0.00175608 0 0.00175618 3.3 0.0017560999999999998 3.3 0.0017561999999999999 0 0.00175612 0 0.00175622 3.3 0.00175614 3.3 0.00175624 0 0.0017561599999999999 0 0.00175626 3.3 0.00175618 3.3 0.00175628 0 0.0017561999999999999 0 0.0017563 3.3 0.00175622 3.3 0.00175632 0 0.0017562399999999998 0 0.00175634 3.3 0.00175626 3.3 0.00175636 0 0.0017562799999999998 0 0.0017563799999999999 3.3 0.0017563 3.3 0.0017564 0 0.0017563199999999998 0 0.0017564199999999999 3.3 0.00175634 3.3 0.00175644 0 0.00175636 0 0.00175646 3.3 0.0017563799999999999 3.3 0.00175648 0 0.0017564 0 0.0017565 3.3 0.0017564199999999999 3.3 0.00175652 0 0.00175644 0 0.00175654 3.3 0.0017564599999999998 3.3 0.00175656 0 0.00175648 0 0.00175658 3.3 0.0017564999999999998 3.3 0.0017565999999999999 0 0.00175652 0 0.00175662 3.3 0.00175654 3.3 0.00175664 0 0.00175656 0 0.00175666 3.3 0.00175658 3.3 0.00175668 0 0.0017565999999999999 0 0.0017567 3.3 0.00175662 3.3 0.00175672 0 0.0017566399999999999 0 0.00175674 3.3 0.00175666 3.3 0.00175676 0 0.0017566799999999998 0 0.0017567799999999999 3.3 0.0017567 3.3 0.0017568 0 0.0017567199999999998 0 0.0017568199999999999 3.3 0.00175674 3.3 0.00175684 0 0.00175676 0 0.00175686 3.3 0.0017567799999999999 3.3 0.00175688 0 0.0017568 0 0.0017569 3.3 0.0017568199999999999 3.3 0.00175692 0 0.00175684 0 0.00175694 3.3 0.0017568599999999998 3.3 0.00175696 0 0.00175688 0 0.00175698 3.3 0.0017568999999999998 3.3 0.0017569999999999999 0 0.00175692 0 0.00175702 3.3 0.0017569399999999998 3.3 0.0017570399999999999 0 0.00175696 0 0.00175706 3.3 0.00175698 3.3 0.00175708 0 0.0017569999999999999 0 0.0017571 3.3 0.00175702 3.3 0.00175712 0 0.0017570399999999999 0 0.00175714 3.3 0.00175706 3.3 0.00175716 0 0.0017570799999999998 0 0.00175718 3.3 0.0017571 3.3 0.0017572 0 0.0017571199999999998 0 0.0017572199999999999 3.3 0.00175714 3.3 0.00175724 0 0.00175716 0 0.00175726 3.3 0.00175718 3.3 0.00175728 0 0.0017572 0 0.0017573 3.3 0.0017572199999999999 3.3 0.00175732 0 0.00175724 0 0.00175734 3.3 0.0017572599999999999 3.3 0.00175736 0 0.00175728 0 0.00175738 3.3 0.0017572999999999998 3.3 0.0017573999999999999 0 0.00175732 0 0.00175742 3.3 0.0017573399999999998 3.3 0.0017574399999999999 0 0.00175736 0 0.00175746 3.3 0.00175738 3.3 0.00175748 0 0.0017573999999999999 0 0.0017575 3.3 0.00175742 3.3 0.00175752 0 0.0017574399999999999 0 0.00175754 3.3 0.00175746 3.3 0.00175756 0 0.0017574799999999998 0 0.00175758 3.3 0.0017575 3.3 0.0017576 0 0.0017575199999999998 0 0.0017576199999999999 3.3 0.00175754 3.3 0.00175764 0 0.0017575599999999998 0 0.0017576599999999999 3.3 0.00175758 3.3 0.00175768 0 0.0017576 0 0.0017577 3.3 0.0017576199999999999 3.3 0.00175772 0 0.00175764 0 0.00175774 3.3 0.0017576599999999999 3.3 0.00175776 0 0.00175768 0 0.00175778 3.3 0.0017576999999999998 3.3 0.0017578 0 0.00175772 0 0.00175782 3.3 0.0017577399999999998 3.3 0.0017578399999999999 0 0.00175776 0 0.00175786 3.3 0.0017577799999999998 3.3 0.0017578799999999999 0 0.0017578 0 0.0017579 3.3 0.00175782 3.3 0.00175792 0 0.0017578399999999999 0 0.00175794 3.3 0.00175786 3.3 0.00175796 0 0.0017578799999999999 0 0.00175798 3.3 0.0017579 3.3 0.001758 0 0.0017579199999999998 0 0.00175802 3.3 0.00175794 3.3 0.00175804 0 0.0017579599999999998 0 0.0017580599999999999 3.3 0.00175798 3.3 0.00175808 0 0.001758 0 0.0017581 3.3 0.00175802 3.3 0.00175812 0 0.00175804 0 0.00175814 3.3 0.0017580599999999999 3.3 0.00175816 0 0.00175808 0 0.00175818 3.3 0.0017580999999999999 3.3 0.0017582 0 0.00175812 0 0.00175822 3.3 0.0017581399999999998 3.3 0.0017582399999999999 0 0.00175816 0 0.00175826 3.3 0.0017581799999999998 3.3 0.0017582799999999999 0 0.0017582 0 0.0017583 3.3 0.00175822 3.3 0.00175832 0 0.0017582399999999999 0 0.00175834 3.3 0.00175826 3.3 0.00175836 0 0.0017582799999999999 0 0.00175838 3.3 0.0017583 3.3 0.0017584 0 0.0017583199999999998 0 0.00175842 3.3 0.00175834 3.3 0.00175844 0 0.0017583599999999998 0 0.0017584599999999999 3.3 0.00175838 3.3 0.00175848 0 0.0017583999999999998 0 0.0017584999999999999 3.3 0.00175842 3.3 0.00175852 0 0.00175844 0 0.00175854 3.3 0.0017584599999999999 3.3 0.00175856 0 0.00175848 0 0.00175858 3.3 0.0017584999999999999 3.3 0.0017586 0 0.00175852 0 0.00175862 3.3 0.0017585399999999998 3.3 0.00175864 0 0.00175856 0 0.00175866 3.3 0.0017585799999999998 3.3 0.0017586799999999999 0 0.0017586 0 0.0017587 3.3 0.0017586199999999998 3.3 0.0017587199999999999 0 0.00175864 0 0.00175874 3.3 0.00175866 3.3 0.00175876 0 0.0017586799999999999 0 0.00175878 3.3 0.0017587 3.3 0.0017588 0 0.0017587199999999999 0 0.00175882 3.3 0.00175874 3.3 0.00175884 0 0.0017587599999999998 0 0.00175886 3.3 0.00175878 3.3 0.00175888 0 0.0017587999999999998 0 0.0017588999999999999 3.3 0.00175882 3.3 0.00175892 0 0.00175884 0 0.00175894 3.3 0.00175886 3.3 0.00175896 0 0.00175888 0 0.00175898 3.3 0.0017588999999999999 3.3 0.001759 0 0.00175892 0 0.00175902 3.3 0.0017589399999999999 3.3 0.00175904 0 0.00175896 0 0.00175906 3.3 0.0017589799999999998 3.3 0.0017590799999999999 0 0.001759 0 0.0017591 3.3 0.0017590199999999998 3.3 0.0017591199999999999 0 0.00175904 0 0.00175914 3.3 0.00175906 3.3 0.00175916 0 0.0017590799999999999 0 0.00175918 3.3 0.0017591 3.3 0.0017592 0 0.0017591199999999999 0 0.00175922 3.3 0.00175914 3.3 0.00175924 0 0.0017591599999999998 0 0.00175926 3.3 0.00175918 3.3 0.00175928 0 0.0017591999999999998 0 0.0017592999999999999 3.3 0.00175922 3.3 0.00175932 0 0.0017592399999999998 0 0.0017593399999999999 3.3 0.00175926 3.3 0.00175936 0 0.00175928 0 0.00175938 3.3 0.0017592999999999999 3.3 0.0017594 0 0.00175932 0 0.00175942 3.3 0.0017593399999999999 3.3 0.00175944 0 0.00175936 0 0.00175946 3.3 0.0017593799999999998 3.3 0.00175948 0 0.0017594 0 0.0017595 3.3 0.0017594199999999998 3.3 0.0017595199999999999 0 0.00175944 0 0.00175954 3.3 0.0017594599999999998 3.3 0.0017595599999999999 0 0.00175948 0 0.00175958 3.3 0.0017595 3.3 0.0017596 0 0.0017595199999999999 0 0.00175962 3.3 0.00175954 3.3 0.00175964 0 0.0017595599999999999 0 0.00175966 3.3 0.00175958 3.3 0.00175968 0 0.0017595999999999998 0 0.0017597 3.3 0.00175962 3.3 0.00175972 0 0.0017596399999999998 0 0.0017597399999999999 3.3 0.00175966 3.3 0.00175976 0 0.00175968 0 0.00175978 3.3 0.0017597 3.3 0.0017598 0 0.00175972 0 0.00175982 3.3 0.0017597399999999999 3.3 0.00175984 0 0.00175976 0 0.00175986 3.3 0.0017597799999999999 3.3 0.00175988 0 0.0017598 0 0.0017599 3.3 0.0017598199999999998 3.3 0.0017599199999999999 0 0.00175984 0 0.00175994 3.3 0.0017598599999999998 3.3 0.0017599599999999999 0 0.00175988 0 0.00175998 3.3 0.0017599 3.3 0.00176 0 0.0017599199999999999 0 0.00176002 3.3 0.00175994 3.3 0.00176004 0 0.0017599599999999999 0 0.00176006 3.3 0.00175998 3.3 0.00176008 0 0.0017599999999999998 0 0.0017601 3.3 0.00176002 3.3 0.00176012 0 0.0017600399999999998 0 0.0017601399999999999 3.3 0.00176006 3.3 0.00176016 0 0.0017600799999999998 0 0.0017601799999999999 3.3 0.0017601 3.3 0.0017602 0 0.00176012 0 0.00176022 3.3 0.0017601399999999999 3.3 0.00176024 0 0.00176016 0 0.00176026 3.3 0.0017601799999999999 3.3 0.00176028 0 0.0017602 0 0.0017603 3.3 0.0017602199999999998 3.3 0.00176032 0 0.00176024 0 0.00176034 3.3 0.0017602599999999998 3.3 0.0017603599999999999 0 0.00176028 0 0.00176038 3.3 0.0017603 3.3 0.0017604 0 0.00176032 0 0.00176042 3.3 0.00176034 3.3 0.00176044 0 0.0017603599999999999 0 0.00176046 3.3 0.00176038 3.3 0.00176048 0 0.0017603999999999999 0 0.0017605 3.3 0.00176042 3.3 0.00176052 0 0.0017604399999999998 0 0.0017605399999999999 3.3 0.00176046 3.3 0.00176056 0 0.0017604799999999998 0 0.0017605799999999999 3.3 0.0017605 3.3 0.0017606 0 0.00176052 0 0.00176062 3.3 0.0017605399999999999 3.3 0.00176064 0 0.00176056 0 0.00176066 3.3 0.0017605799999999999 3.3 0.00176068 0 0.0017606 0 0.0017607 3.3 0.0017606199999999999 3.3 0.00176072 0 0.00176064 0 0.00176074 3.3 0.0017606599999999998 3.3 0.0017607599999999999 0 0.00176068 0 0.00176078 3.3 0.0017606999999999998 3.3 0.0017607999999999999 0 0.00176072 0 0.00176082 3.3 0.00176074 3.3 0.00176084 0 0.0017607599999999999 0 0.00176086 3.3 0.00176078 3.3 0.00176088 0 0.0017607999999999999 0 0.0017609 3.3 0.00176082 3.3 0.00176092 0 0.0017608399999999998 0 0.00176094 3.3 0.00176086 3.3 0.00176096 0 0.0017608799999999998 0 0.0017609799999999999 3.3 0.0017609 3.3 0.001761 0 0.0017609199999999998 0 0.0017610199999999999 3.3 0.00176094 3.3 0.00176104 0 0.00176096 0 0.00176106 3.3 0.0017609799999999999 3.3 0.00176108 0 0.001761 0 0.0017611 3.3 0.0017610199999999999 3.3 0.00176112 0 0.00176104 0 0.00176114 3.3 0.0017610599999999998 3.3 0.00176116 0 0.00176108 0 0.00176118 3.3 0.0017610999999999998 3.3 0.0017611999999999999 0 0.00176112 0 0.00176122 3.3 0.00176114 3.3 0.00176124 0 0.00176116 0 0.00176126 3.3 0.00176118 3.3 0.00176128 0 0.0017611999999999999 0 0.0017613 3.3 0.00176122 3.3 0.00176132 0 0.0017612399999999999 0 0.00176134 3.3 0.00176126 3.3 0.00176136 0 0.0017612799999999998 0 0.0017613799999999999 3.3 0.0017613 3.3 0.0017614 0 0.0017613199999999998 0 0.0017614199999999999 3.3 0.00176134 3.3 0.00176144 0 0.00176136 0 0.00176146 3.3 0.0017613799999999999 3.3 0.00176148 0 0.0017614 0 0.0017615 3.3 0.0017614199999999999 3.3 0.00176152 0 0.00176144 0 0.00176154 3.3 0.0017614599999999998 3.3 0.00176156 0 0.00176148 0 0.00176158 3.3 0.0017614999999999998 3.3 0.0017615999999999999 0 0.00176152 0 0.00176162 3.3 0.0017615399999999998 3.3 0.0017616399999999999 0 0.00176156 0 0.00176166 3.3 0.00176158 3.3 0.00176168 0 0.0017615999999999999 0 0.0017617 3.3 0.00176162 3.3 0.00176172 0 0.0017616399999999999 0 0.00176174 3.3 0.00176166 3.3 0.00176176 0 0.0017616799999999998 0 0.00176178 3.3 0.0017617 3.3 0.0017618 0 0.0017617199999999998 0 0.0017618199999999999 3.3 0.00176174 3.3 0.00176184 0 0.0017617599999999998 0 0.0017618599999999999 3.3 0.00176178 3.3 0.00176188 0 0.0017618 0 0.0017619 3.3 0.0017618199999999999 3.3 0.00176192 0 0.00176184 0 0.00176194 3.3 0.0017618599999999999 3.3 0.00176196 0 0.00176188 0 0.00176198 3.3 0.0017618999999999998 3.3 0.001762 0 0.00176192 0 0.00176202 3.3 0.0017619399999999998 3.3 0.0017620399999999999 0 0.00176196 0 0.00176206 3.3 0.00176198 3.3 0.00176208 0 0.001762 0 0.0017621 3.3 0.00176202 3.3 0.00176212 0 0.0017620399999999999 0 0.00176214 3.3 0.00176206 3.3 0.00176216 0 0.0017620799999999999 0 0.00176218 3.3 0.0017621 3.3 0.0017622 0 0.0017621199999999998 0 0.0017622199999999999 3.3 0.00176214 3.3 0.00176224 0 0.0017621599999999998 0 0.0017622599999999999 3.3 0.00176218 3.3 0.00176228 0 0.0017622 0 0.0017623 3.3 0.0017622199999999999 3.3 0.00176232 0 0.00176224 0 0.00176234 3.3 0.0017622599999999999 3.3 0.00176236 0 0.00176228 0 0.00176238 3.3 0.0017622999999999998 3.3 0.0017624 0 0.00176232 0 0.00176242 3.3 0.0017623399999999998 3.3 0.0017624399999999999 0 0.00176236 0 0.00176246 3.3 0.0017623799999999998 3.3 0.0017624799999999999 0 0.0017624 0 0.0017625 3.3 0.00176242 3.3 0.00176252 0 0.0017624399999999999 0 0.00176254 3.3 0.00176246 3.3 0.00176256 0 0.0017624799999999999 0 0.00176258 3.3 0.0017625 3.3 0.0017626 0 0.0017625199999999998 0 0.00176262 3.3 0.00176254 3.3 0.00176264 0 0.0017625599999999998 0 0.0017626599999999999 3.3 0.00176258 3.3 0.00176268 0 0.0017625999999999998 0 0.0017626999999999999 3.3 0.00176262 3.3 0.00176272 0 0.00176264 0 0.00176274 3.3 0.0017626599999999999 3.3 0.00176276 0 0.00176268 0 0.00176278 3.3 0.0017626999999999999 3.3 0.0017628 0 0.00176272 0 0.00176282 3.3 0.0017627399999999998 3.3 0.00176284 0 0.00176276 0 0.00176286 3.3 0.0017627799999999998 3.3 0.0017628799999999999 0 0.0017628 0 0.0017629 3.3 0.00176282 3.3 0.00176292 0 0.00176284 0 0.00176294 3.3 0.00176286 3.3 0.00176296 0 0.0017628799999999999 0 0.00176298 3.3 0.0017629 3.3 0.001763 0 0.0017629199999999999 0 0.00176302 3.3 0.00176294 3.3 0.00176304 0 0.0017629599999999998 0 0.0017630599999999999 3.3 0.00176298 3.3 0.00176308 0 0.0017629999999999998 0 0.0017630999999999999 3.3 0.00176302 3.3 0.00176312 0 0.00176304 0 0.00176314 3.3 0.0017630599999999999 3.3 0.00176316 0 0.00176308 0 0.00176318 3.3 0.0017630999999999999 3.3 0.0017632 0 0.00176312 0 0.00176322 3.3 0.0017631399999999998 3.3 0.00176324 0 0.00176316 0 0.00176326 3.3 0.0017631799999999998 3.3 0.0017632799999999999 0 0.0017632 0 0.0017633 3.3 0.0017632199999999998 3.3 0.0017633199999999999 0 0.00176324 0 0.00176334 3.3 0.00176326 3.3 0.00176336 0 0.0017632799999999999 0 0.00176338 3.3 0.0017633 3.3 0.0017634 0 0.0017633199999999999 0 0.00176342 3.3 0.00176334 3.3 0.00176344 0 0.0017633599999999998 0 0.00176346 3.3 0.00176338 3.3 0.00176348 0 0.0017633999999999998 0 0.0017634999999999999 3.3 0.00176342 3.3 0.00176352 0 0.00176344 0 0.00176354 3.3 0.00176346 3.3 0.00176356 0 0.00176348 0 0.00176358 3.3 0.0017634999999999999 3.3 0.0017636 0 0.00176352 0 0.00176362 3.3 0.0017635399999999999 3.3 0.00176364 0 0.00176356 0 0.00176366 3.3 0.0017635799999999998 3.3 0.00176368 0 0.0017636 0 0.0017637 3.3 0.0017636199999999998 3.3 0.0017637199999999999 0 0.00176364 0 0.00176374 3.3 0.00176366 3.3 0.00176376 0 0.00176368 0 0.00176378 3.3 0.0017637 3.3 0.0017638 0 0.0017637199999999999 0 0.00176382 3.3 0.00176374 3.3 0.00176384 0 0.0017637599999999999 0 0.00176386 3.3 0.00176378 3.3 0.00176388 0 0.0017637999999999998 0 0.0017638999999999999 3.3 0.00176382 3.3 0.00176392 0 0.0017638399999999998 0 0.0017639399999999999 3.3 0.00176386 3.3 0.00176396 0 0.00176388 0 0.00176398 3.3 0.0017638999999999999 3.3 0.001764 0 0.00176392 0 0.00176402 3.3 0.0017639399999999999 3.3 0.00176404 0 0.00176396 0 0.00176406 3.3 0.0017639799999999998 3.3 0.00176408 0 0.001764 0 0.0017641 3.3 0.0017640199999999998 3.3 0.0017641199999999999 0 0.00176404 0 0.00176414 3.3 0.0017640599999999998 3.3 0.0017641599999999999 0 0.00176408 0 0.00176418 3.3 0.0017641 3.3 0.0017642 0 0.0017641199999999999 0 0.00176422 3.3 0.00176414 3.3 0.00176424 0 0.0017641599999999999 0 0.00176426 3.3 0.00176418 3.3 0.00176428 0 0.0017641999999999998 0 0.0017643 3.3 0.00176422 3.3 0.00176432 0 0.0017642399999999998 0 0.0017643399999999999 3.3 0.00176426 3.3 0.00176436 0 0.00176428 0 0.00176438 3.3 0.0017643 3.3 0.0017644 0 0.00176432 0 0.00176442 3.3 0.0017643399999999999 3.3 0.00176444 0 0.00176436 0 0.00176446 3.3 0.0017643799999999999 3.3 0.00176448 0 0.0017644 0 0.0017645 3.3 0.0017644199999999998 3.3 0.0017645199999999999 0 0.00176444 0 0.00176454 3.3 0.0017644599999999998 3.3 0.0017645599999999999 0 0.00176448 0 0.00176458 3.3 0.0017645 3.3 0.0017646 0 0.0017645199999999999 0 0.00176462 3.3 0.00176454 3.3 0.00176464 0 0.0017645599999999999 0 0.00176466 3.3 0.00176458 3.3 0.00176468 0 0.0017645999999999998 0 0.0017647 3.3 0.00176462 3.3 0.00176472 0 0.0017646399999999998 0 0.0017647399999999999 3.3 0.00176466 3.3 0.00176476 0 0.0017646799999999998 0 0.0017647799999999999 3.3 0.0017647 3.3 0.0017648 0 0.00176472 0 0.00176482 3.3 0.0017647399999999999 3.3 0.00176484 0 0.00176476 0 0.00176486 3.3 0.0017647799999999999 3.3 0.00176488 0 0.0017648 0 0.0017649 3.3 0.0017648199999999998 3.3 0.00176492 0 0.00176484 0 0.00176494 3.3 0.0017648599999999998 3.3 0.0017649599999999999 0 0.00176488 0 0.00176498 3.3 0.0017648999999999998 3.3 0.0017649999999999999 0 0.00176492 0 0.00176502 3.3 0.00176494 3.3 0.00176504 0 0.0017649599999999999 0 0.00176506 3.3 0.00176498 3.3 0.00176508 0 0.0017649999999999999 0 0.0017651 3.3 0.00176502 3.3 0.00176512 0 0.0017650399999999998 0 0.00176514 3.3 0.00176506 3.3 0.00176516 0 0.0017650799999999998 0 0.0017651799999999999 3.3 0.0017651 3.3 0.0017652 0 0.00176512 0 0.00176522 3.3 0.00176514 3.3 0.00176524 0 0.00176516 0 0.00176526 3.3 0.0017651799999999999 3.3 0.00176528 0 0.0017652 0 0.0017653 3.3 0.0017652199999999999 3.3 0.00176532 0 0.00176524 0 0.00176534 3.3 0.0017652599999999998 3.3 0.0017653599999999999 0 0.00176528 0 0.00176538 3.3 0.0017652999999999998 3.3 0.0017653999999999999 0 0.00176532 0 0.00176542 3.3 0.00176534 3.3 0.00176544 0 0.0017653599999999999 0 0.00176546 3.3 0.00176538 3.3 0.00176548 0 0.0017653999999999999 0 0.0017655 3.3 0.00176542 3.3 0.00176552 0 0.0017654399999999998 0 0.00176554 3.3 0.00176546 3.3 0.00176556 0 0.0017654799999999998 0 0.0017655799999999999 3.3 0.0017655 3.3 0.0017656 0 0.0017655199999999998 0 0.0017656199999999999 3.3 0.00176554 3.3 0.00176564 0 0.00176556 0 0.00176566 3.3 0.0017655799999999999 3.3 0.00176568 0 0.0017656 0 0.0017657 3.3 0.0017656199999999999 3.3 0.00176572 0 0.00176564 0 0.00176574 3.3 0.0017656599999999998 3.3 0.00176576 0 0.00176568 0 0.00176578 3.3 0.0017656999999999998 3.3 0.0017657999999999999 0 0.00176572 0 0.00176582 3.3 0.0017657399999999998 3.3 0.0017658399999999999 0 0.00176576 0 0.00176586 3.3 0.00176578 3.3 0.00176588 0 0.0017657999999999999 0 0.0017659 3.3 0.00176582 3.3 0.00176592 0 0.0017658399999999999 0 0.00176594 3.3 0.00176586 3.3 0.00176596 0 0.0017658799999999998 0 0.00176598 3.3 0.0017659 3.3 0.001766 0 0.0017659199999999998 0 0.0017660199999999999 3.3 0.00176594 3.3 0.00176604 0 0.00176596 0 0.00176606 3.3 0.00176598 3.3 0.00176608 0 0.001766 0 0.0017661 3.3 0.0017660199999999999 3.3 0.00176612 0 0.00176604 0 0.00176614 3.3 0.0017660599999999999 3.3 0.00176616 0 0.00176608 0 0.00176618 3.3 0.0017660999999999998 3.3 0.0017661999999999999 0 0.00176612 0 0.00176622 3.3 0.0017661399999999998 3.3 0.0017662399999999999 0 0.00176616 0 0.00176626 3.3 0.00176618 3.3 0.00176628 0 0.0017661999999999999 0 0.0017663 3.3 0.00176622 3.3 0.00176632 0 0.0017662399999999999 0 0.00176634 3.3 0.00176626 3.3 0.00176636 0 0.0017662799999999998 0 0.00176638 3.3 0.0017663 3.3 0.0017664 0 0.0017663199999999998 0 0.0017664199999999999 3.3 0.00176634 3.3 0.00176644 0 0.0017663599999999998 0 0.0017664599999999999 3.3 0.00176638 3.3 0.00176648 0 0.0017664 0 0.0017665 3.3 0.0017664199999999999 3.3 0.00176652 0 0.00176644 0 0.00176654 3.3 0.0017664599999999999 3.3 0.00176656 0 0.00176648 0 0.00176658 3.3 0.0017664999999999998 3.3 0.0017666 0 0.00176652 0 0.00176662 3.3 0.0017665399999999998 3.3 0.0017666399999999999 0 0.00176656 0 0.00176666 3.3 0.0017665799999999998 3.3 0.0017666799999999999 0 0.0017666 0 0.0017667 3.3 0.00176662 3.3 0.00176672 0 0.0017666399999999999 0 0.00176674 3.3 0.00176666 3.3 0.00176676 0 0.0017666799999999999 0 0.00176678 3.3 0.0017667 3.3 0.0017668 0 0.0017667199999999998 0 0.00176682 3.3 0.00176674 3.3 0.00176684 0 0.0017667599999999998 0 0.0017668599999999999 3.3 0.00176678 3.3 0.00176688 0 0.0017668 0 0.0017669 3.3 0.00176682 3.3 0.00176692 0 0.00176684 0 0.00176694 3.3 0.0017668599999999999 3.3 0.00176696 0 0.00176688 0 0.00176698 3.3 0.0017668999999999999 3.3 0.001767 0 0.00176692 0 0.00176702 3.3 0.0017669399999999998 3.3 0.0017670399999999999 0 0.00176696 0 0.00176706 3.3 0.0017669799999999998 3.3 0.0017670799999999999 0 0.001767 0 0.0017671 3.3 0.00176702 3.3 0.00176712 0 0.0017670399999999999 0 0.00176714 3.3 0.00176706 3.3 0.00176716 0 0.0017670799999999999 0 0.00176718 3.3 0.0017671 3.3 0.0017672 0 0.0017671199999999998 0 0.00176722 3.3 0.00176714 3.3 0.00176724 0 0.0017671599999999998 0 0.0017672599999999999 3.3 0.00176718 3.3 0.00176728 0 0.0017671999999999998 0 0.0017672999999999999 3.3 0.00176722 3.3 0.00176732 0 0.00176724 0 0.00176734 3.3 0.0017672599999999999 3.3 0.00176736 0 0.00176728 0 0.00176738 3.3 0.0017672999999999999 3.3 0.0017674 0 0.00176732 0 0.00176742 3.3 0.0017673399999999998 3.3 0.00176744 0 0.00176736 0 0.00176746 3.3 0.0017673799999999998 3.3 0.0017674799999999999 0 0.0017674 0 0.0017675 3.3 0.00176742 3.3 0.00176752 0 0.00176744 0 0.00176754 3.3 0.00176746 3.3 0.00176756 0 0.0017674799999999999 0 0.00176758 3.3 0.0017675 3.3 0.0017676 0 0.0017675199999999999 0 0.00176762 3.3 0.00176754 3.3 0.00176764 0 0.0017675599999999998 0 0.0017676599999999999 3.3 0.00176758 3.3 0.00176768 0 0.0017675999999999998 0 0.0017676999999999999 3.3 0.00176762 3.3 0.00176772 0 0.00176764 0 0.00176774 3.3 0.0017676599999999999 3.3 0.00176776 0 0.00176768 0 0.00176778 3.3 0.0017676999999999999 3.3 0.0017678 0 0.00176772 0 0.00176782 3.3 0.0017677399999999998 3.3 0.00176784 0 0.00176776 0 0.00176786 3.3 0.0017677799999999998 3.3 0.0017678799999999999 0 0.0017678 0 0.0017679 3.3 0.0017678199999999998 3.3 0.0017679199999999999 0 0.00176784 0 0.00176794 3.3 0.00176786 3.3 0.00176796 0 0.0017678799999999999 0 0.00176798 3.3 0.0017679 3.3 0.001768 0 0.0017679199999999999 0 0.00176802 3.3 0.00176794 3.3 0.00176804 0 0.0017679599999999998 0 0.00176806 3.3 0.00176798 3.3 0.00176808 0 0.0017679999999999998 0 0.0017680999999999999 3.3 0.00176802 3.3 0.00176812 0 0.0017680399999999998 0 0.0017681399999999999 3.3 0.00176806 3.3 0.00176816 0 0.00176808 0 0.00176818 3.3 0.0017680999999999999 3.3 0.0017682 0 0.00176812 0 0.00176822 3.3 0.0017681399999999999 3.3 0.00176824 0 0.00176816 0 0.00176826 3.3 0.0017681799999999998 3.3 0.00176828 0 0.0017682 0 0.0017683 3.3 0.0017682199999999998 3.3 0.0017683199999999999 0 0.00176824 0 0.00176834 3.3 0.00176826 3.3 0.00176836 0 0.00176828 0 0.00176838 3.3 0.0017683 3.3 0.0017684 0 0.0017683199999999999 0 0.00176842 3.3 0.00176834 3.3 0.00176844 0 0.0017683599999999999 0 0.00176846 3.3 0.00176838 3.3 0.00176848 0 0.0017683999999999998 0 0.0017684999999999999 3.3 0.00176842 3.3 0.00176852 0 0.0017684399999999998 0 0.0017685399999999999 3.3 0.00176846 3.3 0.00176856 0 0.00176848 0 0.00176858 3.3 0.0017684999999999999 3.3 0.0017686 0 0.00176852 0 0.00176862 3.3 0.0017685399999999999 3.3 0.00176864 0 0.00176856 0 0.00176866 3.3 0.0017685799999999998 3.3 0.00176868 0 0.0017686 0 0.0017687 3.3 0.0017686199999999998 3.3 0.0017687199999999999 0 0.00176864 0 0.00176874 3.3 0.0017686599999999998 3.3 0.0017687599999999999 0 0.00176868 0 0.00176878 3.3 0.0017687 3.3 0.0017688 0 0.0017687199999999999 0 0.00176882 3.3 0.00176874 3.3 0.00176884 0 0.0017687599999999999 0 0.00176886 3.3 0.00176878 3.3 0.00176888 0 0.0017687999999999998 0 0.0017689 3.3 0.00176882 3.3 0.00176892 0 0.0017688399999999998 0 0.0017689399999999999 3.3 0.00176886 3.3 0.00176896 0 0.0017688799999999998 0 0.0017689799999999999 3.3 0.0017689 3.3 0.001769 0 0.00176892 0 0.00176902 3.3 0.0017689399999999999 3.3 0.00176904 0 0.00176896 0 0.00176906 3.3 0.0017689799999999999 3.3 0.00176908 0 0.001769 0 0.0017691 3.3 0.0017690199999999998 3.3 0.00176912 0 0.00176904 0 0.00176914 3.3 0.0017690599999999998 3.3 0.0017691599999999999 0 0.00176908 0 0.00176918 3.3 0.0017691 3.3 0.0017692 0 0.00176912 0 0.00176922 3.3 0.00176914 3.3 0.00176924 0 0.0017691599999999999 0 0.00176926 3.3 0.00176918 3.3 0.00176928 0 0.0017691999999999999 0 0.0017693 3.3 0.00176922 3.3 0.00176932 0 0.0017692399999999998 0 0.0017693399999999999 3.3 0.00176926 3.3 0.00176936 0 0.0017692799999999998 0 0.0017693799999999999 3.3 0.0017693 3.3 0.0017694 0 0.00176932 0 0.00176942 3.3 0.0017693399999999999 3.3 0.00176944 0 0.00176936 0 0.00176946 3.3 0.0017693799999999999 3.3 0.00176948 0 0.0017694 0 0.0017695 3.3 0.0017694199999999998 3.3 0.00176952 0 0.00176944 0 0.00176954 3.3 0.0017694599999999998 3.3 0.0017695599999999999 0 0.00176948 0 0.00176958 3.3 0.0017694999999999998 3.3 0.0017695999999999999 0 0.00176952 0 0.00176962 3.3 0.00176954 3.3 0.00176964 0 0.0017695599999999999 0 0.00176966 3.3 0.00176958 3.3 0.00176968 0 0.0017695999999999999 0 0.0017697 3.3 0.00176962 3.3 0.00176972 0 0.0017696399999999998 0 0.00176974 3.3 0.00176966 3.3 0.00176976 0 0.0017696799999999998 0 0.0017697799999999999 3.3 0.0017697 3.3 0.0017698 0 0.0017697199999999998 0 0.0017698199999999999 3.3 0.00176974 3.3 0.00176984 0 0.00176976 0 0.00176986 3.3 0.0017697799999999999 3.3 0.00176988 0 0.0017698 0 0.0017699 3.3 0.0017698199999999999 3.3 0.00176992 0 0.00176984 0 0.00176994 3.3 0.0017698599999999998 3.3 0.00176996 0 0.00176988 0 0.00176998 3.3 0.0017698999999999998 3.3 0.0017699999999999999 0 0.00176992 0 0.00177002 3.3 0.00176994 3.3 0.00177004 0 0.00176996 0 0.00177006 3.3 0.00176998 3.3 0.00177008 0 0.0017699999999999999 0 0.0017701 3.3 0.00177002 3.3 0.00177012 0 0.0017700399999999999 0 0.00177014 3.3 0.00177006 3.3 0.00177016 0 0.0017700799999999998 0 0.0017701799999999999 3.3 0.0017701 3.3 0.0017702 0 0.0017701199999999998 0 0.0017702199999999999 3.3 0.00177014 3.3 0.00177024 0 0.00177016 0 0.00177026 3.3 0.0017701799999999999 3.3 0.00177028 0 0.0017702 0 0.0017703 3.3 0.0017702199999999999 3.3 0.00177032 0 0.00177024 0 0.00177034 3.3 0.0017702599999999998 3.3 0.00177036 0 0.00177028 0 0.00177038 3.3 0.0017702999999999998 3.3 0.0017703999999999999 0 0.00177032 0 0.00177042 3.3 0.0017703399999999998 3.3 0.0017704399999999999 0 0.00177036 0 0.00177046 3.3 0.00177038 3.3 0.00177048 0 0.0017703999999999999 0 0.0017705 3.3 0.00177042 3.3 0.00177052 0 0.0017704399999999999 0 0.00177054 3.3 0.00177046 3.3 0.00177056 0 0.0017704799999999998 0 0.00177058 3.3 0.0017705 3.3 0.0017706 0 0.0017705199999999998 0 0.0017706199999999999 3.3 0.00177054 3.3 0.00177064 0 0.00177056 0 0.00177066 3.3 0.00177058 3.3 0.00177068 0 0.0017706 0 0.0017707 3.3 0.0017706199999999999 3.3 0.00177072 0 0.00177064 0 0.00177074 3.3 0.0017706599999999999 3.3 0.00177076 0 0.00177068 0 0.00177078 3.3 0.0017706999999999998 3.3 0.0017707999999999999 0 0.00177072 0 0.00177082 3.3 0.0017707399999999998 3.3 0.0017708399999999999 0 0.00177076 0 0.00177086 3.3 0.00177078 3.3 0.00177088 0 0.0017707999999999999 0 0.0017709 3.3 0.00177082 3.3 0.00177092 0 0.0017708399999999999 0 0.00177094 3.3 0.00177086 3.3 0.00177096 0 0.0017708799999999999 0 0.00177098 3.3 0.0017709 3.3 0.001771 0 0.0017709199999999998 0 0.0017710199999999999 3.3 0.00177094 3.3 0.00177104 0 0.0017709599999999998 0 0.0017710599999999999 3.3 0.00177098 3.3 0.00177108 0 0.001771 0 0.0017711 3.3 0.0017710199999999999 3.3 0.00177112 0 0.00177104 0 0.00177114 3.3 0.0017710599999999999 3.3 0.00177116 0 0.00177108 0 0.00177118 3.3 0.0017710999999999998 3.3 0.0017712 0 0.00177112 0 0.00177122 3.3 0.0017711399999999998 3.3 0.0017712399999999999 0 0.00177116 0 0.00177126 3.3 0.0017711799999999998 3.3 0.0017712799999999999 0 0.0017712 0 0.0017713 3.3 0.00177122 3.3 0.00177132 0 0.0017712399999999999 0 0.00177134 3.3 0.00177126 3.3 0.00177136 0 0.0017712799999999999 0 0.00177138 3.3 0.0017713 3.3 0.0017714 0 0.0017713199999999998 0 0.00177142 3.3 0.00177134 3.3 0.00177144 0 0.0017713599999999998 0 0.0017714599999999999 3.3 0.00177138 3.3 0.00177148 0 0.0017714 0 0.0017715 3.3 0.00177142 3.3 0.00177152 0 0.00177144 0 0.00177154 3.3 0.0017714599999999999 3.3 0.00177156 0 0.00177148 0 0.00177158 3.3 0.0017714999999999999 3.3 0.0017716 0 0.00177152 0 0.00177162 3.3 0.0017715399999999998 3.3 0.0017716399999999999 0 0.00177156 0 0.00177166 3.3 0.0017715799999999998 3.3 0.0017716799999999999 0 0.0017716 0 0.0017717 3.3 0.00177162 3.3 0.00177172 0 0.0017716399999999999 0 0.00177174 3.3 0.00177166 3.3 0.00177176 0 0.0017716799999999999 0 0.00177178 3.3 0.0017717 3.3 0.0017718 0 0.0017717199999999998 0 0.00177182 3.3 0.00177174 3.3 0.00177184 0 0.0017717599999999998 0 0.0017718599999999999 3.3 0.00177178 3.3 0.00177188 0 0.0017717999999999998 0 0.0017718999999999999 3.3 0.00177182 3.3 0.00177192 0 0.00177184 0 0.00177194 3.3 0.0017718599999999999 3.3 0.00177196 0 0.00177188 0 0.00177198 3.3 0.0017718999999999999 3.3 0.001772 0 0.00177192 0 0.00177202 3.3 0.0017719399999999998 3.3 0.00177204 0 0.00177196 0 0.00177206 3.3 0.0017719799999999998 3.3 0.0017720799999999999 0 0.001772 0 0.0017721 3.3 0.0017720199999999998 3.3 0.0017721199999999999 0 0.00177204 0 0.00177214 3.3 0.00177206 3.3 0.00177216 0 0.0017720799999999999 0 0.00177218 3.3 0.0017721 3.3 0.0017722 0 0.0017721199999999999 0 0.00177222 3.3 0.00177214 3.3 0.00177224 0 0.0017721599999999998 0 0.00177226 3.3 0.00177218 3.3 0.00177228 0 0.0017721999999999998 0 0.0017722999999999999 3.3 0.00177222 3.3 0.00177232 0 0.00177224 0 0.00177234 3.3 0.00177226 3.3 0.00177236 0 0.00177228 0 0.00177238 3.3 0.0017722999999999999 3.3 0.0017724 0 0.00177232 0 0.00177242 3.3 0.0017723399999999999 3.3 0.00177244 0 0.00177236 0 0.00177246 3.3 0.0017723799999999998 3.3 0.0017724799999999999 0 0.0017724 0 0.0017725 3.3 0.0017724199999999998 3.3 0.0017725199999999999 0 0.00177244 0 0.00177254 3.3 0.00177246 3.3 0.00177256 0 0.0017724799999999999 0 0.00177258 3.3 0.0017725 3.3 0.0017726 0 0.0017725199999999999 0 0.00177262 3.3 0.00177254 3.3 0.00177264 0 0.0017725599999999998 0 0.00177266 3.3 0.00177258 3.3 0.00177268 0 0.0017725999999999998 0 0.0017726999999999999 3.3 0.00177262 3.3 0.00177272 0 0.0017726399999999998 0 0.0017727399999999999 3.3 0.00177266 3.3 0.00177276 0 0.00177268 0 0.00177278 3.3 0.0017726999999999999 3.3 0.0017728 0 0.00177272 0 0.00177282 3.3 0.0017727399999999999 3.3 0.00177284 0 0.00177276 0 0.00177286 3.3 0.0017727799999999998 3.3 0.00177288 0 0.0017728 0 0.0017729 3.3 0.0017728199999999998 3.3 0.0017729199999999999 0 0.00177284 0 0.00177294 3.3 0.0017728599999999998 3.3 0.0017729599999999999 0 0.00177288 0 0.00177298 3.3 0.0017729 3.3 0.001773 0 0.0017729199999999999 0 0.00177302 3.3 0.00177294 3.3 0.00177304 0 0.0017729599999999999 0 0.00177306 3.3 0.00177298 3.3 0.00177308 0 0.0017729999999999998 0 0.0017731 3.3 0.00177302 3.3 0.00177312 0 0.0017730399999999998 0 0.0017731399999999999 3.3 0.00177306 3.3 0.00177316 0 0.00177308 0 0.00177318 3.3 0.0017731 3.3 0.0017732 0 0.00177312 0 0.00177322 3.3 0.0017731399999999999 3.3 0.00177324 0 0.00177316 0 0.00177326 3.3 0.0017731799999999999 3.3 0.00177328 0 0.0017732 0 0.0017733 3.3 0.0017732199999999998 3.3 0.0017733199999999999 0 0.00177324 0 0.00177334 3.3 0.0017732599999999998 3.3 0.0017733599999999999 0 0.00177328 0 0.00177338 3.3 0.0017733 3.3 0.0017734 0 0.0017733199999999999 0 0.00177342 3.3 0.00177334 3.3 0.00177344 0 0.0017733599999999999 0 0.00177346 3.3 0.00177338 3.3 0.00177348 0 0.0017733999999999998 0 0.0017735 3.3 0.00177342 3.3 0.00177352 0 0.0017734399999999998 0 0.0017735399999999999 3.3 0.00177346 3.3 0.00177356 0 0.0017734799999999998 0 0.0017735799999999999 3.3 0.0017735 3.3 0.0017736 0 0.00177352 0 0.00177362 3.3 0.0017735399999999999 3.3 0.00177364 0 0.00177356 0 0.00177366 3.3 0.0017735799999999999 3.3 0.00177368 0 0.0017736 0 0.0017737 3.3 0.0017736199999999998 3.3 0.00177372 0 0.00177364 0 0.00177374 3.3 0.0017736599999999998 3.3 0.0017737599999999999 0 0.00177368 0 0.00177378 3.3 0.0017736999999999998 3.3 0.0017737999999999999 0 0.00177372 0 0.00177382 3.3 0.00177374 3.3 0.00177384 0 0.0017737599999999999 0 0.00177386 3.3 0.00177378 3.3 0.00177388 0 0.0017737999999999999 0 0.0017739 3.3 0.00177382 3.3 0.00177392 0 0.0017738399999999998 0 0.00177394 3.3 0.00177386 3.3 0.00177396 0 0.0017738799999999998 0 0.0017739799999999999 3.3 0.0017739 3.3 0.001774 0 0.00177392 0 0.00177402 3.3 0.00177394 3.3 0.00177404 0 0.00177396 0 0.00177406 3.3 0.0017739799999999999 3.3 0.00177408 0 0.001774 0 0.0017741 3.3 0.0017740199999999999 3.3 0.00177412 0 0.00177404 0 0.00177414 3.3 0.0017740599999999998 3.3 0.0017741599999999999 0 0.00177408 0 0.00177418 3.3 0.0017740999999999998 3.3 0.0017741999999999999 0 0.00177412 0 0.00177422 3.3 0.00177414 3.3 0.00177424 0 0.0017741599999999999 0 0.00177426 3.3 0.00177418 3.3 0.00177428 0 0.0017741999999999999 0 0.0017743 3.3 0.00177422 3.3 0.00177432 0 0.0017742399999999998 0 0.00177434 3.3 0.00177426 3.3 0.00177436 0 0.0017742799999999998 0 0.0017743799999999999 3.3 0.0017743 3.3 0.0017744 0 0.0017743199999999998 0 0.0017744199999999999 3.3 0.00177434 3.3 0.00177444 0 0.00177436 0 0.00177446 3.3 0.0017743799999999999 3.3 0.00177448 0 0.0017744 0 0.0017745 3.3 0.0017744199999999999 3.3 0.00177452 0 0.00177444 0 0.00177454 3.3 0.0017744599999999998 3.3 0.00177456 0 0.00177448 0 0.00177458 3.3 0.0017744999999999998 3.3 0.0017745999999999999 0 0.00177452 0 0.00177462 3.3 0.00177454 3.3 0.00177464 0 0.00177456 0 0.00177466 3.3 0.00177458 3.3 0.00177468 0 0.0017745999999999999 0 0.0017747 3.3 0.00177462 3.3 0.00177472 0 0.0017746399999999999 0 0.00177474 3.3 0.00177466 3.3 0.00177476 0 0.0017746799999999998 0 0.0017747799999999999 3.3 0.0017747 3.3 0.0017748 0 0.0017747199999999998 0 0.0017748199999999999 3.3 0.00177474 3.3 0.00177484 0 0.00177476 0 0.00177486 3.3 0.0017747799999999999 3.3 0.00177488 0 0.0017748 0 0.0017749 3.3 0.0017748199999999999 3.3 0.00177492 0 0.00177484 0 0.00177494 3.3 0.0017748599999999998 3.3 0.00177496 0 0.00177488 0 0.00177498 3.3 0.0017748999999999998 3.3 0.0017749999999999999 0 0.00177492 0 0.00177502 3.3 0.0017749399999999998 3.3 0.0017750399999999999 0 0.00177496 0 0.00177506 3.3 0.00177498 3.3 0.00177508 0 0.0017749999999999999 0 0.0017751 3.3 0.00177502 3.3 0.00177512 0 0.0017750399999999999 0 0.00177514 3.3 0.00177506 3.3 0.00177516 0 0.0017750799999999998 0 0.00177518 3.3 0.0017751 3.3 0.0017752 0 0.0017751199999999998 0 0.0017752199999999999 3.3 0.00177514 3.3 0.00177524 0 0.0017751599999999998 0 0.0017752599999999999 3.3 0.00177518 3.3 0.00177528 0 0.0017752 0 0.0017753 3.3 0.0017752199999999999 3.3 0.00177532 0 0.00177524 0 0.00177534 3.3 0.0017752599999999999 3.3 0.00177536 0 0.00177528 0 0.00177538 3.3 0.0017752999999999998 3.3 0.0017754 0 0.00177532 0 0.00177542 3.3 0.0017753399999999998 3.3 0.0017754399999999999 0 0.00177536 0 0.00177546 3.3 0.00177538 3.3 0.00177548 0 0.0017754 0 0.0017755 3.3 0.00177542 3.3 0.00177552 0 0.0017754399999999999 0 0.00177554 3.3 0.00177546 3.3 0.00177556 0 0.0017754799999999999 0 0.00177558 3.3 0.0017755 3.3 0.0017756 0 0.0017755199999999998 0 0.0017756199999999999 3.3 0.00177554 3.3 0.00177564 0 0.0017755599999999998 0 0.0017756599999999999 3.3 0.00177558 3.3 0.00177568 0 0.0017756 0 0.0017757 3.3 0.0017756199999999999 3.3 0.00177572 0 0.00177564 0 0.00177574 3.3 0.0017756599999999999 3.3 0.00177576 0 0.00177568 0 0.00177578 3.3 0.0017756999999999998 3.3 0.0017758 0 0.00177572 0 0.00177582 3.3 0.0017757399999999998 3.3 0.0017758399999999999 0 0.00177576 0 0.00177586 3.3 0.0017757799999999998 3.3 0.0017758799999999999 0 0.0017758 0 0.0017759 3.3 0.00177582 3.3 0.00177592 0 0.0017758399999999999 0 0.00177594 3.3 0.00177586 3.3 0.00177596 0 0.0017758799999999999 0 0.00177598 3.3 0.0017759 3.3 0.001776 0 0.0017759199999999998 0 0.00177602 3.3 0.00177594 3.3 0.00177604 0 0.0017759599999999998 0 0.0017760599999999999 3.3 0.00177598 3.3 0.00177608 0 0.0017759999999999998 0 0.0017760999999999999 3.3 0.00177602 3.3 0.00177612 0 0.00177604 0 0.00177614 3.3 0.0017760599999999999 3.3 0.00177616 0 0.00177608 0 0.00177618 3.3 0.0017760999999999999 3.3 0.0017762 0 0.00177612 0 0.00177622 3.3 0.0017761399999999998 3.3 0.00177624 0 0.00177616 0 0.00177626 3.3 0.0017761799999999998 3.3 0.0017762799999999999 0 0.0017762 0 0.0017763 3.3 0.00177622 3.3 0.00177632 0 0.00177624 0 0.00177634 3.3 0.00177626 3.3 0.00177636 0 0.0017762799999999999 0 0.00177638 3.3 0.0017763 3.3 0.0017764 0 0.0017763199999999999 0 0.00177642 3.3 0.00177634 3.3 0.00177644 0 0.0017763599999999998 0 0.0017764599999999999 3.3 0.00177638 3.3 0.00177648 0 0.0017763999999999998 0 0.0017764999999999999 3.3 0.00177642 3.3 0.00177652 0 0.00177644 0 0.00177654 3.3 0.0017764599999999999 3.3 0.00177656 0 0.00177648 0 0.00177658 3.3 0.0017764999999999999 3.3 0.0017766 0 0.00177652 0 0.00177662 3.3 0.0017765399999999998 3.3 0.00177664 0 0.00177656 0 0.00177666 3.3 0.0017765799999999998 3.3 0.0017766799999999999 0 0.0017766 0 0.0017767 3.3 0.0017766199999999998 3.3 0.0017767199999999999 0 0.00177664 0 0.00177674 3.3 0.00177666 3.3 0.00177676 0 0.0017766799999999999 0 0.00177678 3.3 0.0017767 3.3 0.0017768 0 0.0017767199999999999 0 0.00177682 3.3 0.00177674 3.3 0.00177684 0 0.0017767599999999998 0 0.00177686 3.3 0.00177678 3.3 0.00177688 0 0.0017767999999999998 0 0.0017768999999999999 3.3 0.00177682 3.3 0.00177692 0 0.0017768399999999998 0 0.0017769399999999999 3.3 0.00177686 3.3 0.00177696 0 0.00177688 0 0.00177698 3.3 0.0017768999999999999 3.3 0.001777 0 0.00177692 0 0.00177702 3.3 0.0017769399999999999 3.3 0.00177704 0 0.00177696 0 0.00177706 3.3 0.0017769799999999998 3.3 0.00177708 0 0.001777 0 0.0017771 3.3 0.0017770199999999998 3.3 0.0017771199999999999 0 0.00177704 0 0.00177714 3.3 0.00177706 3.3 0.00177716 0 0.00177708 0 0.00177718 3.3 0.0017771 3.3 0.0017772 0 0.0017771199999999999 0 0.00177722 3.3 0.00177714 3.3 0.00177724 0 0.0017771599999999999 0 0.00177726 3.3 0.00177718 3.3 0.00177728 0 0.0017771999999999998 0 0.0017772999999999999 3.3 0.00177722 3.3 0.00177732 0 0.0017772399999999998 0 0.0017773399999999999 3.3 0.00177726 3.3 0.00177736 0 0.00177728 0 0.00177738 3.3 0.0017772999999999999 3.3 0.0017774 0 0.00177732 0 0.00177742 3.3 0.0017773399999999999 3.3 0.00177744 0 0.00177736 0 0.00177746 3.3 0.0017773799999999998 3.3 0.00177748 0 0.0017774 0 0.0017775 3.3 0.0017774199999999998 3.3 0.0017775199999999999 0 0.00177744 0 0.00177754 3.3 0.0017774599999999998 3.3 0.0017775599999999999 0 0.00177748 0 0.00177758 3.3 0.0017775 3.3 0.0017776 0 0.0017775199999999999 0 0.00177762 3.3 0.00177754 3.3 0.00177764 0 0.0017775599999999999 0 0.00177766 3.3 0.00177758 3.3 0.00177768 0 0.0017775999999999998 0 0.0017777 3.3 0.00177762 3.3 0.00177772 0 0.0017776399999999998 0 0.0017777399999999999 3.3 0.00177766 3.3 0.00177776 0 0.00177768 0 0.00177778 3.3 0.0017777 3.3 0.0017778 0 0.00177772 0 0.00177782 3.3 0.0017777399999999999 3.3 0.00177784 0 0.00177776 0 0.00177786 3.3 0.0017777799999999999 3.3 0.00177788 0 0.0017778 0 0.0017779 3.3 0.0017778199999999998 3.3 0.0017779199999999999 0 0.00177784 0 0.00177794 3.3 0.0017778599999999998 3.3 0.0017779599999999999 0 0.00177788 0 0.00177798 3.3 0.0017779 3.3 0.001778 0 0.0017779199999999999 0 0.00177802 3.3 0.00177794 3.3 0.00177804 0 0.0017779599999999999 0 0.00177806 3.3 0.00177798 3.3 0.00177808 0 0.0017779999999999998 0 0.0017781 3.3 0.00177802 3.3 0.00177812 0 0.0017780399999999998 0 0.0017781399999999999 3.3 0.00177806 3.3 0.00177816 0 0.0017780799999999998 0 0.0017781799999999999 3.3 0.0017781 3.3 0.0017782 0 0.00177812 0 0.00177822 3.3 0.0017781399999999999 3.3 0.00177824 0 0.00177816 0 0.00177826 3.3 0.0017781799999999999 3.3 0.00177828 0 0.0017782 0 0.0017783 3.3 0.0017782199999999998 3.3 0.00177832 0 0.00177824 0 0.00177834 3.3 0.0017782599999999998 3.3 0.0017783599999999999 0 0.00177828 0 0.00177838 3.3 0.0017782999999999998 3.3 0.0017783999999999999 0 0.00177832 0 0.00177842 3.3 0.00177834 3.3 0.00177844 0 0.0017783599999999999 0 0.00177846 3.3 0.00177838 3.3 0.00177848 0 0.0017783999999999999 0 0.0017785 3.3 0.00177842 3.3 0.00177852 0 0.0017784399999999998 0 0.00177854 3.3 0.00177846 3.3 0.00177856 0 0.0017784799999999998 0 0.0017785799999999999 3.3 0.0017785 3.3 0.0017786 0 0.00177852 0 0.00177862 3.3 0.00177854 3.3 0.00177864 0 0.00177856 0 0.00177866 3.3 0.0017785799999999999 3.3 0.00177868 0 0.0017786 0 0.0017787 3.3 0.0017786199999999999 3.3 0.00177872 0 0.00177864 0 0.00177874 3.3 0.0017786599999999998 3.3 0.0017787599999999999 0 0.00177868 0 0.00177878 3.3 0.0017786999999999998 3.3 0.0017787999999999999 0 0.00177872 0 0.00177882 3.3 0.00177874 3.3 0.00177884 0 0.0017787599999999999 0 0.00177886 3.3 0.00177878 3.3 0.00177888 0 0.0017787999999999999 0 0.0017789 3.3 0.00177882 3.3 0.00177892 0 0.0017788399999999998 0 0.00177894 3.3 0.00177886 3.3 0.00177896 0 0.0017788799999999998 0 0.0017789799999999999 3.3 0.0017789 3.3 0.001779 0 0.0017789199999999998 0 0.0017790199999999999 3.3 0.00177894 3.3 0.00177904 0 0.00177896 0 0.00177906 3.3 0.0017789799999999999 3.3 0.00177908 0 0.001779 0 0.0017791 3.3 0.0017790199999999999 3.3 0.00177912 0 0.00177904 0 0.00177914 3.3 0.0017790599999999998 3.3 0.00177916 0 0.00177908 0 0.00177918 3.3 0.0017790999999999998 3.3 0.0017791999999999999 0 0.00177912 0 0.00177922 3.3 0.0017791399999999998 3.3 0.0017792399999999999 0 0.00177916 0 0.00177926 3.3 0.00177918 3.3 0.00177928 0 0.0017791999999999999 0 0.0017793 3.3 0.00177922 3.3 0.00177932 0 0.0017792399999999999 0 0.00177934 3.3 0.00177926 3.3 0.00177936 0 0.0017792799999999998 0 0.00177938 3.3 0.0017793 3.3 0.0017794 0 0.0017793199999999998 0 0.0017794199999999999 3.3 0.00177934 3.3 0.00177944 0 0.00177936 0 0.00177946 3.3 0.00177938 3.3 0.00177948 0 0.0017794 0 0.0017795 3.3 0.0017794199999999999 3.3 0.00177952 0 0.00177944 0 0.00177954 3.3 0.0017794599999999999 3.3 0.00177956 0 0.00177948 0 0.00177958 3.3 0.0017794999999999998 3.3 0.0017795999999999999 0 0.00177952 0 0.00177962 3.3 0.0017795399999999998 3.3 0.0017796399999999999 0 0.00177956 0 0.00177966 3.3 0.00177958 3.3 0.00177968 0 0.0017795999999999999 0 0.0017797 3.3 0.00177962 3.3 0.00177972 0 0.0017796399999999999 0 0.00177974 3.3 0.00177966 3.3 0.00177976 0 0.0017796799999999998 0 0.00177978 3.3 0.0017797 3.3 0.0017798 0 0.0017797199999999998 0 0.0017798199999999999 3.3 0.00177974 3.3 0.00177984 0 0.0017797599999999998 0 0.0017798599999999999 3.3 0.00177978 3.3 0.00177988 0 0.0017798 0 0.0017799 3.3 0.0017798199999999999 3.3 0.00177992 0 0.00177984 0 0.00177994 3.3 0.0017798599999999999 3.3 0.00177996 0 0.00177988 0 0.00177998 3.3 0.0017798999999999998 3.3 0.00178 0 0.00177992 0 0.00178002 3.3 0.0017799399999999998 3.3 0.0017800399999999999 0 0.00177996 0 0.00178006 3.3 0.0017799799999999998 3.3 0.0017800799999999999 0 0.00178 0 0.0017801 3.3 0.00178002 3.3 0.00178012 0 0.0017800399999999999 0 0.00178014 3.3 0.00178006 3.3 0.00178016 0 0.0017800799999999999 0 0.00178018 3.3 0.0017801 3.3 0.0017802 0 0.0017801199999999998 0 0.00178022 3.3 0.00178014 3.3 0.00178024 0 0.0017801599999999998 0 0.0017802599999999999 3.3 0.00178018 3.3 0.00178028 0 0.0017802 0 0.0017803 3.3 0.00178022 3.3 0.00178032 0 0.00178024 0 0.00178034 3.3 0.0017802599999999999 3.3 0.00178036 0 0.00178028 0 0.00178038 3.3 0.0017802999999999999 3.3 0.0017804 0 0.00178032 0 0.00178042 3.3 0.0017803399999999998 3.3 0.0017804399999999999 0 0.00178036 0 0.00178046 3.3 0.0017803799999999998 3.3 0.0017804799999999999 0 0.0017804 0 0.0017805 3.3 0.00178042 3.3 0.00178052 0 0.0017804399999999999 0 0.00178054 3.3 0.00178046 3.3 0.00178056 0 0.0017804799999999999 0 0.00178058 3.3 0.0017805 3.3 0.0017806 0 0.0017805199999999998 0 0.00178062 3.3 0.00178054 3.3 0.00178064 0 0.0017805599999999998 0 0.0017806599999999999 3.3 0.00178058 3.3 0.00178068 0 0.0017805999999999998 0 0.0017806999999999999 3.3 0.00178062 3.3 0.00178072 0 0.00178064 0 0.00178074 3.3 0.0017806599999999999 3.3 0.00178076 0 0.00178068 0 0.00178078 3.3 0.0017806999999999999 3.3 0.0017808 0 0.00178072 0 0.00178082 3.3 0.0017807399999999998 3.3 0.00178084 0 0.00178076 0 0.00178086 3.3 0.0017807799999999998 3.3 0.0017808799999999999 0 0.0017808 0 0.0017809 3.3 0.00178082 3.3 0.00178092 0 0.00178084 0 0.00178094 3.3 0.00178086 3.3 0.00178096 0 0.0017808799999999999 0 0.00178098 3.3 0.0017809 3.3 0.001781 0 0.0017809199999999999 0 0.00178102 3.3 0.00178094 3.3 0.00178104 0 0.0017809599999999998 0 0.0017810599999999999 3.3 0.00178098 3.3 0.00178108 0 0.0017809999999999998 0 0.0017810999999999999 3.3 0.00178102 3.3 0.00178112 0 0.00178104 0 0.00178114 3.3 0.0017810599999999999 3.3 0.00178116 0 0.00178108 0 0.00178118 3.3 0.0017810999999999999 3.3 0.0017812 0 0.00178112 0 0.00178122 3.3 0.0017811399999999999 3.3 0.00178124 0 0.00178116 0 0.00178126 3.3 0.0017811799999999998 3.3 0.0017812799999999999 0 0.0017812 0 0.0017813 3.3 0.0017812199999999998 3.3 0.0017813199999999999 0 0.00178124 0 0.00178134 3.3 0.00178126 3.3 0.00178136 0 0.0017812799999999999 0 0.00178138 3.3 0.0017813 3.3 0.0017814 0 0.0017813199999999999 0 0.00178142 3.3 0.00178134 3.3 0.00178144 0 0.0017813599999999998 0 0.00178146 3.3 0.00178138 3.3 0.00178148 0 0.0017813999999999998 0 0.0017814999999999999 3.3 0.00178142 3.3 0.00178152 0 0.0017814399999999998 0 0.0017815399999999999 3.3 0.00178146 3.3 0.00178156 0 0.00178148 0 0.00178158 3.3 0.0017814999999999999 3.3 0.0017816 0 0.00178152 0 0.00178162 3.3 0.0017815399999999999 3.3 0.00178164 0 0.00178156 0 0.00178166 3.3 0.0017815799999999998 3.3 0.00178168 0 0.0017816 0 0.0017817 3.3 0.0017816199999999998 3.3 0.0017817199999999999 0 0.00178164 0 0.00178174 3.3 0.00178166 3.3 0.00178176 0 0.00178168 0 0.00178178 3.3 0.0017817 3.3 0.0017818 0 0.0017817199999999999 0 0.00178182 3.3 0.00178174 3.3 0.00178184 0 0.0017817599999999999 0 0.00178186 3.3 0.00178178 3.3 0.00178188 0 0.0017817999999999998 0 0.0017818999999999999 3.3 0.00178182 3.3 0.00178192 0 0.0017818399999999998 0 0.0017819399999999999 3.3 0.00178186 3.3 0.00178196 0 0.00178188 0 0.00178198 3.3 0.0017818999999999999 3.3 0.001782 0 0.00178192 0 0.00178202 3.3 0.0017819399999999999 3.3 0.00178204 0 0.00178196 0 0.00178206 3.3 0.0017819799999999998 3.3 0.00178208 0 0.001782 0 0.0017821 3.3 0.0017820199999999998 3.3 0.0017821199999999999 0 0.00178204 0 0.00178214 3.3 0.0017820599999999998 3.3 0.0017821599999999999 0 0.00178208 0 0.00178218 3.3 0.0017821 3.3 0.0017822 0 0.0017821199999999999 0 0.00178222 3.3 0.00178214 3.3 0.00178224 0 0.0017821599999999999 0 0.00178226 3.3 0.00178218 3.3 0.00178228 0 0.0017821999999999998 0 0.0017823 3.3 0.00178222 3.3 0.00178232 0 0.0017822399999999998 0 0.0017823399999999999 3.3 0.00178226 3.3 0.00178236 0 0.0017822799999999998 0 0.0017823799999999999 3.3 0.0017823 3.3 0.0017824 0 0.00178232 0 0.00178242 3.3 0.0017823399999999999 3.3 0.00178244 0 0.00178236 0 0.00178246 3.3 0.0017823799999999999 3.3 0.00178248 0 0.0017824 0 0.0017825 3.3 0.0017824199999999998 3.3 0.00178252 0 0.00178244 0 0.00178254 3.3 0.0017824599999999998 3.3 0.0017825599999999999 0 0.00178248 0 0.00178258 3.3 0.0017825 3.3 0.0017826 0 0.00178252 0 0.00178262 3.3 0.00178254 3.3 0.00178264 0 0.0017825599999999999 0 0.00178266 3.3 0.00178258 3.3 0.00178268 0 0.0017825999999999999 0 0.0017827 3.3 0.00178262 3.3 0.00178272 0 0.0017826399999999998 0 0.0017827399999999999 3.3 0.00178266 3.3 0.00178276 0 0.0017826799999999998 0 0.0017827799999999999 3.3 0.0017827 3.3 0.0017828 0 0.00178272 0 0.00178282 3.3 0.0017827399999999999 3.3 0.00178284 0 0.00178276 0 0.00178286 3.3 0.0017827799999999999 3.3 0.00178288 0 0.0017828 0 0.0017829 3.3 0.0017828199999999998 3.3 0.00178292 0 0.00178284 0 0.00178294 3.3 0.0017828599999999998 3.3 0.0017829599999999999 0 0.00178288 0 0.00178298 3.3 0.0017828999999999998 3.3 0.0017829999999999999 0 0.00178292 0 0.00178302 3.3 0.00178294 3.3 0.00178304 0 0.0017829599999999999 0 0.00178306 3.3 0.00178298 3.3 0.00178308 0 0.0017829999999999999 0 0.0017831 3.3 0.00178302 3.3 0.00178312 0 0.0017830399999999998 0 0.00178314 3.3 0.00178306 3.3 0.00178316 0 0.0017830799999999998 0 0.0017831799999999999 3.3 0.0017831 3.3 0.0017832 0 0.0017831199999999998 0 0.0017832199999999999 3.3 0.00178314 3.3 0.00178324 0 0.00178316 0 0.00178326 3.3 0.0017831799999999999 3.3 0.00178328 0 0.0017832 0 0.0017833 3.3 0.0017832199999999999 3.3 0.00178332 0 0.00178324 0 0.00178334 3.3 0.0017832599999999998 3.3 0.00178336 0 0.00178328 0 0.00178338 3.3 0.0017832999999999998 3.3 0.0017833999999999999 0 0.00178332 0 0.00178342 3.3 0.00178334 3.3 0.00178344 0 0.00178336 0 0.00178346 3.3 0.00178338 3.3 0.00178348 0 0.0017833999999999999 0 0.0017835 3.3 0.00178342 3.3 0.00178352 0 0.0017834399999999999 0 0.00178354 3.3 0.00178346 3.3 0.00178356 0 0.0017834799999999998 0 0.0017835799999999999 3.3 0.0017835 3.3 0.0017836 0 0.0017835199999999998 0 0.0017836199999999999 3.3 0.00178354 3.3 0.00178364 0 0.00178356 0 0.00178366 3.3 0.0017835799999999999 3.3 0.00178368 0 0.0017836 0 0.0017837 3.3 0.0017836199999999999 3.3 0.00178372 0 0.00178364 0 0.00178374 3.3 0.0017836599999999998 3.3 0.00178376 0 0.00178368 0 0.00178378 3.3 0.0017836999999999998 3.3 0.0017837999999999999 0 0.00178372 0 0.00178382 3.3 0.0017837399999999998 3.3 0.0017838399999999999 0 0.00178376 0 0.00178386 3.3 0.00178378 3.3 0.00178388 0 0.0017837999999999999 0 0.0017839 3.3 0.00178382 3.3 0.00178392 0 0.0017838399999999999 0 0.00178394 3.3 0.00178386 3.3 0.00178396 0 0.0017838799999999998 0 0.00178398 3.3 0.0017839 3.3 0.001784 0 0.0017839199999999998 0 0.0017840199999999999 3.3 0.00178394 3.3 0.00178404 0 0.0017839599999999998 0 0.0017840599999999999 3.3 0.00178398 3.3 0.00178408 0 0.001784 0 0.0017841 3.3 0.0017840199999999999 3.3 0.00178412 0 0.00178404 0 0.00178414 3.3 0.0017840599999999999 3.3 0.00178416 0 0.00178408 0 0.00178418 3.3 0.0017840999999999998 3.3 0.0017842 0 0.00178412 0 0.00178422 3.3 0.0017841399999999998 3.3 0.0017842399999999999 0 0.00178416 0 0.00178426 3.3 0.00178418 3.3 0.00178428 0 0.0017842 0 0.0017843 3.3 0.00178422 3.3 0.00178432 0 0.0017842399999999999 0 0.00178434 3.3 0.00178426 3.3 0.00178436 0 0.0017842799999999999 0 0.00178438 3.3 0.0017843 3.3 0.0017844 0 0.0017843199999999998 0 0.0017844199999999999 3.3 0.00178434 3.3 0.00178444 0 0.0017843599999999998 0 0.0017844599999999999 3.3 0.00178438 3.3 0.00178448 0 0.0017844 0 0.0017845 3.3 0.0017844199999999999 3.3 0.00178452 0 0.00178444 0 0.00178454 3.3 0.0017844599999999999 3.3 0.00178456 0 0.00178448 0 0.00178458 3.3 0.0017844999999999998 3.3 0.0017846 0 0.00178452 0 0.00178462 3.3 0.0017845399999999998 3.3 0.0017846399999999999 0 0.00178456 0 0.00178466 3.3 0.0017845799999999998 3.3 0.0017846799999999999 0 0.0017846 0 0.0017847 3.3 0.00178462 3.3 0.00178472 0 0.0017846399999999999 0 0.00178474 3.3 0.00178466 3.3 0.00178476 0 0.0017846799999999999 0 0.00178478 3.3 0.0017847 3.3 0.0017848 0 0.0017847199999999998 0 0.00178482 3.3 0.00178474 3.3 0.00178484 0 0.0017847599999999998 0 0.0017848599999999999 3.3 0.00178478 3.3 0.00178488 0 0.0017848 0 0.0017849 3.3 0.00178482 3.3 0.00178492 0 0.00178484 0 0.00178494 3.3 0.0017848599999999999 3.3 0.00178496 0 0.00178488 0 0.00178498 3.3 0.0017848999999999999 3.3 0.001785 0 0.00178492 0 0.00178502 3.3 0.0017849399999999998 3.3 0.0017850399999999999 0 0.00178496 0 0.00178506 3.3 0.0017849799999999998 3.3 0.0017850799999999999 0 0.001785 0 0.0017851 3.3 0.00178502 3.3 0.00178512 0 0.0017850399999999999 0 0.00178514 3.3 0.00178506 3.3 0.00178516 0 0.0017850799999999999 0 0.00178518 3.3 0.0017851 3.3 0.0017852 0 0.0017851199999999998 0 0.00178522 3.3 0.00178514 3.3 0.00178524 0 0.0017851599999999998 0 0.0017852599999999999 3.3 0.00178518 3.3 0.00178528 0 0.0017851999999999998 0 0.0017852999999999999 3.3 0.00178522 3.3 0.00178532 0 0.00178524 0 0.00178534 3.3 0.0017852599999999999 3.3 0.00178536 0 0.00178528 0 0.00178538 3.3 0.0017852999999999999 3.3 0.0017854 0 0.00178532 0 0.00178542 3.3 0.0017853399999999998 3.3 0.00178544 0 0.00178536 0 0.00178546 3.3 0.0017853799999999998 3.3 0.0017854799999999999 0 0.0017854 0 0.0017855 3.3 0.0017854199999999998 3.3 0.0017855199999999999 0 0.00178544 0 0.00178554 3.3 0.00178546 3.3 0.00178556 0 0.0017854799999999999 0 0.00178558 3.3 0.0017855 3.3 0.0017856 0 0.0017855199999999999 0 0.00178562 3.3 0.00178554 3.3 0.00178564 0 0.0017855599999999998 0 0.00178566 3.3 0.00178558 3.3 0.00178568 0 0.0017855999999999998 0 0.0017856999999999999 3.3 0.00178562 3.3 0.00178572 0 0.00178564 0 0.00178574 3.3 0.00178566 3.3 0.00178576 0 0.00178568 0 0.00178578 3.3 0.0017856999999999999 3.3 0.0017858 0 0.00178572 0 0.00178582 3.3 0.0017857399999999999 3.3 0.00178584 0 0.00178576 0 0.00178586 3.3 0.0017857799999999998 3.3 0.0017858799999999999 0 0.0017858 0 0.0017859 3.3 0.0017858199999999998 3.3 0.0017859199999999999 0 0.00178584 0 0.00178594 3.3 0.00178586 3.3 0.00178596 0 0.0017858799999999999 0 0.00178598 3.3 0.0017859 3.3 0.001786 0 0.0017859199999999999 0 0.00178602 3.3 0.00178594 3.3 0.00178604 0 0.0017859599999999998 0 0.00178606 3.3 0.00178598 3.3 0.00178608 0 0.0017859999999999998 0 0.0017860999999999999 3.3 0.00178602 3.3 0.00178612 0 0.0017860399999999998 0 0.0017861399999999999 3.3 0.00178606 3.3 0.00178616 0 0.00178608 0 0.00178618 3.3 0.0017860999999999999 3.3 0.0017862 0 0.00178612 0 0.00178622 3.3 0.0017861399999999999 3.3 0.00178624 0 0.00178616 0 0.00178626 3.3 0.0017861799999999998 3.3 0.00178628 0 0.0017862 0 0.0017863 3.3 0.0017862199999999998 3.3 0.0017863199999999999 0 0.00178624 0 0.00178634 3.3 0.0017862599999999998 3.3 0.0017863599999999999 0 0.00178628 0 0.00178638 3.3 0.0017863 3.3 0.0017864 0 0.0017863199999999999 0 0.00178642 3.3 0.00178634 3.3 0.00178644 0 0.0017863599999999999 0 0.00178646 3.3 0.00178638 3.3 0.00178648 0 0.0017863999999999998 0 0.0017865 3.3 0.00178642 3.3 0.00178652 0 0.0017864399999999998 0 0.0017865399999999999 3.3 0.00178646 3.3 0.00178656 0 0.00178648 0 0.00178658 3.3 0.0017865 3.3 0.0017866 0 0.00178652 0 0.00178662 3.3 0.0017865399999999999 3.3 0.00178664 0 0.00178656 0 0.00178666 3.3 0.0017865799999999999 3.3 0.00178668 0 0.0017866 0 0.0017867 3.3 0.0017866199999999998 3.3 0.0017867199999999999 0 0.00178664 0 0.00178674 3.3 0.0017866599999999998 3.3 0.0017867599999999999 0 0.00178668 0 0.00178678 3.3 0.0017867 3.3 0.0017868 0 0.0017867199999999999 0 0.00178682 3.3 0.00178674 3.3 0.00178684 0 0.0017867599999999999 0 0.00178686 3.3 0.00178678 3.3 0.00178688 0 0.0017867999999999998 0 0.0017869 3.3 0.00178682 3.3 0.00178692 0 0.0017868399999999998 0 0.0017869399999999999 3.3 0.00178686 3.3 0.00178696 0 0.0017868799999999998 0 0.0017869799999999999 3.3 0.0017869 3.3 0.001787 0 0.00178692 0 0.00178702 3.3 0.0017869399999999999 3.3 0.00178704 0 0.00178696 0 0.00178706 3.3 0.0017869799999999999 3.3 0.00178708 0 0.001787 0 0.0017871 3.3 0.0017870199999999998 3.3 0.00178712 0 0.00178704 0 0.00178714 3.3 0.0017870599999999998 3.3 0.0017871599999999999 0 0.00178708 0 0.00178718 3.3 0.0017870999999999998 3.3 0.0017871999999999999 0 0.00178712 0 0.00178722 3.3 0.00178714 3.3 0.00178724 0 0.0017871599999999999 0 0.00178726 3.3 0.00178718 3.3 0.00178728 0 0.0017871999999999999 0 0.0017873 3.3 0.00178722 3.3 0.00178732 0 0.0017872399999999998 0 0.00178734 3.3 0.00178726 3.3 0.00178736 0 0.0017872399999999998 0 0.00178734 3.3)

* resetn - 1 transitions
V_resetn resetn 0 PWL(0 0 1.3999999999999998e-07 0 2.4e-07 3.3)

* spi_miso - 3405 transitions
V_spi_miso spi_miso 0 PWL(0 0 1.9020000000000002e-06 0 2.002e-06 3.3 2.142e-06 3.3 2.242e-06 0 4.302e-06 0 4.4019999999999995e-06 3.3 4.542e-06 3.3 4.642e-06 0 4.6620000000000004e-06 0 4.762e-06 3.3 5.022e-06 3.3 5.122e-06 0 5.862e-06 0 5.962e-06 3.3 5.982e-06 3.3 6.0819999999999995e-06 0 6.822e-06 0 6.922e-06 3.3 6.942e-06 3.3 7.042e-06 0 9.821999999999998e-06 0 9.922e-06 3.3 1.0062e-05 3.3 1.0162e-05 0 1.2342e-05 0 1.2442e-05 3.3 1.2461999999999999e-05 3.3 1.2562e-05 0 1.2702e-05 0 1.2802e-05 3.3 1.2941999999999999e-05 3.3 1.3042e-05 0 1.3782e-05 0 1.3882e-05 3.3 1.3901999999999998e-05 3.3 1.4001999999999999e-05 0 1.4741999999999999e-05 0 1.4842e-05 3.3 1.4862e-05 3.3 1.4962e-05 0 1.5462000000000002e-05 0 1.5562e-05 3.3 1.5582e-05 3.3 1.5682e-05 0 1.5822000000000002e-05 0 1.5922e-05 3.3 1.5982e-05 3.3 1.6082e-05 0 1.7742e-05 0 1.7842e-05 3.3 1.7982e-05 3.3 1.8082e-05 0 1.9902e-05 0 2.0002e-05 3.3 2.0022e-05 3.3 2.0121999999999998e-05 0 2.0262e-05 0 2.0362e-05 3.3 2.0382e-05 3.3 2.0481999999999998e-05 0 2.0622e-05 0 2.0722e-05 3.3 2.0862e-05 3.3 2.0962e-05 0 2.1582e-05 0 2.1682e-05 3.3 2.1702e-05 3.3 2.1802e-05 0 2.1942e-05 0 2.2042e-05 3.3 2.2182000000000002e-05 3.3 2.2282e-05 0 2.3622000000000002e-05 0 2.3722e-05 3.3 2.3742e-05 3.3 2.3842e-05 0 2.5662e-05 0 2.5762e-05 3.3 2.5902e-05 3.3 2.6002e-05 0 2.8182e-05 0 2.8281999999999998e-05 3.3 2.8302e-05 3.3 2.8402e-05 0 2.8542e-05 0 2.8641999999999998e-05 3.3 2.8782e-05 3.3 2.8882e-05 0 2.9502e-05 0 2.9602e-05 3.3 2.9742e-05 3.3 2.9842e-05 0 2.9982000000000002e-05 0 3.0082e-05 3.3 3.0102e-05 3.3 3.0202e-05 0 3.1302e-05 0 3.1402e-05 3.3 3.1422e-05 3.3 3.1522e-05 0 3.3582e-05 0 3.3682e-05 3.3 3.3821999999999996e-05 3.3 3.3922e-05 0 3.6101999999999994e-05 0 3.6201999999999997e-05 3.3 3.6222e-05 3.3 3.6322e-05 0 3.6462e-05 0 3.6562e-05 3.3 3.6701999999999995e-05 3.3 3.6802e-05 0 3.7301999999999996e-05 0 3.7402e-05 3.3 3.7421999999999995e-05 3.3 3.7522e-05 0 3.7541999999999994e-05 0 3.7641999999999996e-05 3.3 3.7902e-05 3.3 3.8002e-05 0 3.9102e-05 0 3.9202e-05 3.3 3.9222e-05 3.3 3.9322e-05 0 3.9461999999999996e-05 0 3.9562e-05 3.3 3.9742e-05 3.3 3.9842e-05 0 4.1502e-05 0 4.1602e-05 3.3 4.1741999999999994e-05 3.3 4.1842e-05 0 4.3661999999999996e-05 0 4.3762e-05 3.3 4.4022e-05 3.3 4.4122e-05 0 4.4142e-05 0 4.4242e-05 3.3 4.4621999999999994e-05 3.3 4.4721999999999996e-05 0 4.5582e-05 0 4.5682e-05 3.3 4.5821999999999996e-05 3.3 4.5922e-05 0 4.7142e-05 0 4.7242e-05 3.3 4.7261999999999996e-05 3.3 4.7362e-05 0 4.7381999999999995e-05 0 4.7482e-05 3.3 4.7662e-05 3.3 4.7762e-05 0 4.9421999999999995e-05 0 4.9522e-05 3.3 4.9662e-05 3.3 4.9762e-05 0 5.1942e-05 0 5.2042e-05 3.3 5.2062e-05 3.3 5.2162e-05 0 5.2301999999999995e-05 0 5.2402e-05 3.3 5.2542e-05 3.3 5.2642e-05 0 5.3382e-05 0 5.3482e-05 3.3 5.3741999999999995e-05 3.3 5.3842e-05 0 5.4341999999999996e-05 0 5.4442e-05 3.3 5.5422e-05 3.3 5.5522e-05 0 5.7341999999999994e-05 0 5.7441999999999997e-05 3.3 5.7582e-05 3.3 5.7682e-05 0 5.9742e-05 0 5.9842e-05 3.3 5.9862e-05 3.3 5.9962e-05 0 6.0221999999999994e-05 0 6.0321999999999996e-05 3.3 6.0462e-05 3.3 6.0562e-05 0 6.0701999999999996e-05 0 6.0802e-05 3.3 6.0821999999999995e-05 3.3 6.0922e-05 0 6.1782e-05 0 6.1882e-05 3.3 6.190199999999999e-05 3.3 6.2002e-05 0 6.2262e-05 0 6.2362e-05 3.3 6.2382e-05 3.3 6.2482e-05 0 6.334199999999999e-05 0 6.3442e-05 3.3 6.7542e-05 3.3 6.7642e-05 0 6.9222e-05 0 6.9322e-05 3.3 6.9462e-05 3.3 6.9562e-05 0 7.1382e-05 0 7.1482e-05 3.3 7.1502e-05 3.3 7.1602e-05 0 7.174199999999999e-05 0 7.1842e-05 3.3 7.1862e-05 3.3 7.1962e-05 0 7.2102e-05 0 7.2202e-05 3.3 7.234199999999999e-05 3.3 7.2442e-05 0 7.3062e-05 0 7.3162e-05 3.3 7.3302e-05 3.3 7.3402e-05 0 7.3902e-05 0 7.4002e-05 3.3 7.402199999999999e-05 3.3 7.412199999999999e-05 0 7.4142e-05 0 7.4242e-05 3.3 7.4262e-05 3.3 7.4362e-05 0 7.7142e-05 0 7.7242e-05 3.3 7.7382e-05 3.3 7.7482e-05 0 8.0022e-05 0 8.0122e-05 3.3 8.0502e-05 3.3 8.0602e-05 0 8.0862e-05 0 8.0962e-05 3.3 8.098199999999999e-05 3.3 8.1082e-05 0 8.1102e-05 0 8.1202e-05 3.3 8.1222e-05 3.3 8.1322e-05 0 8.1942e-05 0 8.2042e-05 3.3 8.2182e-05 3.3 8.2282e-05 0 8.4942e-05 0 8.5042e-05 3.3 8.5182e-05 3.3 8.5282e-05 0 8.7222e-05 0 8.7322e-05 3.3 8.734199999999999e-05 3.3 8.7442e-05 0 8.758199999999999e-05 0 8.768199999999999e-05 3.3 8.7702e-05 3.3 8.7802e-05 0 8.794199999999999e-05 0 8.8042e-05 3.3 8.8062e-05 3.3 8.8162e-05 0 8.818199999999999e-05 0 8.828199999999999e-05 3.3 8.8422e-05 3.3 8.8522e-05 0 8.8542e-05 0 8.8642e-05 3.3 8.8902e-05 3.3 8.9002e-05 0 8.9502e-05 0 8.9602e-05 3.3 8.962199999999999e-05 3.3 8.972199999999999e-05 0 8.9742e-05 0 8.9842e-05 3.3 8.9862e-05 3.3 8.9962e-05 0 9.2742e-05 0 9.2842e-05 3.3 9.2982e-05 3.3 9.3082e-05 0 9.5022e-05 0 9.5122e-05 3.3 9.5262e-05 3.3 9.5362e-05 0 9.5622e-05 0 9.5722e-05 3.3 9.5862e-05 3.3 9.5962e-05 0 9.6342e-05 0 9.6442e-05 3.3 9.6462e-05 3.3 9.6562e-05 0 9.742199999999999e-05 0 9.752199999999999e-05 3.3 9.7542e-05 3.3 9.7642e-05 0 9.7662e-05 0 9.7762e-05 3.3 9.778199999999999e-05 3.3 9.7882e-05 0 9.8742e-05 0 9.8842e-05 3.3 9.8902e-05 3.3 9.9002e-05 0 0.00010066199999999999 0 0.000100762 3.3 0.00010090199999999999 3.3 0.00010100199999999999 0 0.000102822 0 0.000102922 3.3 0.00010318199999999999 3.3 0.00010328199999999999 0 0.000103302 0 0.000103402 3.3 0.00010378199999999999 3.3 0.00010388199999999999 0 0.000104742 0 0.000104842 3.3 0.000104862 3.3 0.000104962 0 0.000105942 0 0.000106042 3.3 0.000106062 3.3 0.000106162 0 0.000106182 0 0.000106282 3.3 0.000106302 3.3 0.000106402 0 0.00010642199999999999 0 0.000106522 3.3 0.000106542 3.3 0.000106642 0 0.00010666199999999999 0 0.00010676199999999999 3.3 0.000106822 3.3 0.000106922 0 0.000108582 0 0.000108682 3.3 0.000108822 3.3 0.000108922 0 0.000110502 0 0.000110602 3.3 0.00011074199999999999 3.3 0.000110842 0 0.000111102 0 0.000111202 3.3 0.000111222 3.3 0.000111322 0 0.000111462 0 0.000111562 3.3 0.000111702 3.3 0.000111802 0 0.000112542 0 0.000112642 3.3 0.00011278199999999999 3.3 0.000112882 0 0.000113502 0 0.000113602 3.3 0.000114582 3.3 0.000114682 0 0.00011650199999999999 0 0.00011660199999999999 3.3 0.000116742 3.3 0.000116842 0 0.000118422 0 0.000118522 3.3 0.000118662 3.3 0.000118762 0 0.000118902 0 0.000119002 3.3 0.000119022 3.3 0.000119122 0 0.00011938199999999999 0 0.00011948199999999999 3.3 0.000119622 3.3 0.000119722 0 0.000119862 0 0.000119962 3.3 0.00011998199999999999 3.3 0.00012008199999999999 0 0.000120702 0 0.000120802 3.3 0.00012082199999999999 3.3 0.00012092199999999999 0 0.000120942 0 0.000121042 3.3 0.000121062 3.3 0.000121162 0 0.00012142199999999999 0 0.00012152199999999999 3.3 0.000121542 3.3 0.000121642 0 0.000128382 0 0.000128482 3.3 0.000128622 3.3 0.000128722 0 0.000130302 0 0.000130402 3.3 0.00013054199999999998 3.3 0.000130642 0 0.000130782 0 0.000130882 3.3 0.000130902 3.3 0.000131002 0 0.000131262 0 0.000131362 3.3 0.000131502 3.3 0.000131602 0 0.000131742 0 0.000131842 3.3 0.000131862 3.3 0.000131962 0 0.00013222199999999998 0 0.00013232199999999998 3.3 0.000132342 3.3 0.000132442 0 0.00013258199999999999 0 0.000132682 3.3 0.000132822 3.3 0.000132922 0 0.000133302 0 0.000133402 3.3 0.00013342199999999998 3.3 0.00013352199999999999 0 0.000134382 0 0.000134482 3.3 0.000138582 3.3 0.000138682 0 0.000140262 0 0.000140362 3.3 0.000140502 3.3 0.000140602 0 0.000142182 0 0.000142282 3.3 0.000142542 3.3 0.000142642 0 0.000142662 0 0.000142762 3.3 0.00014290199999999998 3.3 0.00014300199999999998 0 0.000143022 0 0.000143122 3.3 0.000143382 3.3 0.000143482 0 0.000144222 0 0.000144322 3.3 0.000144342 3.3 0.000144442 0 0.000144462 0 0.000144562 3.3 0.000144582 3.3 0.000144682 0 0.00014818199999999998 0 0.000148282 3.3 0.000148422 3.3 0.000148522 0 0.000150102 0 0.000150202 3.3 0.000150342 3.3 0.000150442 0 0.000150582 0 0.000150682 3.3 0.00015070199999999998 3.3 0.00015080199999999998 0 0.00015106199999999998 0 0.000151162 3.3 0.000151422 3.3 0.000151522 0 0.000151542 0 0.000151642 3.3 0.000151662 3.3 0.000151762 0 0.00015190199999999998 0 0.00015200199999999999 3.3 0.000152022 3.3 0.000152122 0 0.000152262 0 0.000152362 3.3 0.000152382 3.3 0.000152482 0 0.000152502 0 0.000152602 3.3 0.000152622 3.3 0.000152722 0 0.00015310199999999999 0 0.000153202 3.3 0.000153222 3.3 0.000153322 0 0.000154182 0 0.000154282 3.3 0.000154422 3.3 0.000154522 0 0.000156102 0 0.000156202 3.3 0.000156342 3.3 0.000156442 0 0.00015802199999999999 0 0.000158122 3.3 0.000158382 3.3 0.000158482 0 0.000158622 0 0.000158722 3.3 0.000158742 3.3 0.000158842 0 0.000158982 0 0.000159082 3.3 0.000159222 3.3 0.000159322 0 0.000159942 0 0.000160042 3.3 0.00016006199999999999 3.3 0.000160162 0 0.000160182 0 0.000160282 3.3 0.000160302 3.3 0.000160402 0 0.000164022 0 0.000164122 3.3 0.000164262 3.3 0.000164362 0 0.000165942 0 0.000166042 3.3 0.000166182 3.3 0.000166282 0 0.000166422 0 0.000166522 3.3 0.000166542 3.3 0.000166642 0 0.000166902 0 0.000167002 3.3 0.000167262 3.3 0.000167362 0 0.000167382 0 0.000167482 3.3 0.00016750199999999998 3.3 0.00016760199999999999 0 0.000167622 0 0.000167722 3.3 0.000167742 3.3 0.000167842 0 0.000168222 0 0.000168322 3.3 0.00016834199999999998 3.3 0.00016844199999999998 0 0.000168462 0 0.000168562 3.3 0.000168582 3.3 0.000168682 0 0.000168942 0 0.000169042 3.3 0.000169062 3.3 0.000169162 0 0.000170022 0 0.000170122 3.3 0.000170262 3.3 0.000170362 0 0.000171942 0 0.000172042 3.3 0.000172182 3.3 0.000172282 0 0.000173862 0 0.000173962 3.3 0.000174222 3.3 0.000174322 0 0.00017446199999999998 0 0.000174562 3.3 0.000174582 3.3 0.000174682 0 0.000174822 0 0.000174922 3.3 0.000175062 3.3 0.000175162 0 0.000175782 0 0.000175882 3.3 0.000175902 3.3 0.000176002 0 0.000179862 0 0.000179962 3.3 0.000180102 3.3 0.000180202 0 0.000181782 0 0.000181882 3.3 0.000182022 3.3 0.000182122 0 0.00018226199999999998 0 0.00018236199999999999 3.3 0.000182382 3.3 0.000182482 0 0.000182742 0 0.000182842 3.3 0.00018310199999999998 3.3 0.00018320199999999999 0 0.000183222 0 0.000183322 3.3 0.000183342 3.3 0.000183442 0 0.00018346199999999999 0 0.000183562 3.3 0.000183582 3.3 0.000183682 0 0.000184062 0 0.000184162 3.3 0.000184182 3.3 0.000184282 0 0.00018430199999999998 0 0.000184402 3.3 0.000184422 3.3 0.000184522 0 0.000184782 0 0.000184882 3.3 0.000184902 3.3 0.000185002 0 0.000185862 0 0.000185962 3.3 0.000186102 3.3 0.000186202 0 0.000187782 0 0.000187882 3.3 0.00018802199999999998 3.3 0.00018812199999999999 0 0.00018970199999999998 0 0.00018980199999999998 3.3 0.00019006199999999998 3.3 0.00019016199999999999 0 0.000190302 0 0.000190402 3.3 0.000190422 3.3 0.000190522 0 0.000190662 0 0.000190762 3.3 0.00019090199999999998 3.3 0.00019100199999999998 0 0.000191622 0 0.000191722 3.3 0.00019174199999999998 3.3 0.00019184199999999998 0 0.000193062 0 0.000193162 3.3 0.000193182 3.3 0.000193282 0 0.000195702 0 0.000195802 3.3 0.000195942 3.3 0.000196042 0 0.000197622 0 0.000197722 3.3 0.00019786199999999998 3.3 0.00019796199999999999 0 0.000198582 0 0.000198682 3.3 0.000198942 3.3 0.000199042 0 0.00019906199999999999 0 0.000199162 3.3 0.000199182 3.3 0.000199282 0 0.00019954199999999998 0 0.00019964199999999998 3.3 0.000199782 3.3 0.000199882 0 0.000200622 0 0.000200722 3.3 0.00020074199999999998 3.3 0.00020084199999999999 0 0.00020158199999999998 0 0.00020168199999999998 3.3 0.000201702 3.3 0.000201802 0 0.00020362199999999998 0 0.00020372199999999999 3.3 0.000203862 3.3 0.000203962 0 0.000205542 0 0.000205642 3.3 0.000205782 3.3 0.000205882 0 0.000206022 0 0.000206122 3.3 0.000206262 3.3 0.000206362 0 0.00020650199999999998 0 0.00020660199999999998 3.3 0.000206742 3.3 0.000206842 0 0.00020686199999999999 0 0.000206962 3.3 0.000207222 3.3 0.000207322 0 0.000207462 0 0.000207562 3.3 0.00020770199999999998 3.3 0.000207802 0 0.000207822 0 0.000207922 3.3 0.000207942 3.3 0.000208042 0 0.000208062 0 0.000208162 3.3 0.000208182 3.3 0.000208282 0 0.000208422 0 0.000208522 3.3 0.000208662 3.3 0.000208762 0 0.000209622 0 0.000209722 3.3 0.000209782 3.3 0.000209882 0 0.000211542 0 0.000211642 3.3 0.00021178199999999999 3.3 0.000211882 0 0.00021346199999999998 0 0.00021356199999999999 3.3 0.000214062 3.3 0.000214162 0 0.000214422 0 0.000214522 3.3 0.00021466199999999999 3.3 0.000214762 0 0.000215022 0 0.000215122 3.3 0.000215382 3.3 0.000215482 0 0.00021634199999999998 0 0.00021644199999999999 3.3 0.000217422 3.3 0.000217522 0 0.00021754199999999998 0 0.000217642 3.3 0.00021770199999999998 3.3 0.00021780199999999999 0 0.000219462 0 0.000219562 3.3 0.000219702 3.3 0.000219802 0 0.000221382 0 0.000221482 3.3 0.000221622 3.3 0.000221722 0 0.000222342 0 0.000222442 3.3 0.000222702 3.3 0.000222802 0 0.000222822 0 0.000222922 3.3 0.00022294199999999998 3.3 0.00022304199999999998 0 0.00022330199999999998 0 0.00022340199999999999 3.3 0.000223542 3.3 0.000223642 0 0.000224382 0 0.000224482 3.3 0.00022450199999999999 3.3 0.000224602 0 0.00022534199999999998 0 0.000225442 3.3 0.000225462 3.3 0.000225562 0 0.00022738199999999999 0 0.000227482 3.3 0.000227622 3.3 0.000227722 0 0.000229302 0 0.000229402 3.3 0.000229542 3.3 0.000229642 0 0.000229782 0 0.000229882 3.3 0.000230022 3.3 0.000230122 0 0.00023026199999999999 0 0.000230362 3.3 0.000230502 3.3 0.000230602 0 0.000230622 0 0.000230722 3.3 0.000230982 3.3 0.000231082 0 0.000231222 0 0.000231322 3.3 0.000231462 3.3 0.000231562 0 0.000231582 0 0.000231682 3.3 0.000231702 3.3 0.000231802 0 0.000231822 0 0.000231922 3.3 0.00023194199999999998 3.3 0.00023204199999999999 0 0.000232182 0 0.000232282 3.3 0.000232422 3.3 0.000232522 0 0.000233382 0 0.000233482 3.3 0.000233542 3.3 0.000233642 0 0.000235302 0 0.000235402 3.3 0.000235542 3.3 0.000235642 0 0.00023722199999999999 0 0.000237322 3.3 0.000237822 3.3 0.000237922 0 0.000238182 0 0.000238282 3.3 0.000238422 3.3 0.000238522 0 0.000238782 0 0.000238882 3.3 0.000239142 3.3 0.000239242 0 0.00024010199999999999 0 0.000240202 3.3 0.000241182 3.3 0.000241282 0 0.000241302 0 0.000241402 3.3 0.00024146199999999999 3.3 0.000241562 0 0.000243222 0 0.000243322 3.3 0.00024346199999999998 3.3 0.00024356199999999998 0 0.000245142 0 0.000245242 3.3 0.000245382 3.3 0.000245482 0 0.000246102 0 0.000246202 3.3 0.00024646199999999997 3.3 0.000246562 0 0.000246582 0 0.000246682 3.3 0.000246702 3.3 0.000246802 0 0.000247062 0 0.000247162 3.3 0.00024730199999999997 3.3 0.000247402 0 0.00024814199999999997 0 0.00024824199999999997 3.3 0.000248262 3.3 0.000248362 0 0.000249102 0 0.000249202 3.3 0.000249222 3.3 0.000249322 0 0.000251142 0 0.000251242 3.3 0.00025138199999999997 3.3 0.000251482 0 0.00025306199999999997 0 0.00025316199999999997 3.3 0.000253302 3.3 0.000253402 0 0.000253542 0 0.000253642 3.3 0.000253782 3.3 0.000253882 0 0.000254022 0 0.000254122 3.3 0.000254262 3.3 0.000254362 0 0.000254382 0 0.000254482 3.3 0.00025474199999999997 3.3 0.00025484199999999997 0 0.000254982 0 0.000255082 3.3 0.000255222 3.3 0.000255322 0 0.000255342 0 0.000255442 3.3 0.000255462 3.3 0.000255562 0 0.00025558199999999997 0 0.00025568199999999997 3.3 0.000255702 3.3 0.000255802 0 0.000255942 0 0.000256042 3.3 0.000256182 3.3 0.000256282 0 0.00025714199999999997 0 0.000257242 3.3 0.000257302 3.3 0.000257402 0 0.000259062 0 0.000259162 3.3 0.000259302 3.3 0.000259402 0 0.000260982 0 0.000261082 3.3 0.000261582 3.3 0.000261682 0 0.000261942 0 0.000262042 3.3 0.000262182 3.3 0.000262282 0 0.000262542 0 0.000262642 3.3 0.00026290199999999997 3.3 0.000263002 0 0.000263862 0 0.000263962 3.3 0.000264942 3.3 0.000265042 0 0.000265062 0 0.000265162 3.3 0.000265222 3.3 0.000265322 0 0.00026698199999999997 0 0.000267082 3.3 0.000267222 3.3 0.000267322 0 0.000268902 0 0.000269002 3.3 0.000269142 3.3 0.000269242 0 0.000269862 0 0.000269962 3.3 0.000270222 3.3 0.000270322 0 0.00027034199999999997 0 0.00027044199999999997 3.3 0.000270462 3.3 0.000270562 0 0.000270822 0 0.000270922 3.3 0.000271062 3.3 0.000271162 0 0.00027190199999999997 0 0.000272002 3.3 0.000272022 3.3 0.000272122 0 0.000272862 0 0.000272962 3.3 0.000272982 3.3 0.000273082 0 0.000274902 0 0.000275002 3.3 0.000275142 3.3 0.000275242 0 0.000276822 0 0.000276922 3.3 0.000277062 3.3 0.000277162 0 0.000277302 0 0.000277402 3.3 0.000277542 3.3 0.000277642 0 0.000277782 0 0.000277882 3.3 0.000278022 3.3 0.000278122 0 0.000278142 0 0.000278242 3.3 0.00027850199999999997 3.3 0.000278602 0 0.000278742 0 0.000278842 3.3 0.000278982 3.3 0.000279082 0 0.000279102 0 0.000279202 3.3 0.000279222 3.3 0.000279322 0 0.00027934199999999997 0 0.00027944199999999997 3.3 0.000279462 3.3 0.000279562 0 0.000279702 0 0.000279802 3.3 0.000279942 3.3 0.000280042 0 0.000280902 0 0.000281002 3.3 0.000281062 3.3 0.000281162 0 0.000282822 0 0.000282922 3.3 0.000283062 3.3 0.000283162 0 0.000284742 0 0.000284842 3.3 0.000285342 3.3 0.000285442 0 0.000285702 0 0.000285802 3.3 0.00028594199999999997 3.3 0.00028604199999999997 0 0.000286302 0 0.000286402 3.3 0.000286662 3.3 0.000286762 0 0.000287622 0 0.000287722 3.3 0.000288702 3.3 0.000288802 0 0.000288822 0 0.000288922 3.3 0.00028898199999999997 3.3 0.00028908199999999997 0 0.000290742 0 0.000290842 3.3 0.000290982 3.3 0.000291082 0 0.000292662 0 0.000292762 3.3 0.000292902 3.3 0.000293002 0 0.000293622 0 0.000293722 3.3 0.000293982 3.3 0.000294082 0 0.00029410199999999997 0 0.00029420199999999997 3.3 0.000294222 3.3 0.000294322 0 0.000294582 0 0.000294682 3.3 0.000294822 3.3 0.000294922 0 0.000295662 0 0.000295762 3.3 0.00029578199999999997 3.3 0.00029588199999999997 0 0.00029662199999999997 0 0.00029672199999999997 3.3 0.000296742 3.3 0.000296842 0 0.000298662 0 0.000298762 3.3 0.000298902 3.3 0.000299002 0 0.000300582 0 0.000300682 3.3 0.000300822 3.3 0.000300922 0 0.000301062 0 0.000301162 3.3 0.000301302 3.3 0.000301402 0 0.00030154199999999997 0 0.00030164199999999997 3.3 0.000301782 3.3 0.000301882 0 0.000301902 0 0.000302002 3.3 0.000302262 3.3 0.000302362 0 0.000302502 0 0.000302602 3.3 0.000302742 3.3 0.000302842 0 0.000302862 0 0.000302962 3.3 0.000302982 3.3 0.000303082 0 0.00030310199999999997 0 0.000303202 3.3 0.000303222 3.3 0.000303322 0 0.000303462 0 0.000303562 3.3 0.000303702 3.3 0.000303802 0 0.000304662 0 0.000304762 3.3 0.000304822 3.3 0.000304922 0 0.000306582 0 0.000306682 3.3 0.000306822 3.3 0.000306922 0 0.000308502 0 0.000308602 3.3 0.000309102 3.3 0.000309202 0 0.000309462 0 0.000309562 3.3 0.00030970199999999997 3.3 0.00030980199999999997 0 0.000310062 0 0.000310162 3.3 0.000310422 3.3 0.000310522 0 0.00031138199999999997 0 0.00031148199999999997 3.3 0.000312462 3.3 0.000312562 0 0.000312582 0 0.000312682 3.3 0.00031274199999999997 3.3 0.00031284199999999997 0 0.000314502 0 0.000314602 3.3 0.000314742 3.3 0.000314842 0 0.000316422 0 0.000316522 3.3 0.000316662 3.3 0.000316762 0 0.000317382 0 0.000317482 3.3 0.000317742 3.3 0.000317842 0 0.000317862 0 0.000317962 3.3 0.00031798199999999997 3.3 0.00031808199999999997 0 0.000318342 0 0.000318442 3.3 0.000318582 3.3 0.000318682 0 0.000319422 0 0.000319522 3.3 0.00031954199999999997 3.3 0.000319642 0 0.00032038199999999997 0 0.00032048199999999997 3.3 0.000320502 3.3 0.000320602 0 0.000322422 0 0.000322522 3.3 0.000322662 3.3 0.000322762 0 0.000324342 0 0.000324442 3.3 0.000324582 3.3 0.000324682 0 0.000324822 0 0.000324922 3.3 0.000325062 3.3 0.000325162 0 0.00032530199999999997 0 0.00032540199999999997 3.3 0.000325542 3.3 0.000325642 0 0.000325662 0 0.000325762 3.3 0.000326022 3.3 0.000326122 0 0.000326262 0 0.000326362 3.3 0.000326502 3.3 0.000326602 0 0.000326622 0 0.000326722 3.3 0.000326742 3.3 0.000326842 0 0.000326862 0 0.000326962 3.3 0.00032698199999999997 3.3 0.00032708199999999997 0 0.000327222 0 0.000327322 3.3 0.000327462 3.3 0.000327562 0 0.000328422 0 0.000328522 3.3 0.000328582 3.3 0.000328682 0 0.000330342 0 0.000330442 3.3 0.000330582 3.3 0.000330682 0 0.000332262 0 0.000332362 3.3 0.000332862 3.3 0.000332962 0 0.000333222 0 0.000333322 3.3 0.00033346199999999997 3.3 0.000333562 0 0.000333822 0 0.000333922 3.3 0.000334182 3.3 0.000334282 0 0.00033514199999999997 0 0.00033524199999999997 3.3 0.000336222 3.3 0.000336322 0 0.000336342 0 0.000336442 3.3 0.00033650199999999997 3.3 0.000336602 0 0.000338262 0 0.000338362 3.3 0.00033850199999999997 3.3 0.00033860199999999997 0 0.000340182 0 0.000340282 3.3 0.000340422 3.3 0.000340522 0 0.000341142 0 0.000341242 3.3 0.000341502 3.3 0.000341602 0 0.000341622 0 0.000341722 3.3 0.00034174199999999997 3.3 0.00034184199999999997 0 0.000342102 0 0.000342202 3.3 0.000342342 3.3 0.000342442 0 0.000343182 0 0.000343282 3.3 0.000343302 3.3 0.000343402 0 0.00034414199999999997 0 0.000344242 3.3 0.00034426199999999996 3.3 0.00034436199999999997 0 0.000346182 0 0.000346282 3.3 0.000346422 3.3 0.000346522 0 0.000348102 0 0.000348202 3.3 0.00034834199999999997 3.3 0.00034844199999999997 0 0.000348582 0 0.000348682 3.3 0.000348822 3.3 0.000348922 0 0.00034906199999999997 0 0.000349162 3.3 0.000349302 3.3 0.000349402 0 0.000349422 0 0.000349522 3.3 0.000349782 3.3 0.000349882 0 0.000350022 0 0.000350122 3.3 0.000350262 3.3 0.000350362 0 0.000350382 0 0.000350482 3.3 0.000350502 3.3 0.000350602 0 0.000350622 0 0.000350722 3.3 0.00035074199999999997 3.3 0.00035084199999999997 0 0.000350982 0 0.000351082 3.3 0.000351222 3.3 0.000351322 0 0.000352182 0 0.000352282 3.3 0.000352342 3.3 0.000352442 0 0.00035410199999999996 0 0.00035420199999999997 3.3 0.000354342 3.3 0.000354442 0 0.000356022 0 0.000356122 3.3 0.000356622 3.3 0.000356722 0 0.000356982 0 0.000357082 3.3 0.000357222 3.3 0.000357322 0 0.000357582 0 0.000357682 3.3 0.000357942 3.3 0.000358042 0 0.000358902 0 0.000359002 3.3 0.000359982 3.3 0.000360082 0 0.000360102 0 0.000360202 3.3 0.000360262 3.3 0.000360362 0 0.000362022 0 0.000362122 3.3 0.00036226199999999997 3.3 0.00036236199999999997 0 0.00036394199999999997 0 0.00036404199999999997 3.3 0.000364182 3.3 0.000364282 0 0.000364902 0 0.000365002 3.3 0.000365262 3.3 0.000365362 0 0.000365382 0 0.000365482 3.3 0.00036550199999999997 3.3 0.000365602 0 0.000365862 0 0.000365962 3.3 0.000366102 3.3 0.000366202 0 0.000366942 0 0.000367042 3.3 0.000367062 3.3 0.000367162 0 0.000367902 0 0.000368002 3.3 0.00036802199999999997 3.3 0.00036812199999999997 0 0.000369942 0 0.000370042 3.3 0.000370182 3.3 0.000370282 0 0.000371862 0 0.000371962 3.3 0.00037210199999999997 3.3 0.00037220199999999997 0 0.000372342 0 0.000372442 3.3 0.000372582 3.3 0.000372682 0 0.000372822 0 0.000372922 3.3 0.000373062 3.3 0.000373162 0 0.000373182 0 0.000373282 3.3 0.000373542 3.3 0.000373642 0 0.00037378199999999997 0 0.00037388199999999997 3.3 0.000374022 3.3 0.000374122 0 0.000374142 0 0.000374242 3.3 0.000374262 3.3 0.000374362 0 0.000374382 0 0.000374482 3.3 0.000374502 3.3 0.000374602 0 0.000374742 0 0.000374842 3.3 0.000374982 3.3 0.000375082 0 0.000375942 0 0.000376042 3.3 0.000376102 3.3 0.000376202 0 0.00037786199999999997 0 0.00037796199999999997 3.3 0.000378102 3.3 0.000378202 0 0.000379782 0 0.000379882 3.3 0.00038038199999999996 3.3 0.00038048199999999997 0 0.000380742 0 0.000380842 3.3 0.000380982 3.3 0.000381082 0 0.000381342 0 0.000381442 3.3 0.000381702 3.3 0.000381802 0 0.000382662 0 0.000382762 3.3 0.000383742 3.3 0.000383842 0 0.000383862 0 0.000383962 3.3 0.000384022 3.3 0.000384122 0 0.000385782 0 0.000385882 3.3 0.00038602199999999997 3.3 0.000386122 0 0.00038770199999999997 0 0.00038780199999999997 3.3 0.000387942 3.3 0.000388042 0 0.000388662 0 0.000388762 3.3 0.000389022 3.3 0.000389122 0 0.000389142 0 0.000389242 3.3 0.000389262 3.3 0.000389362 0 0.000389622 0 0.000389722 3.3 0.000389862 3.3 0.000389962 0 0.000390702 0 0.000390802 3.3 0.000390822 3.3 0.000390922 0 0.000391662 0 0.000391762 3.3 0.00039178199999999997 3.3 0.00039188199999999997 0 0.000393702 0 0.000393802 3.3 0.000393942 3.3 0.000394042 0 0.000395622 0 0.000395722 3.3 0.00039586199999999997 3.3 0.000395962 0 0.000396102 0 0.000396202 3.3 0.000396342 3.3 0.000396442 0 0.000396582 0 0.000396682 3.3 0.00039682199999999996 3.3 0.00039692199999999996 0 0.000396942 0 0.000397042 3.3 0.000397302 3.3 0.000397402 0 0.00039754199999999997 0 0.00039764199999999997 3.3 0.000397782 3.3 0.000397882 0 0.000397902 0 0.000398002 3.3 0.000398022 3.3 0.000398122 0 0.000398142 0 0.000398242 3.3 0.000398262 3.3 0.000398362 0 0.000398502 0 0.000398602 3.3 0.000398742 3.3 0.000398842 0 0.000399702 0 0.000399802 3.3 0.000399862 3.3 0.000399962 0 0.00040162199999999997 0 0.000401722 3.3 0.000401862 3.3 0.000401962 0 0.000403542 0 0.000403642 3.3 0.00040414199999999997 3.3 0.00040424199999999997 0 0.000404502 0 0.000404602 3.3 0.000404742 3.3 0.000404842 0 0.000405102 0 0.000405202 3.3 0.000405462 3.3 0.000405562 0 0.000406422 0 0.000406522 3.3 0.000407502 3.3 0.000407602 0 0.000407622 0 0.000407722 3.3 0.000407782 3.3 0.000407882 0 0.000409542 0 0.000409642 3.3 0.000409782 3.3 0.000409882 0 0.00041146199999999997 0 0.000411562 3.3 0.000411702 3.3 0.000411802 0 0.00041242199999999996 0 0.00041252199999999996 3.3 0.000412782 3.3 0.000412882 0 0.000412902 0 0.000413002 3.3 0.000413022 3.3 0.000413122 0 0.000413382 0 0.000413482 3.3 0.000413622 3.3 0.000413722 0 0.000414462 0 0.000414562 3.3 0.000414582 3.3 0.000414682 0 0.000415422 0 0.000415522 3.3 0.000415542 3.3 0.000415642 0 0.000417462 0 0.000417562 3.3 0.000417702 3.3 0.000417802 0 0.000419382 0 0.000419482 3.3 0.000419622 3.3 0.000419722 0 0.000419862 0 0.000419962 3.3 0.000420102 3.3 0.000420202 0 0.000420342 0 0.000420442 3.3 0.00042058199999999997 3.3 0.00042068199999999997 0 0.000420702 0 0.000420802 3.3 0.000421062 3.3 0.000421162 0 0.00042130199999999997 0 0.000421402 3.3 0.000421542 3.3 0.000421642 0 0.000421662 0 0.000421762 3.3 0.000421782 3.3 0.000421882 0 0.000421902 0 0.000422002 3.3 0.000422022 3.3 0.000422122 0 0.00042226199999999996 0 0.00042236199999999997 3.3 0.000422502 3.3 0.000422602 0 0.000423462 0 0.000423562 3.3 0.00042362199999999996 3.3 0.00042372199999999997 0 0.000425382 0 0.000425482 3.3 0.000425622 3.3 0.000425722 0 0.000427302 0 0.000427402 3.3 0.00042790199999999997 3.3 0.00042800199999999997 0 0.000428262 0 0.000428362 3.3 0.000428502 3.3 0.000428602 0 0.000428862 0 0.000428962 3.3 0.000429222 3.3 0.000429322 0 0.000430182 0 0.000430282 3.3 0.00043126199999999996 3.3 0.00043136199999999997 0 0.000431382 0 0.000431482 3.3 0.000431542 3.3 0.000431642 0 0.000433302 0 0.000433402 3.3 0.000433542 3.3 0.000433642 0 0.000435222 0 0.000435322 3.3 0.000435462 3.3 0.000435562 0 0.00043618199999999997 0 0.00043628199999999997 3.3 0.000436542 3.3 0.000436642 0 0.000436662 0 0.000436762 3.3 0.000436782 3.3 0.000436882 0 0.000437142 0 0.000437242 3.3 0.000437382 3.3 0.000437482 0 0.000438222 0 0.000438322 3.3 0.000438342 3.3 0.000438442 0 0.000439182 0 0.000439282 3.3 0.000439302 3.3 0.000439402 0 0.000441222 0 0.000441322 3.3 0.000441462 3.3 0.000441562 0 0.000443142 0 0.000443242 3.3 0.000443382 3.3 0.000443482 0 0.00044362199999999996 0 0.00044372199999999996 3.3 0.000443862 3.3 0.000443962 0 0.000444102 0 0.000444202 3.3 0.00044434199999999997 3.3 0.00044444199999999997 0 0.000444462 0 0.000444562 3.3 0.000444822 3.3 0.000444922 0 0.000445062 0 0.000445162 3.3 0.000445302 3.3 0.000445402 0 0.000445422 0 0.000445522 3.3 0.000445542 3.3 0.000445642 0 0.000445662 0 0.000445762 3.3 0.000445782 3.3 0.000445882 0 0.00044602199999999997 0 0.00044612199999999997 3.3 0.000446262 3.3 0.000446362 0 0.000447222 0 0.000447322 3.3 0.00044738199999999997 3.3 0.00044748199999999997 0 0.000449142 0 0.000449242 3.3 0.000449382 3.3 0.000449482 0 0.000451062 0 0.000451162 3.3 0.00045166199999999997 3.3 0.000451762 0 0.000452022 0 0.000452122 3.3 0.000452262 3.3 0.000452362 0 0.00045262199999999996 0 0.00045272199999999997 3.3 0.000452982 3.3 0.000453082 0 0.000453942 0 0.000454042 3.3 0.00045502199999999997 3.3 0.00045512199999999997 0 0.000455142 0 0.000455242 3.3 0.000455302 3.3 0.000455402 0 0.000457062 0 0.000457162 3.3 0.000457302 3.3 0.000457402 0 0.000458982 0 0.000459082 3.3 0.00045922199999999996 3.3 0.00045932199999999996 0 0.00045994199999999997 0 0.00046004199999999997 3.3 0.000460302 3.3 0.000460402 0 0.000460422 0 0.000460522 3.3 0.000460542 3.3 0.000460642 0 0.000460902 0 0.000461002 3.3 0.000461142 3.3 0.000461242 0 0.000461982 0 0.000462082 3.3 0.000462102 3.3 0.000462202 0 0.000462942 0 0.000463042 3.3 0.000463062 3.3 0.000463162 0 0.000464982 0 0.000465082 3.3 0.000465222 3.3 0.000465322 0 0.000466902 0 0.000467002 3.3 0.000467142 3.3 0.000467242 0 0.00046738199999999996 0 0.00046748199999999997 3.3 0.000467622 3.3 0.000467722 0 0.000467862 0 0.000467962 3.3 0.00046810199999999997 3.3 0.000468202 0 0.00046822199999999996 0 0.00046832199999999997 3.3 0.000468582 3.3 0.000468682 0 0.000468822 0 0.000468922 3.3 0.00046906199999999996 3.3 0.00046916199999999996 0 0.000469182 0 0.000469282 3.3 0.000469302 3.3 0.000469402 0 0.000469422 0 0.000469522 3.3 0.000469542 3.3 0.000469642 0 0.00046978199999999997 0 0.00046988199999999997 3.3 0.000470022 3.3 0.000470122 0 0.000470982 0 0.000471082 3.3 0.00047114199999999997 3.3 0.00047124199999999997 0 0.000472902 0 0.000473002 3.3 0.00047314199999999996 3.3 0.00047324199999999997 0 0.00047482199999999996 0 0.00047492199999999996 3.3 0.000475422 3.3 0.000475522 0 0.000475782 0 0.000475882 3.3 0.000476022 3.3 0.000476122 0 0.00047638199999999997 0 0.00047648199999999997 3.3 0.000476742 3.3 0.000476842 0 0.000477702 0 0.000477802 3.3 0.00047878199999999997 3.3 0.000478882 0 0.00047890199999999996 0 0.00047900199999999997 3.3 0.000479062 3.3 0.000479162 0 0.000480822 0 0.000480922 3.3 0.000481062 3.3 0.000481162 0 0.000482742 0 0.000482842 3.3 0.00048298199999999996 3.3 0.00048308199999999997 0 0.00048370199999999997 0 0.000483802 3.3 0.000484062 3.3 0.000484162 0 0.000484182 0 0.000484282 3.3 0.000484302 3.3 0.000484402 0 0.00048466199999999996 0 0.00048476199999999996 3.3 0.000484902 3.3 0.000485002 0 0.000485742 0 0.000485842 3.3 0.000485862 3.3 0.000485962 0 0.000486702 0 0.000486802 3.3 0.000486822 3.3 0.000486922 0 0.000488742 0 0.000488842 3.3 0.000488982 3.3 0.000489082 0 0.000490662 0 0.000490762 3.3 0.0004909020000000001 3.3 0.000491002 0 0.0004911420000000001 0 0.000491242 3.3 0.0004913820000000001 3.3 0.000491482 0 0.000491622 0 0.000491722 3.3 0.000491862 3.3 0.000491962 0 0.0004919820000000001 0 0.000492082 3.3 0.000492342 3.3 0.0004924419999999999 0 0.0004925820000000001 0 0.000492682 3.3 0.0004928220000000001 3.3 0.000492922 0 0.000492942 0 0.000493042 3.3 0.0004930620000000001 3.3 0.000493162 0 0.000493182 0 0.0004932819999999999 3.3 0.000493302 3.3 0.000493402 0 0.000493542 0 0.000493642 3.3 0.000493782 3.3 0.000493882 0 0.0004947420000000001 0 0.000494842 3.3 0.0004949020000000001 3.3 0.000495002 0 0.000496662 0 0.000496762 3.3 0.000496902 3.3 0.000497002 0 0.000498582 0 0.000498682 3.3 0.000499182 3.3 0.000499282 0 0.0004995420000000001 0 0.000499642 3.3 0.000499782 3.3 0.000499882 0 0.0005001420000000001 0 0.000500242 3.3 0.000500502 3.3 0.000500602 0 0.000501462 0 0.000501562 3.3 0.000502542 3.3 0.000502642 0 0.0005026620000000001 0 0.000502762 3.3 0.000502822 3.3 0.0005029219999999999 0 0.0005045820000000001 0 0.000504682 3.3 0.000504822 3.3 0.000504922 0 0.000506502 0 0.000506602 3.3 0.000506742 3.3 0.000506842 0 0.0005074620000000001 0 0.000507562 3.3 0.000507822 3.3 0.000507922 0 0.000507942 0 0.000508042 3.3 0.000508062 3.3 0.0005081619999999999 0 0.000508422 0 0.000508522 3.3 0.000508662 3.3 0.000508762 0 0.000509502 0 0.000509602 3.3 0.000509622 3.3 0.000509722 0 0.000510462 0 0.000510562 3.3 0.0005105820000000001 3.3 0.000510682 0 0.0005125020000000001 0 0.000512602 3.3 0.0005127420000000001 3.3 0.000512842 0 0.0005144220000000001 0 0.000514522 3.3 0.000514662 3.3 0.000514762 0 0.000514902 0 0.000515002 3.3 0.000515142 3.3 0.000515242 0 0.000515382 0 0.0005154819999999999 3.3 0.0005156220000000001 3.3 0.000515722 0 0.000515742 0 0.000515842 3.3 0.000516102 3.3 0.000516202 0 0.000516342 0 0.000516442 3.3 0.000516582 3.3 0.000516682 0 0.0005167020000000001 0 0.000516802 3.3 0.000516822 3.3 0.000516922 0 0.000516942 0 0.000517042 3.3 0.000517062 3.3 0.0005171619999999999 0 0.0005173020000000001 0 0.000517402 3.3 0.0005175420000000001 3.3 0.000517642 0 0.000518502 0 0.000518602 3.3 0.000518662 3.3 0.000518762 0 0.0005204220000000001 0 0.000520522 3.3 0.0005206620000000001 3.3 0.000520762 0 0.0005223420000000001 0 0.000522442 3.3 0.0005229420000000001 3.3 0.000523042 0 0.000523302 0 0.000523402 3.3 0.000523542 3.3 0.0005236419999999999 0 0.000523902 0 0.000524002 3.3 0.0005242620000000001 3.3 0.000524362 0 0.000525222 0 0.0005253219999999999 3.3 0.0005263020000000001 3.3 0.000526402 0 0.000526422 0 0.000526522 3.3 0.000526582 3.3 0.000526682 0 0.000528342 0 0.000528442 3.3 0.000528582 3.3 0.0005286819999999999 0 0.0005302620000000001 0 0.000530362 3.3 0.0005305020000000001 3.3 0.000530602 0 0.000531222 0 0.000531322 3.3 0.0005315820000000001 3.3 0.000531682 0 0.000531702 0 0.000531802 3.3 0.000531822 3.3 0.000531922 0 0.0005321820000000001 0 0.000532282 3.3 0.0005324220000000001 3.3 0.000532522 0 0.0005332620000000001 0 0.000533362 3.3 0.000533382 3.3 0.0005334819999999999 0 0.000534222 0 0.0005343219999999999 3.3 0.000534342 3.3 0.000534442 0 0.000536262 0 0.000536362 3.3 0.000536502 3.3 0.000536602 0 0.000538182 0 0.000538282 3.3 0.000538422 3.3 0.0005385219999999999 0 0.0005386620000000001 0 0.000538762 3.3 0.0005389020000000001 3.3 0.000539002 0 0.000539142 0 0.000539242 3.3 0.000539382 3.3 0.000539482 0 0.0005395020000000001 0 0.000539602 3.3 0.000539862 3.3 0.000539962 0 0.0005401020000000001 0 0.000540202 3.3 0.0005403420000000001 3.3 0.000540442 0 0.000540462 0 0.000540562 3.3 0.0005405820000000001 3.3 0.000540682 0 0.000540702 0 0.000540802 3.3 0.000540822 3.3 0.000540922 0 0.000541062 0 0.000541162 3.3 0.000541302 3.3 0.000541402 0 0.0005422620000000001 0 0.000542362 3.3 0.0005424220000000001 3.3 0.000542522 0 0.000544182 0 0.000544282 3.3 0.000544422 3.3 0.000544522 0 0.000546102 0 0.000546202 3.3 0.000546702 3.3 0.000546802 0 0.0005470620000000001 0 0.000547162 3.3 0.000547302 3.3 0.000547402 0 0.0005476620000000001 0 0.000547762 3.3 0.000548022 3.3 0.000548122 0 0.000548982 0 0.000549082 3.3 0.000550062 3.3 0.000550162 0 0.0005501820000000001 0 0.000550282 3.3 0.000550342 3.3 0.0005504419999999999 0 0.0005521020000000001 0 0.000552202 3.3 0.000552342 3.3 0.000552442 0 0.000554022 0 0.000554122 3.3 0.000554262 3.3 0.000554362 0 0.0005549820000000001 0 0.000555082 3.3 0.000555342 3.3 0.000555442 0 0.0005554620000000001 0 0.000555562 3.3 0.000555582 3.3 0.0005556819999999999 0 0.000555942 0 0.000556042 3.3 0.000556182 3.3 0.000556282 0 0.000557022 0 0.000557122 3.3 0.000557142 3.3 0.000557242 0 0.000557982 0 0.000558082 3.3 0.000558102 3.3 0.0005582019999999999 0 0.0005600220000000001 0 0.000560122 3.3 0.0005602620000000001 3.3 0.000560362 0 0.0005619420000000001 0 0.000562042 3.3 0.000562182 3.3 0.000562282 0 0.000562422 0 0.000562522 3.3 0.000562662 3.3 0.000562762 0 0.000562902 0 0.000563002 3.3 0.0005631420000000001 3.3 0.000563242 0 0.000563262 0 0.000563362 3.3 0.0005636220000000001 3.3 0.000563722 0 0.000563862 0 0.000563962 3.3 0.000564102 3.3 0.000564202 0 0.0005642220000000001 0 0.000564322 3.3 0.000564342 3.3 0.000564442 0 0.0005644620000000001 0 0.000564562 3.3 0.000564582 3.3 0.0005646819999999999 0 0.0005648220000000001 0 0.000564922 3.3 0.0005650620000000001 3.3 0.000565162 0 0.000566022 0 0.000566122 3.3 0.000566182 3.3 0.000566282 0 0.000567942 0 0.0005680419999999999 3.3 0.0005681820000000001 3.3 0.000568282 0 0.0005698620000000001 0 0.000569962 3.3 0.000570462 3.3 0.0005705619999999999 0 0.000570822 0 0.000570922 3.3 0.000571062 3.3 0.000571162 0 0.000571422 0 0.000571522 3.3 0.0005717820000000001 3.3 0.000571882 0 0.000572742 0 0.000572842 3.3 0.0005738220000000001 3.3 0.000573922 0 0.000573942 0 0.000574042 3.3 0.000574102 3.3 0.000574202 0 0.000575862 0 0.000575962 3.3 0.000576102 3.3 0.0005762019999999999 0 0.000577782 0 0.0005778819999999999 3.3 0.0005780220000000001 3.3 0.000578122 0 0.000578742 0 0.000578842 3.3 0.0005791020000000001 3.3 0.000579202 0 0.000579222 0 0.000579322 3.3 0.000579342 3.3 0.000579442 0 0.0005797020000000001 0 0.000579802 3.3 0.0005799420000000001 3.3 0.000580042 0 0.0005807820000000001 0 0.000580882 3.3 0.000580902 3.3 0.000581002 0 0.000581742 0 0.000581842 3.3 0.000581862 3.3 0.000581962 0 0.000583782 0 0.000583882 3.3 0.000584022 3.3 0.000584122 0 0.000585702 0 0.000585802 3.3 0.000585942 3.3 0.0005860419999999999 0 0.0005861820000000001 0 0.000586282 3.3 0.0005864220000000001 3.3 0.000586522 0 0.0005866620000000001 0 0.000586762 3.3 0.000586902 3.3 0.000587002 0 0.0005870220000000001 0 0.000587122 3.3 0.000587382 3.3 0.000587482 0 0.000587622 0 0.0005877219999999999 3.3 0.0005878620000000001 3.3 0.000587962 0 0.000587982 0 0.000588082 3.3 0.0005881020000000001 3.3 0.000588202 0 0.000588222 0 0.000588322 3.3 0.000588342 3.3 0.000588442 0 0.000588582 0 0.000588682 3.3 0.000588822 3.3 0.000588922 0 0.0005897820000000001 0 0.000589882 3.3 0.0005899420000000001 3.3 0.000590042 0 0.000591702 0 0.000591802 3.3 0.000591942 3.3 0.000592042 0 0.000593622 0 0.000593722 3.3 0.000594222 3.3 0.000594322 0 0.0005945820000000001 0 0.000594682 3.3 0.0005948220000000001 3.3 0.000594922 0 0.0005951820000000001 0 0.000595282 3.3 0.000595542 3.3 0.000595642 0 0.0005965020000000001 0 0.000596602 3.3 0.000597582 3.3 0.000597682 0 0.0005977020000000001 0 0.000597802 3.3 0.000597862 3.3 0.000597962 0 0.0005996220000000001 0 0.000599722 3.3 0.000599862 3.3 0.000599962 0 0.000601542 0 0.000601642 3.3 0.000601782 3.3 0.000601882 0 0.000602502 0 0.0006026019999999999 3.3 0.000602862 3.3 0.000602962 0 0.0006029820000000001 0 0.000603082 3.3 0.000603102 3.3 0.000603202 0 0.000603462 0 0.000603562 3.3 0.000603702 3.3 0.000603802 0 0.000604542 0 0.000604642 3.3 0.0006046620000000001 3.3 0.000604762 0 0.0006055020000000001 0 0.000605602 3.3 0.000605622 3.3 0.0006057219999999999 0 0.0006075420000000001 0 0.000607642 3.3 0.0006077820000000001 3.3 0.000607882 0 0.0006094620000000001 0 0.000609562 3.3 0.000609702 3.3 0.000609802 0 0.000609942 0 0.000610042 3.3 0.000610182 3.3 0.000610282 0 0.000610422 0 0.000610522 3.3 0.000610662 3.3 0.0006107619999999999 0 0.000610782 0 0.000610882 3.3 0.0006111420000000001 3.3 0.000611242 0 0.000611382 0 0.000611482 3.3 0.000611622 3.3 0.000611722 0 0.0006117420000000001 0 0.000611842 3.3 0.000611862 3.3 0.000611962 0 0.0006119820000000001 0 0.000612082 3.3 0.000612102 3.3 0.000612202 0 0.000612342 0 0.0006124419999999999 3.3 0.0006125820000000001 3.3 0.000612682 0 0.000613542 0 0.000613642 3.3 0.000613702 3.3 0.000613802 0 0.000615462 0 0.0006155619999999999 3.3 0.0006157020000000001 3.3 0.000615802 0 0.0006173820000000001 0 0.000617482 3.3 0.000617982 3.3 0.0006180819999999999 0 0.000618342 0 0.000618442 3.3 0.000618582 3.3 0.000618682 0 0.000618942 0 0.000619042 3.3 0.0006193020000000001 3.3 0.000619402 0 0.000620262 0 0.000620362 3.3 0.000621342 3.3 0.0006214419999999999 0 0.000621462 0 0.000621562 3.3 0.0006216220000000001 3.3 0.000621722 0 0.000623382 0 0.000623482 3.3 0.000623622 3.3 0.000623722 0 0.000625302 0 0.000625402 3.3 0.0006255420000000001 3.3 0.000625642 0 0.000626262 0 0.000626362 3.3 0.0006266220000000001 3.3 0.000626722 0 0.000626742 0 0.000626842 3.3 0.0006268620000000001 3.3 0.000626962 0 0.0006272220000000001 0 0.000627322 3.3 0.0006274620000000001 3.3 0.000627562 0 0.0006283020000000001 0 0.000628402 3.3 0.000628422 3.3 0.000628522 0 0.000629262 0 0.000629362 3.3 0.000629382 3.3 0.000629482 0 0.000631302 0 0.000631402 3.3 0.000631542 3.3 0.000631642 0 0.000633222 0 0.000633322 3.3 0.000633462 3.3 0.000633562 0 0.000633702 0 0.0006338019999999999 3.3 0.0006339420000000001 3.3 0.000634042 0 0.0006341820000000001 0 0.000634282 3.3 0.000634422 3.3 0.000634522 0 0.0006345420000000001 0 0.000634642 3.3 0.000634902 3.3 0.000635002 0 0.000635142 0 0.000635242 3.3 0.0006353820000000001 3.3 0.000635482 0 0.000635502 0 0.000635602 3.3 0.0006356220000000001 3.3 0.000635722 0 0.000635742 0 0.000635842 3.3 0.0006358620000000001 3.3 0.000635962 0 0.000636102 0 0.000636202 3.3 0.000636342 3.3 0.000636442 0 0.0006373020000000001 0 0.000637402 3.3 0.000637462 3.3 0.0006375619999999999 0 0.000639222 0 0.000639322 3.3 0.000639462 3.3 0.000639562 0 0.000641142 0 0.000641242 3.3 0.000641742 3.3 0.000641842 0 0.0006421020000000001 0 0.000642202 3.3 0.0006423420000000001 3.3 0.000642442 0 0.000642702 0 0.0006428019999999999 3.3 0.000643062 3.3 0.000643162 0 0.0006440220000000001 0 0.000644122 3.3 0.000645102 3.3 0.000645202 0 0.0006452220000000001 0 0.000645322 3.3 0.000645382 3.3 0.000645482 0 0.0006471420000000001 0 0.000647242 3.3 0.0006473820000000001 3.3 0.000647482 0 0.0006490620000000001 0 0.000649162 3.3 0.000649302 3.3 0.000649402 0 0.000650022 0 0.0006501219999999999 3.3 0.000650382 3.3 0.000650482 0 0.0006505020000000001 0 0.000650602 3.3 0.000650622 3.3 0.000650722 0 0.000650982 0 0.000651082 3.3 0.000651222 3.3 0.000651322 0 0.000652062 0 0.000652162 3.3 0.0006521820000000001 3.3 0.000652282 0 0.0006530220000000001 0 0.000653122 3.3 0.000653142 3.3 0.000653242 0 0.0006550620000000001 0 0.000655162 3.3 0.0006553020000000001 3.3 0.000655402 0 0.0006569820000000001 0 0.000657082 3.3 0.0006572220000000001 3.3 0.000657322 0 0.000657462 0 0.000657562 3.3 0.000657702 3.3 0.000657802 0 0.000657942 0 0.000658042 3.3 0.000658182 3.3 0.0006582819999999999 0 0.000658302 0 0.000658402 3.3 0.0006586620000000001 3.3 0.000658762 0 0.0006589020000000001 0 0.000659002 3.3 0.000659142 3.3 0.000659242 0 0.0006592620000000001 0 0.000659362 3.3 0.000659382 3.3 0.000659482 0 0.0006595020000000001 0 0.000659602 3.3 0.000659622 3.3 0.000659722 0 0.000659862 0 0.0006599619999999999 3.3 0.0006601020000000001 3.3 0.000660202 0 0.000661062 0 0.000661162 3.3 0.000661222 3.3 0.000661322 0 0.000662982 0 0.000663082 3.3 0.000663222 3.3 0.0006633219999999999 0 0.000664902 0 0.0006650019999999999 3.3 0.000665502 3.3 0.000665602 0 0.000665862 0 0.000665962 3.3 0.000666102 3.3 0.000666202 0 0.000666462 0 0.000666562 3.3 0.0006668220000000001 3.3 0.000666922 0 0.000667782 0 0.000667882 3.3 0.000668862 3.3 0.0006689619999999999 0 0.000668982 0 0.000669082 3.3 0.0006691420000000001 3.3 0.000669242 0 0.000670902 0 0.000671002 3.3 0.000671142 3.3 0.000671242 0 0.000672822 0 0.000672922 3.3 0.000673062 3.3 0.0006731619999999999 0 0.000673782 0 0.000673882 3.3 0.0006741420000000001 3.3 0.000674242 0 0.000674262 0 0.000674362 3.3 0.0006743820000000001 3.3 0.000674482 0 0.000674742 0 0.0006748419999999999 3.3 0.0006749820000000001 3.3 0.000675082 0 0.0006758220000000001 0 0.000675922 3.3 0.000675942 3.3 0.000676042 0 0.000676782 0 0.000676882 3.3 0.0006769020000000001 3.3 0.000677002 0 0.000678822 0 0.000678922 3.3 0.000679062 3.3 0.000679162 0 0.000680742 0 0.000680842 3.3 0.000680982 3.3 0.000681082 0 0.000681222 0 0.0006813219999999999 3.3 0.0006814620000000001 3.3 0.000681562 0 0.0006817020000000001 0 0.000681802 3.3 0.000681942 3.3 0.000682042 0 0.000682062 0 0.0006821619999999999 3.3 0.000682422 3.3 0.000682522 0 0.000682662 0 0.000682762 3.3 0.000682902 3.3 0.0006830019999999999 0 0.000683022 0 0.000683122 3.3 0.0006831420000000001 3.3 0.000683242 0 0.000683262 0 0.000683362 3.3 0.0006833820000000001 3.3 0.000683482 0 0.000683622 0 0.000683722 3.3 0.000683862 3.3 0.000683962 0 0.0006848220000000001 0 0.000684922 3.3 0.000684982 3.3 0.0006850819999999999 0 0.0006867420000000001 0 0.000686842 3.3 0.000686982 3.3 0.000687082 0 0.000688662 0 0.000688762 3.3 0.0006892620000000001 3.3 0.000689362 0 0.0006896220000000001 0 0.000689722 3.3 0.0006898620000000001 3.3 0.000689962 0 0.000690222 0 0.0006903219999999999 3.3 0.000690582 3.3 0.000690682 0 0.0006915420000000001 0 0.000691642 3.3 0.000692622 3.3 0.000692722 0 0.000692742 0 0.0006928419999999999 3.3 0.000692902 3.3 0.000693002 0 0.0006946620000000001 0 0.000694762 3.3 0.0006949020000000001 3.3 0.000695002 0 0.0006965820000000001 0 0.000696682 3.3 0.000696822 3.3 0.000696922 0 0.000697542 0 0.0006976419999999999 3.3 0.000697902 3.3 0.000698002 0 0.0006980220000000001 0 0.000698122 3.3 0.000698142 3.3 0.000698242 0 0.000698502 0 0.000698602 3.3 0.000698742 3.3 0.000698842 0 0.000699582 0 0.000699682 3.3 0.0006997020000000001 3.3 0.000699802 0 0.0007005420000000001 0 0.000700642 3.3 0.000700662 3.3 0.000700762 0 0.000702582 0 0.0007026819999999999 3.3 0.0007028220000000001 3.3 0.000702922 0 0.0007045020000000001 0 0.000704602 3.3 0.0007047420000000001 3.3 0.000704842 0 0.000704982 0 0.000705082 3.3 0.000705222 3.3 0.000705322 0 0.000705462 0 0.000705562 3.3 0.000705702 3.3 0.000705802 0 0.000705822 0 0.000705922 3.3 0.0007061820000000001 3.3 0.000706282 0 0.0007064220000000001 0 0.000706522 3.3 0.000706662 3.3 0.000706762 0 0.0007067820000000001 0 0.000706882 3.3 0.000706902 3.3 0.000707002 0 0.0007070220000000001 0 0.000707122 3.3 0.000707142 3.3 0.000707242 0 0.000707382 0 0.000707482 3.3 0.0007076220000000001 3.3 0.000707722 0 0.000708582 0 0.000708682 3.3 0.000708742 3.3 0.000708842 0 0.000710502 0 0.000710602 3.3 0.000710742 3.3 0.0007108419999999999 0 0.000712422 0 0.0007125219999999999 3.3 0.000713022 3.3 0.000713122 0 0.000713382 0 0.000713482 3.3 0.000713622 3.3 0.000713722 0 0.000713982 0 0.000714082 3.3 0.0007143420000000001 3.3 0.000714442 0 0.000715302 0 0.000715402 3.3 0.000716382 3.3 0.000716482 0 0.000716502 0 0.000716602 3.3 0.0007166620000000001 3.3 0.000716762 0 0.000718422 0 0.000718522 3.3 0.000718662 3.3 0.000718762 0 0.000720342 0 0.000720442 3.3 0.000720582 3.3 0.0007206819999999999 0 0.0007213020000000001 0 0.000721402 3.3 0.0007216620000000001 3.3 0.000721762 0 0.000721782 0 0.000721882 3.3 0.0007219020000000001 3.3 0.000722002 0 0.000722262 0 0.0007223619999999999 3.3 0.0007225020000000001 3.3 0.000722602 0 0.0007233420000000001 0 0.000723442 3.3 0.000723462 3.3 0.000723562 0 0.000724302 0 0.000724402 3.3 0.0007244220000000001 3.3 0.000724522 0 0.000726342 0 0.000726442 3.3 0.000726582 3.3 0.000726682 0 0.000728262 0 0.000728362 3.3 0.000728502 3.3 0.000728602 0 0.000728742 0 0.0007288419999999999 3.3 0.0007289820000000001 3.3 0.000729082 0 0.0007292220000000001 0 0.000729322 3.3 0.0007294620000000001 3.3 0.000729562 0 0.000729582 0 0.0007296819999999999 3.3 0.000729942 3.3 0.000730042 0 0.000730182 0 0.000730282 3.3 0.000730422 3.3 0.0007305219999999999 0 0.000730542 0 0.000730642 3.3 0.0007306620000000001 3.3 0.000730762 0 0.000730782 0 0.000730882 3.3 0.0007309020000000001 3.3 0.000731002 0 0.0007311420000000001 0 0.000731242 3.3 0.000731382 3.3 0.000731482 0 0.0007323420000000001 0 0.000732442 3.3 0.000732502 3.3 0.000732602 0 0.0007342620000000001 0 0.000734362 3.3 0.000734502 3.3 0.000734602 0 0.000736182 0 0.000736282 3.3 0.0007367820000000001 3.3 0.000736882 0 0.000737142 0 0.0007372419999999999 3.3 0.0007373820000000001 3.3 0.000737482 0 0.000737742 0 0.000737842 3.3 0.000738102 3.3 0.000738202 0 0.0007390620000000001 0 0.000739162 3.3 0.0007401420000000001 3.3 0.000740242 0 0.000740262 0 0.0007403619999999999 3.3 0.000740422 3.3 0.000740522 0 0.0007421820000000001 0 0.000742282 3.3 0.0007424220000000001 3.3 0.000742522 0 0.0007441020000000001 0 0.000744202 3.3 0.000744342 3.3 0.000744442 0 0.000745062 0 0.000745162 3.3 0.000745422 3.3 0.000745522 0 0.0007455420000000001 0 0.000745642 3.3 0.000745662 3.3 0.000745762 0 0.000746022 0 0.000746122 3.3 0.000746262 3.3 0.000746362 0 0.000747102 0 0.000747202 3.3 0.0007472220000000001 3.3 0.000747322 0 0.0007480620000000001 0 0.000748162 3.3 0.000748182 3.3 0.000748282 0 0.000750102 0 0.0007502019999999999 3.3 0.0007503420000000001 3.3 0.000750442 0 0.0007520220000000001 0 0.000752122 3.3 0.0007522620000000001 3.3 0.000752362 0 0.000752502 0 0.000752602 3.3 0.000752742 3.3 0.000752842 0 0.000752982 0 0.000753082 3.3 0.000753222 3.3 0.000753322 0 0.000753342 0 0.000753442 3.3 0.0007537020000000001 3.3 0.000753802 0 0.0007539420000000001 0 0.000754042 3.3 0.000754182 3.3 0.000754282 0 0.000754302 0 0.0007544019999999999 3.3 0.000754422 3.3 0.000754522 0 0.0007545420000000001 0 0.000754642 3.3 0.000754662 3.3 0.000754762 0 0.000754902 0 0.000755002 3.3 0.000755142 3.3 0.0007552419999999999 0 0.000756102 0 0.000756202 3.3 0.0007562620000000001 3.3 0.000756362 0 0.000758022 0 0.000758122 3.3 0.000758262 3.3 0.000758362 0 0.000759942 0 0.0007600419999999999 3.3 0.000760542 3.3 0.000760642 0 0.000760902 0 0.000761002 3.3 0.000761142 3.3 0.000761242 0 0.0007615020000000001 0 0.000761602 3.3 0.0007618620000000001 3.3 0.000761962 0 0.000762822 0 0.000762922 3.3 0.000763902 3.3 0.000764002 0 0.000764022 0 0.000764122 3.3 0.0007641820000000001 3.3 0.000764282 0 0.000765942 0 0.000766042 3.3 0.000766182 3.3 0.000766282 0 0.000767862 0 0.000767962 3.3 0.000768102 3.3 0.000768202 0 0.0007688220000000001 0 0.000768922 3.3 0.0007691820000000001 3.3 0.000769282 0 0.000769302 0 0.000769402 3.3 0.0007694220000000001 3.3 0.000769522 0 0.000769782 0 0.0007698819999999999 3.3 0.0007700220000000001 3.3 0.000770122 0 0.0007708620000000001 0 0.000770962 3.3 0.000770982 3.3 0.000771082 0 0.000771822 0 0.000771922 3.3 0.0007719420000000001 3.3 0.000772042 0 0.000773862 0 0.000773962 3.3 0.000774102 3.3 0.000774202 0 0.000775782 0 0.000775882 3.3 0.000776022 3.3 0.000776122 0 0.000776262 0 0.000776362 3.3 0.000776502 3.3 0.0007766019999999999 0 0.0007767420000000001 0 0.000776842 3.3 0.0007769820000000001 3.3 0.000777082 0 0.000777102 0 0.000777202 3.3 0.000777462 3.3 0.000777562 0 0.000777702 0 0.000777802 3.3 0.000777942 3.3 0.000778042 0 0.000778062 0 0.000778162 3.3 0.000778182 3.3 0.0007782819999999999 0 0.000778302 0 0.000778402 3.3 0.0007784220000000001 3.3 0.000778522 0 0.0007786620000000001 0 0.000778762 3.3 0.000778902 3.3 0.000779002 0 0.0007798620000000001 0 0.000779962 3.3 0.000780022 3.3 0.000780122 0 0.0007817820000000001 0 0.000781882 3.3 0.0007820220000000001 3.3 0.000782122 0 0.000783702 0 0.000783802 3.3 0.0007843020000000001 3.3 0.000784402 0 0.000784662 0 0.0007847619999999999 3.3 0.0007849020000000001 3.3 0.000785002 0 0.000785262 0 0.000785362 3.3 0.000785622 3.3 0.000785722 0 0.0007865820000000001 0 0.000786682 3.3 0.0007876620000000001 3.3 0.000787762 0 0.000787782 0 0.000787882 3.3 0.000787942 3.3 0.000788042 0 0.000789702 0 0.0007898019999999999 3.3 0.0007899420000000001 3.3 0.000790042 0 0.0007916220000000001 0 0.000791722 3.3 0.0007918620000000001 3.3 0.000791962 0 0.000792582 0 0.000792682 3.3 0.000792942 3.3 0.000793042 0 0.0007930620000000001 0 0.000793162 3.3 0.000793182 3.3 0.000793282 0 0.000793542 0 0.000793642 3.3 0.000793782 3.3 0.000793882 0 0.000794622 0 0.000794722 3.3 0.0007947420000000001 3.3 0.000794842 0 0.0007955820000000001 0 0.000795682 3.3 0.000795702 3.3 0.000795802 0 0.000797622 0 0.000797722 3.3 0.000797862 3.3 0.0007979619999999999 0 0.000799542 0 0.0007996419999999999 3.3 0.0007997820000000001 3.3 0.000799882 0 0.0008000220000000001 0 0.000800122 3.3 0.000800262 3.3 0.000800362 0 0.000800502 0 0.000800602 3.3 0.000800742 3.3 0.000800842 0 0.0008008620000000001 0 0.000800962 3.3 0.0008012220000000001 3.3 0.000801322 0 0.0008014620000000001 0 0.000801562 3.3 0.0008017020000000001 3.3 0.000801802 0 0.000801822 0 0.0008019219999999999 3.3 0.000801942 3.3 0.000802042 0 0.0008020620000000001 0 0.000802162 3.3 0.000802182 3.3 0.000802282 0 0.000802422 0 0.000802522 3.3 0.000802662 3.3 0.0008027619999999999 0 0.000803622 0 0.000803722 3.3 0.0008037820000000001 3.3 0.000803882 0 0.000805542 0 0.000805642 3.3 0.000805782 3.3 0.000805882 0 0.000807462 0 0.000807562 3.3 0.000808062 3.3 0.000808162 0 0.000808422 0 0.000808522 3.3 0.000808662 3.3 0.000808762 0 0.0008090220000000001 0 0.000809122 3.3 0.000809382 3.3 0.0008094819999999999 0 0.000810342 0 0.000810442 3.3 0.000811422 3.3 0.000811522 0 0.0008115420000000001 0 0.000811642 3.3 0.0008117020000000001 3.3 0.000811802 0 0.000813462 0 0.000813562 3.3 0.000813702 3.3 0.000813802 0 0.000815382 0 0.000815482 3.3 0.000815622 3.3 0.000815722 0 0.0008163420000000001 0 0.000816442 3.3 0.000816702 3.3 0.0008168019999999999 0 0.000816822 0 0.000816922 3.3 0.0008169420000000001 3.3 0.000817042 0 0.000817302 0 0.000817402 3.3 0.000817542 3.3 0.0008176419999999999 0 0.000818382 0 0.0008184819999999999 3.3 0.000818502 3.3 0.000818602 0 0.000819342 0 0.000819442 3.3 0.0008194620000000001 3.3 0.000819562 0 0.0008213820000000001 0 0.000821482 3.3 0.000821622 3.3 0.000821722 0 0.000823302 0 0.000823402 3.3 0.000823542 3.3 0.000823642 0 0.000823782 0 0.000823882 3.3 0.000824022 3.3 0.0008241219999999999 0 0.0008242620000000001 0 0.000824362 3.3 0.0008245020000000001 3.3 0.000824602 0 0.000824622 0 0.000824722 3.3 0.000824982 3.3 0.000825082 0 0.000825222 0 0.000825322 3.3 0.000825462 3.3 0.000825562 0 0.000825582 0 0.000825682 3.3 0.000825702 3.3 0.0008258019999999999 0 0.000825822 0 0.000825922 3.3 0.0008259420000000001 3.3 0.000826042 0 0.0008261820000000001 0 0.000826282 3.3 0.000826422 3.3 0.000826522 0 0.000827382 0 0.0008274819999999999 3.3 0.000827542 3.3 0.000827642 0 0.0008293020000000001 0 0.000829402 3.3 0.0008295420000000001 3.3 0.000829642 0 0.0008312220000000001 0 0.000831322 3.3 0.0008318220000000001 3.3 0.000831922 0 0.000832182 0 0.0008322819999999999 3.3 0.0008324220000000001 3.3 0.000832522 0 0.000832782 0 0.000832882 3.3 0.000833142 3.3 0.000833242 0 0.0008341020000000001 0 0.000834202 3.3 0.0008351820000000001 3.3 0.000835282 0 0.000835302 0 0.000835402 3.3 0.000835462 3.3 0.000835562 0 0.000837222 0 0.0008373219999999999 3.3 0.0008374620000000001 3.3 0.000837562 0 0.0008391420000000001 0 0.000839242 3.3 0.0008393820000000001 3.3 0.000839482 0 0.000840102 0 0.000840202 3.3 0.000840462 3.3 0.000840562 0 0.000840582 0 0.0008406819999999999 3.3 0.000840702 3.3 0.000840802 0 0.0008410620000000001 0 0.000841162 3.3 0.000841302 3.3 0.000841402 0 0.000842142 0 0.000842242 3.3 0.0008422620000000001 3.3 0.000842362 0 0.0008431020000000001 0 0.000843202 3.3 0.000843222 3.3 0.000843322 0 0.000845142 0 0.000845242 3.3 0.000845382 3.3 0.0008454819999999999 0 0.000847062 0 0.0008471619999999999 3.3 0.0008473020000000001 3.3 0.000847402 0 0.0008475420000000001 0 0.000847642 3.3 0.000847782 3.3 0.000847882 0 0.000848022 0 0.000848122 3.3 0.000848262 3.3 0.000848362 0 0.0008483820000000001 0 0.000848482 3.3 0.000848742 3.3 0.0008488419999999999 0 0.0008489820000000001 0 0.000849082 3.3 0.0008492220000000001 3.3 0.000849322 0 0.000849342 0 0.000849442 3.3 0.000849462 3.3 0.000849562 0 0.000849582 0 0.0008496819999999999 3.3 0.000849702 3.3 0.000849802 0 0.000849942 0 0.000850042 3.3 0.000850182 3.3 0.000850282 0 0.000851142 0 0.000851242 3.3 0.0008513020000000001 3.3 0.000851402 0 0.000853062 0 0.000853162 3.3 0.000853302 3.3 0.000853402 0 0.000854982 0 0.000855082 3.3 0.000855582 3.3 0.000855682 0 0.000855942 0 0.000856042 3.3 0.000856182 3.3 0.000856282 0 0.0008565420000000001 0 0.000856642 3.3 0.000856902 3.3 0.0008570019999999999 0 0.000857862 0 0.000857962 3.3 0.000858942 3.3 0.000859042 0 0.0008590620000000001 0 0.000859162 3.3 0.000859222 3.3 0.0008593219999999999 0 0.000860982 0 0.000861082 3.3 0.000861222 3.3 0.000861322 0 0.000862902 0 0.000863002 3.3 0.000863142 3.3 0.000863242 0 0.0008638620000000001 0 0.000863962 3.3 0.000864222 3.3 0.0008643219999999999 0 0.000864342 0 0.000864442 3.3 0.0008644620000000001 3.3 0.000864562 0 0.000864822 0 0.000864922 3.3 0.000865062 3.3 0.0008651619999999999 0 0.000865902 0 0.0008660019999999999 3.3 0.000866022 3.3 0.000866122 0 0.000866862 0 0.000866962 3.3 0.0008669820000000001 3.3 0.000867082 0 0.0008689020000000001 0 0.000869002 3.3 0.000869142 3.3 0.000869242 0 0.000870822 0 0.000870922 3.3 0.000871062 3.3 0.000871162 0 0.000871302 0 0.000871402 3.3 0.000871542 3.3 0.000871642 0 0.000871782 0 0.0008718819999999999 3.3 0.0008720220000000001 3.3 0.000872122 0 0.000872142 0 0.000872242 3.3 0.000872502 3.3 0.000872602 0 0.000872742 0 0.000872842 3.3 0.000872982 3.3 0.000873082 0 0.0008731020000000001 0 0.000873202 3.3 0.000873222 3.3 0.0008733219999999999 0 0.000873342 0 0.000873442 3.3 0.0008734620000000001 3.3 0.000873562 0 0.0008737020000000001 0 0.000873802 3.3 0.0008739420000000001 3.3 0.000874042 0 0.000874902 0 0.0008750019999999999 3.3 0.000875062 3.3 0.000875162 0 0.0008768220000000001 0 0.000876922 3.3 0.0008770620000000001 3.3 0.000877162 0 0.0008787420000000001 0 0.000878842 3.3 0.0008793420000000001 3.3 0.000879442 0 0.000879702 0 0.000879802 3.3 0.000879942 3.3 0.0008800419999999999 0 0.000880302 0 0.000880402 3.3 0.000880662 3.3 0.000880762 0 0.000881622 0 0.0008817219999999999 3.3 0.0008827020000000001 3.3 0.000882802 0 0.000882822 0 0.000882922 3.3 0.000882982 3.3 0.000883082 0 0.000884742 0 0.0008848419999999999 3.3 0.0008849820000000001 3.3 0.000885082 0 0.0008866620000000001 0 0.000886762 3.3 0.0008869020000000001 3.3 0.000887002 0 0.000887622 0 0.000887722 3.3 0.000887982 3.3 0.000888082 0 0.000888102 0 0.0008882019999999999 3.3 0.000888222 3.3 0.000888322 0 0.0008885820000000001 0 0.000888682 3.3 0.000888822 3.3 0.000888922 0 0.000889662 0 0.000889762 3.3 0.000889782 3.3 0.0008898819999999999 0 0.000890622 0 0.0008907219999999999 3.3 0.000890742 3.3 0.000890842 0 0.000892662 0 0.000892762 3.3 0.000892902 3.3 0.0008930019999999999 0 0.000894582 0 0.0008946819999999999 3.3 0.0008948220000000001 3.3 0.000894922 0 0.0008950620000000001 0 0.000895162 3.3 0.0008953020000000001 3.3 0.000895402 0 0.000895542 0 0.000895642 3.3 0.000895782 3.3 0.000895882 0 0.0008959020000000001 0 0.000896002 3.3 0.000896262 3.3 0.0008963619999999999 0 0.0008965020000000001 0 0.000896602 3.3 0.0008967420000000001 3.3 0.000896842 0 0.000896862 0 0.000896962 3.3 0.000896982 3.3 0.000897082 0 0.000897102 0 0.0008972019999999999 3.3 0.000897222 3.3 0.000897322 0 0.000897462 0 0.000897562 3.3 0.000897702 3.3 0.000897802 0 0.000898662 0 0.000898762 3.3 0.0008988220000000001 3.3 0.000898922 0 0.000900582 0 0.000900682 3.3 0.000900822 3.3 0.000900922 0 0.000902502 0 0.000902602 3.3 0.000903102 3.3 0.000903202 0 0.0009034620000000001 0 0.000903562 3.3 0.000903702 3.3 0.000903802 0 0.0009040620000000001 0 0.000904162 3.3 0.000904422 3.3 0.0009045219999999999 0 0.000905382 0 0.000905482 3.3 0.000906462 3.3 0.000906562 0 0.0009065820000000001 0 0.000906682 3.3 0.000906742 3.3 0.0009068419999999999 0 0.000908502 0 0.000908602 3.3 0.000908742 3.3 0.000908842 0 0.000910422 0 0.000910522 3.3 0.000910662 3.3 0.000910762 0 0.0009113820000000001 0 0.000911482 3.3 0.000911742 3.3 0.000911842 0 0.000911862 0 0.000911962 3.3 0.000911982 3.3 0.0009120819999999999 0 0.000912342 0 0.000912442 3.3 0.000912582 3.3 0.000912682 0 0.000913422 0 0.0009135219999999999 3.3 0.000913542 3.3 0.000913642 0 0.000914382 0 0.000914482 3.3 0.000914502 3.3 0.0009146019999999999 0 0.0009164220000000001 0 0.000916522 3.3 0.000916662 3.3 0.000916762 0 0.000918342 0 0.000918442 3.3 0.000918582 3.3 0.000918682 0 0.000918822 0 0.000918922 3.3 0.000919062 3.3 0.000919162 0 0.000919302 0 0.0009194019999999999 3.3 0.0009195420000000001 3.3 0.000919642 0 0.000919662 0 0.000919762 3.3 0.000920022 3.3 0.000920122 0 0.000920262 0 0.000920362 3.3 0.000920502 3.3 0.000920602 0 0.0009206220000000001 0 0.000920722 3.3 0.000920742 3.3 0.000920842 0 0.000920862 0 0.000920962 3.3 0.000920982 3.3 0.0009210819999999999 0 0.0009212220000000001 0 0.000921322 3.3 0.0009214620000000001 3.3 0.000921562 0 0.000922422 0 0.000922522 3.3 0.000922582 3.3 0.000922682 0 0.000924342 0 0.0009244419999999999 3.3 0.0009245820000000001 3.3 0.000924682 0 0.0009262620000000001 0 0.000926362 3.3 0.0009268620000000001 3.3 0.000926962 0 0.000927222 0 0.000927322 3.3 0.000927462 3.3 0.0009275619999999999 0 0.000927822 0 0.000927922 3.3 0.000928182 3.3 0.000928282 0 0.000929142 0 0.0009292419999999999 3.3 0.0009302220000000001 3.3 0.000930322 0 0.000930342 0 0.000930442 3.3 0.000930502 3.3 0.000930602 0 0.000932262 0 0.000932362 3.3 0.000932502 3.3 0.0009326019999999999 0 0.000934182 0 0.0009342819999999999 3.3 0.0009344220000000001 3.3 0.000934522 0 0.000935142 0 0.000935242 3.3 0.0009355020000000001 3.3 0.000935602 0 0.000935622 0 0.0009357219999999999 3.3 0.000935742 3.3 0.000935842 0 0.0009361020000000001 0 0.000936202 3.3 0.0009363420000000001 3.3 0.000936442 0 0.000937182 0 0.000937282 3.3 0.000937302 3.3 0.0009374019999999999 0 0.000938142 0 0.0009382419999999999 3.3 0.000938262 3.3 0.000938362 0 0.000940182 0 0.000940282 3.3 0.000940422 3.3 0.000940522 0 0.000942102 0 0.000942202 3.3 0.000942342 3.3 0.0009424419999999999 0 0.0009425820000000001 0 0.000942682 3.3 0.0009428220000000001 3.3 0.000942922 0 0.000943062 0 0.000943162 3.3 0.000943302 3.3 0.000943402 0 0.0009434220000000001 0 0.000943522 3.3 0.000943782 3.3 0.000943882 0 0.000944022 0 0.0009441219999999999 3.3 0.0009442620000000001 3.3 0.000944362 0 0.000944382 0 0.000944482 3.3 0.0009445020000000001 3.3 0.000944602 0 0.000944622 0 0.0009447219999999999 3.3 0.000944742 3.3 0.000944842 0 0.000944982 0 0.000945082 3.3 0.000945222 3.3 0.000945322 0 0.0009461820000000001 0 0.000946282 3.3 0.0009463420000000001 3.3 0.000946442 0 0.000948102 0 0.000948202 3.3 0.000948342 3.3 0.000948442 0 0.000950022 0 0.000950122 3.3 0.000950622 3.3 0.000950722 0 0.0009509820000000001 0 0.000951082 3.3 0.000951222 3.3 0.000951322 0 0.0009515820000000001 0 0.000951682 3.3 0.000951942 3.3 0.000952042 0 0.000952902 0 0.000953002 3.3 0.000953982 3.3 0.000954082 0 0.0009541020000000001 0 0.000954202 3.3 0.000954262 3.3 0.0009543619999999999 0 0.0009560220000000001 0 0.000956122 3.3 0.000956262 3.3 0.000956362 0 0.000957942 0 0.000958042 3.3 0.000958182 3.3 0.000958282 0 0.0009589020000000001 0 0.000959002 3.3 0.000959262 3.3 0.000959362 0 0.000959382 0 0.000959482 3.3 0.000959502 3.3 0.0009596019999999999 0 0.000959862 0 0.000959962 3.3 0.000960102 3.3 0.000960202 0 0.000960942 0 0.000961042 3.3 0.000961062 3.3 0.000961162 0 0.000961902 0 0.000962002 3.3 0.000962022 3.3 0.0009621219999999999 0 0.0009639420000000001 0 0.000964042 3.3 0.0009641820000000001 3.3 0.000964282 0 0.0009658620000000001 0 0.000965962 3.3 0.000966102 3.3 0.000966202 0 0.000966342 0 0.000966442 3.3 0.000966582 3.3 0.000966682 0 0.000966822 0 0.0009669219999999999 3.3 0.0009670620000000001 3.3 0.000967162 0 0.000967182 0 0.000967282 3.3 0.0009675420000000001 3.3 0.000967642 0 0.000967782 0 0.000967882 3.3 0.000968022 3.3 0.000968122 0 0.0009681420000000001 0 0.000968242 3.3 0.000968262 3.3 0.000968362 0 0.000968382 0 0.000968482 3.3 0.000968502 3.3 0.0009686019999999999 0 0.0009687420000000001 0 0.000968842 3.3 0.0009689820000000001 3.3 0.000969082 0 0.000969942 0 0.000970042 3.3 0.000970102 3.3 0.000970202 0 0.000971862 0 0.0009719619999999999 3.3 0.0009721020000000001 3.3 0.000972202 0 0.0009737820000000001 0 0.000973882 3.3 0.000974382 3.3 0.0009744819999999999 0 0.000974742 0 0.000974842 3.3 0.000974982 3.3 0.0009750819999999999 0 0.000975342 0 0.000975442 3.3 0.0009757020000000001 3.3 0.000975802 0 0.0009766619999999999 0 0.000976762 3.3 0.000977742 3.3 0.000977842 0 0.000977862 0 0.000977962 3.3 0.0009780219999999998 3.3 0.0009781219999999999 0 0.000979782 0 0.000979882 3.3 0.0009800219999999999 3.3 0.000980122 0 0.0009817019999999999 0 0.000981802 3.3 0.000981942 3.3 0.000982042 0 0.000982662 0 0.000982762 3.3 0.0009830219999999998 3.3 0.000983122 0 0.000983142 0 0.000983242 3.3 0.000983262 3.3 0.000983362 0 0.000983622 0 0.000983722 3.3 0.0009838619999999998 3.3 0.000983962 0 0.0009847019999999998 0 0.000984802 3.3 0.000984822 3.3 0.000984922 0 0.000985662 0 0.000985762 3.3 0.000985782 3.3 0.000985882 0 0.000987702 0 0.000987802 3.3 0.000987942 3.3 0.000988042 0 0.000989622 0 0.000989722 3.3 0.000989862 3.3 0.000989962 0 0.0009901019999999999 0 0.000990202 3.3 0.000990342 3.3 0.000990442 0 0.0009905819999999998 0 0.0009906819999999999 3.3 0.000990822 3.3 0.000990922 0 0.0009909419999999999 0 0.000991042 3.3 0.000991302 3.3 0.000991402 0 0.000991542 0 0.000991642 3.3 0.0009917819999999999 3.3 0.000991882 0 0.000991902 0 0.000992002 3.3 0.000992022 3.3 0.000992122 0 0.000992142 0 0.000992242 3.3 0.0009922619999999998 3.3 0.0009923619999999999 0 0.000992502 0 0.000992602 3.3 0.000992742 3.3 0.000992842 0 0.000993702 0 0.000993802 3.3 0.0009938619999999999 3.3 0.000993962 0 0.0009956219999999998 0 0.0009957219999999999 3.3 0.000995862 3.3 0.000995962 0 0.000997542 0 0.000997642 3.3 0.0009981419999999998 3.3 0.0009982419999999999 0 0.0009985019999999999 0 0.000998602 3.3 0.000998742 3.3 0.000998842 0 0.000999102 0 0.000999202 3.3 0.000999462 3.3 0.000999562 0 0.001000422 0 0.001000522 3.3 0.0010015019999999998 3.3 0.0010016019999999999 0 0.001001622 0 0.001001722 3.3 0.0010017819999999999 3.3 0.001001882 0 0.0010035419999999998 0 0.001003642 3.3 0.001003782 3.3 0.001003882 0 0.001005462 0 0.001005562 3.3 0.001005702 3.3 0.001005802 0 0.0010064219999999999 0 0.001006522 3.3 0.001006782 3.3 0.001006882 0 0.0010069019999999998 0 0.001007002 3.3 0.001007022 3.3 0.001007122 0 0.001007382 0 0.001007482 3.3 0.001007622 3.3 0.001007722 0 0.001008462 0 0.001008562 3.3 0.0010085819999999998 3.3 0.001008682 0 0.0010094219999999998 0 0.001009522 3.3 0.001009542 3.3 0.001009642 0 0.0010114619999999999 0 0.001011562 3.3 0.001011702 3.3 0.001011802 0 0.001013382 0 0.001013482 3.3 0.0010136219999999998 3.3 0.0010137219999999999 0 0.001013862 0 0.001013962 3.3 0.001014102 3.3 0.001014202 0 0.0010143419999999999 0 0.001014442 3.3 0.001014582 3.3 0.001014682 0 0.001014702 0 0.001014802 3.3 0.001015062 3.3 0.001015162 0 0.0010153019999999998 0 0.0010154019999999999 3.3 0.001015542 3.3 0.001015642 0 0.0010156619999999999 0 0.001015762 3.3 0.001015782 3.3 0.001015882 0 0.001015902 0 0.001016002 3.3 0.0010160219999999999 3.3 0.001016122 0 0.001016262 0 0.001016362 3.3 0.0010165019999999999 3.3 0.001016602 0 0.001017462 0 0.001017562 3.3 0.001017622 3.3 0.001017722 0 0.0010193819999999999 0 0.001019482 3.3 0.001019622 3.3 0.001019722 0 0.001021302 0 0.001021402 3.3 0.0010219019999999999 3.3 0.001022002 0 0.001022262 0 0.001022362 3.3 0.001022502 3.3 0.001022602 0 0.0010228619999999998 0 0.0010229619999999999 3.3 0.0010232219999999998 3.3 0.001023322 0 0.001024182 0 0.001024282 3.3 0.0010252619999999999 3.3 0.001025362 0 0.001025382 0 0.001025482 3.3 0.001025542 3.3 0.001025642 0 0.001027302 0 0.001027402 3.3 0.001027542 3.3 0.001027642 0 0.001029222 0 0.001029322 3.3 0.0010294619999999999 3.3 0.001029562 0 0.001030182 0 0.001030282 3.3 0.001030542 3.3 0.001030642 0 0.001030662 0 0.001030762 3.3 0.0010307819999999998 3.3 0.001030882 0 0.0010311419999999999 0 0.001031242 3.3 0.001031382 3.3 0.001031482 0 0.001032222 0 0.001032322 3.3 0.001032342 3.3 0.001032442 0 0.001033182 0 0.001033282 3.3 0.0010333019999999998 3.3 0.0010334019999999999 0 0.001035222 0 0.001035322 3.3 0.001035462 3.3 0.001035562 0 0.001037142 0 0.001037242 3.3 0.0010373819999999999 3.3 0.001037482 0 0.001037622 0 0.001037722 3.3 0.0010378619999999999 3.3 0.001037962 0 0.001038102 0 0.001038202 3.3 0.0010383419999999998 3.3 0.0010384419999999999 0 0.001038462 0 0.001038562 3.3 0.001038822 3.3 0.001038922 0 0.0010390619999999999 0 0.001039162 3.3 0.001039302 3.3 0.001039402 0 0.001039422 0 0.001039522 3.3 0.0010395419999999999 3.3 0.001039642 0 0.001039662 0 0.001039762 3.3 0.001039782 3.3 0.001039882 0 0.0010400219999999998 0 0.0010401219999999999 3.3 0.001040262 3.3 0.001040362 0 0.0010412219999999999 0 0.001041322 3.3 0.001041382 3.3 0.001041482 0 0.001043142 0 0.001043242 3.3 0.0010433819999999998 3.3 0.0010434819999999999 0 0.0010450619999999998 0 0.0010451619999999999 3.3 0.001045662 3.3 0.001045762 0 0.001046022 0 0.001046122 3.3 0.0010462619999999998 3.3 0.001046362 0 0.0010466219999999999 0 0.001046722 3.3 0.001046982 3.3 0.001047082 0 0.0010479419999999998 0 0.001048042 3.3 0.001049022 3.3 0.001049122 0 0.0010491419999999999 0 0.001049242 3.3 0.001049302 3.3 0.001049402 0 0.001051062 0 0.001051162 3.3 0.0010513019999999998 3.3 0.001051402 0 0.0010529819999999998 0 0.0010530819999999999 3.3 0.001053222 3.3 0.001053322 0 0.001053942 0 0.001054042 3.3 0.001054302 3.3 0.001054402 0 0.001054422 0 0.001054522 3.3 0.001054542 3.3 0.001054642 0 0.001054902 0 0.001055002 3.3 0.001055142 3.3 0.001055242 0 0.001055982 0 0.001056082 3.3 0.001056102 3.3 0.001056202 0 0.001056942 0 0.001057042 3.3 0.0010570619999999999 3.3 0.001057162 0 0.001058982 0 0.001059082 3.3 0.0010592219999999999 3.3 0.001059322 0 0.0010609019999999999 0 0.001061002 3.3 0.001061142 3.3 0.001061242 0 0.0010613819999999998 0 0.0010614819999999999 3.3 0.001061622 3.3 0.001061722 0 0.001061862 0 0.001061962 3.3 0.0010621019999999999 3.3 0.001062202 0 0.0010622219999999998 0 0.0010623219999999999 3.3 0.0010625819999999998 3.3 0.001062682 0 0.001062822 0 0.001062922 3.3 0.0010630619999999998 3.3 0.0010631619999999999 0 0.001063182 0 0.001063282 3.3 0.001063302 3.3 0.001063402 0 0.0010634219999999998 0 0.001063522 3.3 0.001063542 3.3 0.001063642 0 0.0010637819999999999 0 0.001063882 3.3 0.001064022 3.3 0.001064122 0 0.001064982 0 0.001065082 3.3 0.0010651419999999998 3.3 0.0010652419999999999 0 0.001066902 0 0.001067002 3.3 0.0010671419999999999 3.3 0.001067242 0 0.0010688219999999999 0 0.001068922 3.3 0.001069422 3.3 0.001069522 0 0.001069782 0 0.001069882 3.3 0.001070022 3.3 0.001070122 0 0.001070382 0 0.001070482 3.3 0.001070742 3.3 0.001070842 0 0.001071702 0 0.001071802 3.3 0.001072782 3.3 0.001072882 0 0.001072902 0 0.001073002 3.3 0.0010730619999999998 3.3 0.001073162 0 0.001074822 0 0.001074922 3.3 0.001075062 3.3 0.001075162 0 0.0010767419999999999 0 0.001076842 3.3 0.001076982 3.3 0.001077082 0 0.0010777019999999998 0 0.0010778019999999999 3.3 0.0010780619999999999 3.3 0.001078162 0 0.001078182 0 0.001078282 3.3 0.001078302 3.3 0.001078402 0 0.001078662 0 0.001078762 3.3 0.0010789019999999999 3.3 0.001079002 0 0.0010797419999999999 0 0.001079842 3.3 0.001079862 3.3 0.001079962 0 0.001080702 0 0.001080802 3.3 0.001080822 3.3 0.001080922 0 0.0010827419999999998 0 0.0010828419999999999 3.3 0.001082982 3.3 0.001083082 0 0.001084662 0 0.001084762 3.3 0.001084902 3.3 0.001085002 0 0.0010851419999999999 0 0.001085242 3.3 0.001085382 3.3 0.001085482 0 0.0010856219999999998 0 0.001085722 3.3 0.001085862 3.3 0.001085962 0 0.0010859819999999999 0 0.001086082 3.3 0.001086342 3.3 0.001086442 0 0.001086582 0 0.001086682 3.3 0.0010868219999999999 3.3 0.001086922 0 0.001086942 0 0.001087042 3.3 0.001087062 3.3 0.001087162 0 0.001087182 0 0.001087282 3.3 0.0010873019999999998 3.3 0.001087402 0 0.001087542 0 0.001087642 3.3 0.001087782 3.3 0.001087882 0 0.001088742 0 0.001088842 3.3 0.0010889019999999999 3.3 0.001089002 0 0.0010906619999999998 0 0.001090762 3.3 0.001090902 3.3 0.001091002 0 0.001092582 0 0.001092682 3.3 0.0010931819999999998 3.3 0.0010932819999999999 0 0.0010935419999999999 0 0.001093642 3.3 0.001093782 3.3 0.001093882 0 0.001094142 0 0.001094242 3.3 0.001094502 3.3 0.001094602 0 0.001095462 0 0.001095562 3.3 0.0010965419999999998 3.3 0.0010966419999999999 0 0.001096662 0 0.001096762 3.3 0.001096822 3.3 0.001096922 0 0.0010985819999999999 0 0.001098682 3.3 0.001098822 3.3 0.001098922 0 0.001100502 0 0.001100602 3.3 0.0011007419999999998 3.3 0.0011008419999999999 0 0.0011014619999999999 0 0.001101562 3.3 0.001101822 3.3 0.001101922 0 0.0011019419999999999 0 0.001102042 3.3 0.001102062 3.3 0.001102162 0 0.0011024219999999998 0 0.0011025219999999999 3.3 0.001102662 3.3 0.001102762 0 0.001103502 0 0.001103602 3.3 0.0011036219999999998 3.3 0.001103722 0 0.0011044619999999998 0 0.001104562 3.3 0.001104582 3.3 0.001104682 0 0.0011065019999999999 0 0.001106602 3.3 0.001106742 3.3 0.001106842 0 0.001108422 0 0.001108522 3.3 0.0011086619999999998 3.3 0.001108762 0 0.001108902 0 0.001109002 3.3 0.001109142 3.3 0.001109242 0 0.001109382 0 0.001109482 3.3 0.001109622 3.3 0.001109722 0 0.001109742 0 0.001109842 3.3 0.001110102 3.3 0.001110202 0 0.0011103419999999998 0 0.001110442 3.3 0.001110582 3.3 0.001110682 0 0.0011107019999999999 0 0.001110802 3.3 0.001110822 3.3 0.001110922 0 0.001110942 0 0.001111042 3.3 0.001111062 3.3 0.001111162 0 0.001111302 0 0.001111402 3.3 0.0011115419999999999 3.3 0.001111642 0 0.001112502 0 0.001112602 3.3 0.001112662 3.3 0.001112762 0 0.001114422 0 0.001114522 3.3 0.001114662 3.3 0.001114762 0 0.001116342 0 0.001116442 3.3 0.0011169419999999999 3.3 0.001117042 0 0.001117302 0 0.001117402 3.3 0.001117542 3.3 0.001117642 0 0.0011179019999999998 0 0.0011180019999999999 3.3 0.0011182619999999999 3.3 0.001118362 0 0.001119222 0 0.001119322 3.3 0.0011203019999999999 3.3 0.001120402 0 0.0011204219999999998 0 0.0011205219999999999 3.3 0.001120582 3.3 0.001120682 0 0.001122342 0 0.001122442 3.3 0.001122582 3.3 0.001122682 0 0.001124262 0 0.001124362 3.3 0.0011245019999999999 3.3 0.001124602 0 0.001125222 0 0.001125322 3.3 0.001125582 3.3 0.001125682 0 0.001125702 0 0.001125802 3.3 0.0011258219999999998 3.3 0.001125922 0 0.0011261819999999999 0 0.001126282 3.3 0.001126422 3.3 0.001126522 0 0.001127262 0 0.001127362 3.3 0.001127382 3.3 0.001127482 0 0.001128222 0 0.001128322 3.3 0.0011283419999999998 3.3 0.001128442 0 0.001130262 0 0.001130362 3.3 0.001130502 3.3 0.001130602 0 0.001132182 0 0.001132282 3.3 0.001132422 3.3 0.001132522 0 0.001132662 0 0.001132762 3.3 0.0011329019999999999 3.3 0.001133002 0 0.001133142 0 0.001133242 3.3 0.0011333819999999998 3.3 0.001133482 0 0.001133502 0 0.001133602 3.3 0.001133862 3.3 0.001133962 0 0.001134102 0 0.001134202 3.3 0.001134342 3.3 0.001134442 0 0.001134462 0 0.001134562 3.3 0.0011345819999999999 3.3 0.001134682 0 0.001134702 0 0.001134802 3.3 0.001134822 3.3 0.001134922 0 0.0011350619999999998 0 0.0011351619999999999 3.3 0.001135302 3.3 0.001135402 0 0.0011362619999999999 0 0.001136362 3.3 0.001136422 3.3 0.001136522 0 0.001138182 0 0.001138282 3.3 0.0011384219999999998 3.3 0.0011385219999999999 0 0.0011401019999999998 0 0.0011402019999999999 3.3 0.001140702 3.3 0.001140802 0 0.001141062 0 0.001141162 3.3 0.0011413019999999999 3.3 0.001141402 0 0.0011416619999999999 0 0.001141762 3.3 0.001142022 3.3 0.001142122 0 0.0011429819999999999 0 0.001143082 3.3 0.001144062 3.3 0.001144162 0 0.0011441819999999999 0 0.001144282 3.3 0.001144342 3.3 0.001144442 0 0.001146102 0 0.001146202 3.3 0.0011463419999999998 3.3 0.001146442 0 0.0011480219999999998 0 0.001148122 3.3 0.001148262 3.3 0.001148362 0 0.001148982 0 0.001149082 3.3 0.001149342 3.3 0.001149442 0 0.001149462 0 0.001149562 3.3 0.001149582 3.3 0.001149682 0 0.001149942 0 0.001150042 3.3 0.001150182 3.3 0.001150282 0 0.001151022 0 0.001151122 3.3 0.001151142 3.3 0.001151242 0 0.001151982 0 0.001152082 3.3 0.001152102 3.3 0.001152202 0 0.001154022 0 0.001154122 3.3 0.0011542619999999999 3.3 0.001154362 0 0.0011559419999999999 0 0.001156042 3.3 0.001156182 3.3 0.001156282 0 0.0011564219999999998 0 0.0011565219999999999 3.3 0.001156662 3.3 0.001156762 0 0.001156902 0 0.001157002 3.3 0.001157142 3.3 0.001157242 0 0.0011572619999999998 0 0.0011573619999999999 3.3 0.0011576219999999999 3.3 0.001157722 0 0.001157862 0 0.001157962 3.3 0.0011581019999999998 3.3 0.0011582019999999999 0 0.001158222 0 0.001158322 3.3 0.001158342 3.3 0.001158442 0 0.0011584619999999999 0 0.001158562 3.3 0.001158582 3.3 0.001158682 0 0.0011588219999999999 0 0.001158922 3.3 0.001159062 3.3 0.001159162 0 0.001160022 0 0.001160122 3.3 0.0011601819999999998 3.3 0.001160282 0 0.001161942 0 0.001162042 3.3 0.0011621819999999999 3.3 0.001162282 0 0.0011638619999999999 0 0.001163962 3.3 0.001164462 3.3 0.001164562 0 0.0011648219999999998 0 0.0011649219999999999 3.3 0.001165062 3.3 0.001165162 0 0.001165422 0 0.001165522 3.3 0.001165782 3.3 0.001165882 0 0.001166742 0 0.001166842 3.3 0.001167822 3.3 0.001167922 0 0.001167942 0 0.001168042 3.3 0.0011681019999999999 3.3 0.001168202 0 0.0011698619999999998 0 0.0011699619999999999 3.3 0.001170102 3.3 0.001170202 0 0.001171782 0 0.001171882 3.3 0.001172022 3.3 0.001172122 0 0.0011727419999999998 0 0.001172842 3.3 0.0011731019999999999 3.3 0.001173202 0 0.001173222 0 0.001173322 3.3 0.001173342 3.3 0.001173442 0 0.001173702 0 0.001173802 3.3 0.0011739419999999999 3.3 0.001174042 0 0.0011747819999999999 0 0.001174882 3.3 0.001174902 3.3 0.001175002 0 0.001175742 0 0.001175842 3.3 0.001175862 3.3 0.001175962 0 0.0011777819999999998 0 0.0011778819999999999 3.3 0.001178022 3.3 0.001178122 0 0.001179702 0 0.001179802 3.3 0.001179942 3.3 0.001180042 0 0.0011801819999999999 0 0.001180282 3.3 0.001180422 3.3 0.001180522 0 0.0011806619999999999 0 0.001180762 3.3 0.001180902 3.3 0.001181002 0 0.0011810219999999999 0 0.001181122 3.3 0.001181382 3.3 0.001181482 0 0.001181622 0 0.001181722 3.3 0.0011818619999999999 3.3 0.001181962 0 0.0011819819999999998 0 0.0011820819999999999 3.3 0.001182102 3.3 0.001182202 0 0.001182222 0 0.001182322 3.3 0.0011823419999999999 3.3 0.001182442 0 0.001182582 0 0.001182682 3.3 0.0011828219999999998 3.3 0.0011829219999999999 0 0.001183782 0 0.001183882 3.3 0.001183942 3.3 0.001184042 0 0.0011857019999999998 0 0.001185802 3.3 0.001185942 3.3 0.001186042 0 0.001187622 0 0.001187722 3.3 0.0011882219999999998 3.3 0.001188322 0 0.0011885819999999999 0 0.001188682 3.3 0.001188822 3.3 0.001188922 0 0.001189182 0 0.001189282 3.3 0.0011895419999999998 3.3 0.0011896419999999999 0 0.001190502 0 0.001190602 3.3 0.0011915819999999998 3.3 0.001191682 0 0.001191702 0 0.001191802 3.3 0.001191862 3.3 0.001191962 0 0.0011936219999999999 0 0.001193722 3.3 0.001193862 3.3 0.001193962 0 0.001195542 0 0.001195642 3.3 0.0011957819999999998 3.3 0.0011958819999999999 0 0.001196502 0 0.001196602 3.3 0.001196862 3.3 0.001196962 0 0.0011969819999999999 0 0.001197082 3.3 0.001197102 3.3 0.001197202 0 0.0011974619999999998 0 0.0011975619999999999 3.3 0.001197702 3.3 0.001197802 0 0.001198542 0 0.001198642 3.3 0.0011986619999999999 3.3 0.001198762 0 0.0011995019999999999 0 0.001199602 3.3 0.001199622 3.3 0.001199722 0 0.0012015419999999999 0 0.001201642 3.3 0.001201782 3.3 0.001201882 0 0.001203462 0 0.001203562 3.3 0.0012037019999999999 3.3 0.001203802 0 0.001203942 0 0.001204042 3.3 0.0012041819999999998 3.3 0.0012042819999999999 0 0.001204422 0 0.001204522 3.3 0.001204662 3.3 0.001204762 0 0.001204782 0 0.001204882 3.3 0.001205142 3.3 0.001205242 0 0.0012053819999999999 0 0.001205482 3.3 0.001205622 3.3 0.001205722 0 0.0012057419999999999 0 0.001205842 3.3 0.0012058619999999998 3.3 0.0012059619999999999 0 0.001205982 0 0.001206082 3.3 0.001206102 3.3 0.001206202 0 0.001206342 0 0.001206442 3.3 0.0012065819999999999 3.3 0.001206682 0 0.0012075419999999998 0 0.0012076419999999999 3.3 0.001207702 3.3 0.001207802 0 0.001209462 0 0.001209562 3.3 0.001209702 3.3 0.001209802 0 0.001211382 0 0.001211482 3.3 0.001211982 3.3 0.001212082 0 0.001212342 0 0.001212442 3.3 0.001212582 3.3 0.001212682 0 0.0012129419999999998 0 0.001213042 3.3 0.0012133019999999999 3.3 0.001213402 0 0.001214262 0 0.001214362 3.3 0.001215342 3.3 0.001215442 0 0.0012154619999999998 0 0.001215562 3.3 0.001215622 3.3 0.001215722 0 0.001217382 0 0.001217482 3.3 0.001217622 3.3 0.001217722 0 0.001219302 0 0.001219402 3.3 0.001219542 3.3 0.001219642 0 0.001220262 0 0.001220362 3.3 0.001220622 3.3 0.001220722 0 0.001220742 0 0.001220842 3.3 0.0012208619999999999 3.3 0.001220962 0 0.0012212219999999999 0 0.001221322 3.3 0.001221462 3.3 0.001221562 0 0.001222302 0 0.001222402 3.3 0.001222422 3.3 0.001222522 0 0.001223262 0 0.001223362 3.3 0.0012233819999999999 3.3 0.001223482 0 0.001225302 0 0.001225402 3.3 0.0012255419999999998 3.3 0.0012256419999999999 0 0.0012272219999999998 0 0.0012273219999999999 3.3 0.001227462 3.3 0.001227562 0 0.001227702 0 0.001227802 3.3 0.0012279419999999999 3.3 0.001228042 0 0.001228182 0 0.001228282 3.3 0.0012284219999999998 3.3 0.001228522 0 0.001228542 0 0.001228642 3.3 0.0012289019999999998 3.3 0.0012290019999999999 0 0.001229142 0 0.001229242 3.3 0.001229382 3.3 0.001229482 0 0.001229502 0 0.001229602 3.3 0.0012296219999999999 3.3 0.001229722 0 0.0012297419999999998 0 0.0012298419999999999 3.3 0.001229862 3.3 0.001229962 0 0.0012301019999999998 0 0.001230202 3.3 0.001230342 3.3 0.001230442 0 0.0012313019999999999 0 0.001231402 3.3 0.001231462 3.3 0.001231562 0 0.001233222 0 0.001233322 3.3 0.0012334619999999998 3.3 0.001233562 0 0.0012351419999999998 0 0.001235242 3.3 0.001235742 3.3 0.001235842 0 0.001236102 0 0.001236202 3.3 0.0012363419999999999 3.3 0.001236442 0 0.001236702 0 0.001236802 3.3 0.001237062 3.3 0.001237162 0 0.0012380219999999999 0 0.001238122 3.3 0.001239102 3.3 0.001239202 0 0.001239222 0 0.001239322 3.3 0.0012393819999999998 3.3 0.0012394819999999999 0 0.001241142 0 0.001241242 3.3 0.0012413819999999999 3.3 0.001241482 0 0.0012430619999999999 0 0.001243162 3.3 0.001243302 3.3 0.001243402 0 0.001244022 0 0.001244122 3.3 0.0012443819999999998 3.3 0.0012444819999999999 0 0.001244502 0 0.001244602 3.3 0.001244622 3.3 0.001244722 0 0.001244982 0 0.001245082 3.3 0.0012452219999999998 3.3 0.0012453219999999999 0 0.0012460619999999998 0 0.0012461619999999999 3.3 0.001246182 3.3 0.001246282 0 0.001247022 0 0.001247122 3.3 0.001247142 3.3 0.001247242 0 0.001249062 0 0.001249162 3.3 0.0012493019999999999 3.3 0.001249402 0 0.0012509819999999999 0 0.001251082 3.3 0.001251222 3.3 0.001251322 0 0.0012514619999999998 0 0.001251562 3.3 0.001251702 3.3 0.001251802 0 0.0012519419999999998 0 0.0012520419999999999 3.3 0.001252182 3.3 0.001252282 0 0.0012523019999999998 0 0.001252402 3.3 0.0012526619999999999 3.3 0.001252762 0 0.001252902 0 0.001253002 3.3 0.0012531419999999998 3.3 0.001253242 0 0.001253262 0 0.001253362 3.3 0.001253382 3.3 0.001253482 0 0.0012535019999999999 0 0.001253602 3.3 0.001253622 3.3 0.001253722 0 0.001253862 0 0.001253962 3.3 0.001254102 3.3 0.001254202 0 0.001255062 0 0.001255162 3.3 0.0012552219999999998 3.3 0.001255322 0 0.001256982 0 0.001257082 3.3 0.001257222 3.3 0.001257322 0 0.001258902 0 0.001259002 3.3 0.001259502 3.3 0.001259602 0 0.0012598619999999998 0 0.0012599619999999999 3.3 0.001260102 3.3 0.001260202 0 0.001260462 0 0.001260562 3.3 0.001260822 3.3 0.001260922 0 0.001261782 0 0.001261882 3.3 0.001262862 3.3 0.001262962 0 0.001262982 0 0.001263082 3.3 0.0012631419999999999 3.3 0.001263242 0 0.0012649019999999998 0 0.0012650019999999999 3.3 0.001265142 3.3 0.001265242 0 0.001266822 0 0.001266922 3.3 0.001267062 3.3 0.001267162 0 0.0012677819999999999 0 0.001267882 3.3 0.0012681419999999999 3.3 0.001268242 0 0.0012682619999999998 0 0.0012683619999999999 3.3 0.001268382 3.3 0.001268482 0 0.001268742 0 0.001268842 3.3 0.0012689819999999999 3.3 0.001269082 0 0.0012698219999999999 0 0.001269922 3.3 0.0012699419999999998 3.3 0.0012700419999999999 0 0.0012707819999999998 0 0.0012708819999999999 3.3 0.001270902 3.3 0.001271002 0 0.0012728219999999998 0 0.001272922 3.3 0.001273062 3.3 0.001273162 0 0.001274742 0 0.001274842 3.3 0.001274982 3.3 0.001275082 0 0.001275222 0 0.001275322 3.3 0.001275462 3.3 0.001275562 0 0.0012757019999999999 0 0.001275802 3.3 0.001275942 3.3 0.001276042 0 0.001276062 0 0.001276162 3.3 0.001276422 3.3 0.001276522 0 0.001276662 0 0.001276762 3.3 0.001276902 3.3 0.001277002 0 0.0012770219999999998 0 0.001277122 3.3 0.001277142 3.3 0.001277242 0 0.001277262 0 0.001277362 3.3 0.0012773819999999999 3.3 0.001277482 0 0.001277622 0 0.001277722 3.3 0.0012778619999999998 3.3 0.0012779619999999999 0 0.001278822 0 0.001278922 3.3 0.001278982 3.3 0.001279082 0 0.0012807419999999999 0 0.001280842 3.3 0.001280982 3.3 0.001281082 0 0.001282662 0 0.001282762 3.3 0.0012832619999999999 3.3 0.001283362 0 0.0012836219999999999 0 0.001283722 3.3 0.001283862 3.3 0.001283962 0 0.001284222 0 0.001284322 3.3 0.0012845819999999998 3.3 0.0012846819999999999 0 0.001285542 0 0.001285642 3.3 0.0012866219999999999 3.3 0.001286722 0 0.001286742 0 0.001286842 3.3 0.001286902 3.3 0.001287002 0 0.0012886619999999999 0 0.001288762 3.3 0.001288902 3.3 0.001289002 0 0.001290582 0 0.001290682 3.3 0.0012908219999999998 3.3 0.001290922 0 0.001291542 0 0.001291642 3.3 0.001291902 3.3 0.001292002 0 0.0012920219999999999 0 0.001292122 3.3 0.0012921419999999998 3.3 0.0012922419999999999 0 0.0012925019999999998 0 0.001292602 3.3 0.001292742 3.3 0.001292842 0 0.001293582 0 0.001293682 3.3 0.0012937019999999999 3.3 0.001293802 0 0.0012945419999999999 0 0.001294642 3.3 0.0012946619999999998 3.3 0.0012947619999999999 0 0.001296582 0 0.001296682 3.3 0.001296822 3.3 0.001296922 0 0.001298502 0 0.001298602 3.3 0.0012987419999999999 3.3 0.001298842 0 0.001298982 0 0.001299082 3.3 0.0012992219999999998 3.3 0.0012993219999999999 0 0.001299462 0 0.001299562 3.3 0.001299702 3.3 0.001299802 0 0.001299822 0 0.001299922 3.3 0.001300182 3.3 0.001300282 0 0.0013004219999999999 0 0.001300522 3.3 0.001300662 3.3 0.001300762 0 0.001300782 0 0.001300882 3.3 0.0013009019999999998 3.3 0.0013010019999999999 0 0.001301022 0 0.001301122 3.3 0.001301142 3.3 0.001301242 0 0.001301382 0 0.001301482 3.3 0.001301622 3.3 0.001301722 0 0.0013025819999999998 0 0.0013026819999999999 3.3 0.001302742 3.3 0.001302842 0 0.001304502 0 0.001304602 3.3 0.001304742 3.3 0.001304842 0 0.001306422 0 0.001306522 3.3 0.001307022 3.3 0.001307122 0 0.001307382 0 0.001307482 3.3 0.0013076219999999998 3.3 0.0013077219999999999 0 0.0013079819999999999 0 0.001308082 3.3 0.0013083419999999999 3.3 0.001308442 0 0.0013093019999999998 0 0.0013094019999999999 3.3 0.001310382 3.3 0.001310482 0 0.0013105019999999998 0 0.001310602 3.3 0.001310662 3.3 0.001310762 0 0.001312422 0 0.001312522 3.3 0.0013126619999999998 3.3 0.0013127619999999999 0 0.0013143419999999998 0 0.0013144419999999999 3.3 0.001314582 3.3 0.001314682 0 0.001315302 0 0.001315402 3.3 0.001315662 3.3 0.001315762 0 0.001315782 0 0.001315882 3.3 0.0013159019999999999 3.3 0.001316002 0 0.001316262 0 0.001316362 3.3 0.001316502 3.3 0.001316602 0 0.001317342 0 0.001317442 3.3 0.001317462 3.3 0.001317562 0 0.001318302 0 0.001318402 3.3 0.0013184219999999999 3.3 0.001318522 0 0.001320342 0 0.001320442 3.3 0.0013205819999999998 3.3 0.0013206819999999999 0 0.0013222619999999998 0 0.0013223619999999999 3.3 0.001322502 3.3 0.001322602 0 0.001322742 0 0.001322842 3.3 0.0013229819999999999 3.3 0.001323082 0 0.001323222 0 0.001323322 3.3 0.0013234619999999999 3.3 0.001323562 0 0.001323582 0 0.001323682 3.3 0.0013239419999999998 3.3 0.0013240419999999999 0 0.001324182 0 0.001324282 3.3 0.001324422 3.3 0.001324522 0 0.001324542 0 0.001324642 3.3 0.0013246619999999999 3.3 0.001324762 0 0.0013247819999999998 0 0.0013248819999999999 3.3 0.001324902 3.3 0.001325002 0 0.0013251419999999999 0 0.001325242 3.3 0.001325382 3.3 0.001325482 0 0.0013263419999999999 0 0.001326442 3.3 0.001326502 3.3 0.001326602 0 0.001328262 0 0.001328362 3.3 0.0013285019999999999 3.3 0.001328602 0 0.0013301819999999998 0 0.001330282 3.3 0.001330782 3.3 0.001330882 0 0.001331142 0 0.001331242 3.3 0.0013313819999999999 3.3 0.001331482 0 0.001331742 0 0.001331842 3.3 0.001332102 3.3 0.001332202 0 0.0013330619999999999 0 0.001333162 3.3 0.001334142 3.3 0.001334242 0 0.001334262 0 0.001334362 3.3 0.0013344219999999998 3.3 0.0013345219999999999 0 0.001336182 0 0.001336282 3.3 0.0013364219999999999 3.3 0.001336522 0 0.0013381019999999999 0 0.001338202 3.3 0.001338342 3.3 0.001338442 0 0.001339062 0 0.001339162 3.3 0.0013394219999999998 3.3 0.001339522 0 0.001339542 0 0.001339642 3.3 0.001339662 3.3 0.001339762 0 0.001340022 0 0.001340122 3.3 0.0013402619999999998 3.3 0.0013403619999999999 0 0.0013411019999999998 0 0.0013412019999999999 3.3 0.001341222 3.3 0.001341322 0 0.001342062 0 0.001342162 3.3 0.001342182 3.3 0.001342282 0 0.001344102 0 0.001344202 3.3 0.0013443419999999999 3.3 0.001344442 0 0.0013460219999999999 0 0.001346122 3.3 0.001346262 3.3 0.001346362 0 0.0013465019999999999 0 0.001346602 3.3 0.001346742 3.3 0.001346842 0 0.0013469819999999998 0 0.0013470819999999999 3.3 0.001347222 3.3 0.001347322 0 0.0013473419999999999 0 0.001347442 3.3 0.0013477019999999999 3.3 0.001347802 0 0.001347942 0 0.001348042 3.3 0.0013481819999999999 3.3 0.001348282 0 0.001348302 0 0.001348402 3.3 0.001348422 3.3 0.001348522 0 0.0013485419999999999 0 0.001348642 3.3 0.0013486619999999998 3.3 0.0013487619999999999 0 0.001348902 0 0.001349002 3.3 0.001349142 3.3 0.001349242 0 0.001350102 0 0.001350202 3.3 0.0013502619999999999 3.3 0.001350362 0 0.0013520219999999998 0 0.0013521219999999999 3.3 0.001352262 3.3 0.001352362 0 0.001353942 0 0.001354042 3.3 0.0013545419999999998 3.3 0.0013546419999999999 0 0.0013549019999999998 0 0.001355002 3.3 0.001355142 3.3 0.001355242 0 0.001355502 0 0.001355602 3.3 0.001355862 3.3 0.001355962 0 0.001356822 0 0.001356922 3.3 0.001357902 3.3 0.001358002 0 0.001358022 0 0.001358122 3.3 0.0013581819999999999 3.3 0.001358282 0 0.0013599419999999998 0 0.001360042 3.3 0.001360182 3.3 0.001360282 0 0.001361862 0 0.001361962 3.3 0.001362102 3.3 0.001362202 0 0.0013628219999999999 0 0.001362922 3.3 0.001363182 3.3 0.001363282 0 0.0013633019999999998 0 0.0013634019999999999 3.3 0.001363422 3.3 0.001363522 0 0.001363782 0 0.001363882 3.3 0.0013640219999999999 3.3 0.001364122 0 0.0013648619999999999 0 0.001364962 3.3 0.0013649819999999998 3.3 0.0013650819999999999 0 0.0013658219999999998 0 0.0013659219999999999 3.3 0.001365942 3.3 0.001366042 0 0.0013678619999999999 0 0.001367962 3.3 0.001368102 3.3 0.001368202 0 0.001369782 0 0.001369882 3.3 0.0013700219999999998 3.3 0.0013701219999999999 0 0.001370262 0 0.001370362 3.3 0.001370502 3.3 0.001370602 0 0.0013707419999999999 0 0.001370842 3.3 0.001370982 3.3 0.001371082 0 0.001371102 0 0.001371202 3.3 0.001371462 3.3 0.001371562 0 0.0013717019999999998 0 0.0013718019999999999 3.3 0.001371942 3.3 0.001372042 0 0.0013720619999999998 0 0.001372162 3.3 0.001372182 3.3 0.001372282 0 0.001372302 0 0.001372402 3.3 0.0013724219999999999 3.3 0.001372522 0 0.001372662 0 0.001372762 3.3 0.0013729019999999998 3.3 0.001373002 0 0.001373862 0 0.001373962 3.3 0.001374022 3.3 0.001374122 0 0.0013757819999999999 0 0.001375882 3.3 0.001376022 3.3 0.001376122 0 0.001377702 0 0.001377802 3.3 0.0013783019999999999 3.3 0.001378402 0 0.001378662 0 0.001378762 3.3 0.001378902 3.3 0.001379002 0 0.001379262 0 0.001379362 3.3 0.0013796219999999998 3.3 0.001379722 0 0.001380582 0 0.001380682 3.3 0.0013816619999999999 3.3 0.001381762 0 0.001381782 0 0.001381882 3.3 0.001381942 3.3 0.001382042 0 0.001383702 0 0.001383802 3.3 0.001383942 3.3 0.001384042 0 0.001385622 0 0.001385722 3.3 0.0013858619999999999 3.3 0.001385962 0 0.001386582 0 0.001386682 3.3 0.001386942 3.3 0.001387042 0 0.0013870619999999999 0 0.001387162 3.3 0.0013871819999999998 3.3 0.0013872819999999999 0 0.0013875419999999999 0 0.001387642 3.3 0.001387782 3.3 0.001387882 0 0.001388622 0 0.001388722 3.3 0.0013887419999999999 3.3 0.001388842 0 0.0013895819999999999 0 0.001389682 3.3 0.0013897019999999998 3.3 0.0013898019999999999 0 0.001391622 0 0.001391722 3.3 0.001391862 3.3 0.001391962 0 0.001393542 0 0.001393642 3.3 0.0013937819999999999 3.3 0.001393882 0 0.001394022 0 0.001394122 3.3 0.0013942619999999998 3.3 0.001394362 0 0.001394502 0 0.001394602 3.3 0.0013947419999999998 3.3 0.0013948419999999999 0 0.001394862 0 0.001394962 3.3 0.001395222 3.3 0.001395322 0 0.0013954619999999999 0 0.001395562 3.3 0.001395702 3.3 0.001395802 0 0.001395822 0 0.001395922 3.3 0.0013959419999999998 3.3 0.001396042 0 0.001396062 0 0.001396162 3.3 0.001396182 3.3 0.001396282 0 0.0013964219999999998 0 0.0013965219999999999 3.3 0.001396662 3.3 0.001396762 0 0.0013976219999999998 0 0.001397722 3.3 0.001397782 3.3 0.001397882 0 0.001399542 0 0.001399642 3.3 0.001399782 3.3 0.001399882 0 0.001401462 0 0.001401562 3.3 0.001402062 3.3 0.001402162 0 0.001402422 0 0.001402522 3.3 0.0014026619999999998 3.3 0.0014027619999999999 0 0.0014030219999999999 0 0.001403122 3.3 0.001403382 3.3 0.001403482 0 0.0014043419999999998 0 0.0014044419999999999 3.3 0.001405422 3.3 0.001405522 0 0.0014055419999999999 0 0.001405642 3.3 0.001405702 3.3 0.001405802 0 0.001407462 0 0.001407562 3.3 0.0014077019999999998 3.3 0.0014078019999999999 0 0.0014093819999999998 0 0.0014094819999999999 3.3 0.001409622 3.3 0.001409722 0 0.001410342 0 0.001410442 3.3 0.001410702 3.3 0.001410802 0 0.001410822 0 0.001410922 3.3 0.0014109419999999999 3.3 0.001411042 0 0.001411302 0 0.001411402 3.3 0.001411542 3.3 0.001411642 0 0.001412382 0 0.001412482 3.3 0.001412502 3.3 0.001412602 0 0.001413342 0 0.001413442 3.3 0.0014134619999999999 3.3 0.001413562 0 0.001415382 0 0.001415482 3.3 0.0014156219999999998 3.3 0.001415722 0 0.0014173019999999998 0 0.001417402 3.3 0.001417542 3.3 0.001417642 0 0.0014177819999999998 0 0.0014178819999999999 3.3 0.001418022 3.3 0.001418122 0 0.001418262 0 0.001418362 3.3 0.0014185019999999999 3.3 0.001418602 0 0.0014186219999999998 0 0.0014187219999999999 3.3 0.0014189819999999998 3.3 0.001419082 0 0.001419222 0 0.001419322 3.3 0.0014194619999999998 3.3 0.0014195619999999999 0 0.001419582 0 0.001419682 3.3 0.001419702 3.3 0.001419802 0 0.0014198219999999998 0 0.001419922 3.3 0.001419942 3.3 0.001420042 0 0.0014201819999999999 0 0.001420282 3.3 0.001420422 3.3 0.001420522 0 0.001421382 0 0.001421482 3.3 0.0014215419999999998 3.3 0.0014216419999999999 0 0.001423302 0 0.001423402 3.3 0.0014235419999999999 3.3 0.001423642 0 0.0014252219999999999 0 0.001425322 3.3 0.001425822 3.3 0.001425922 0 0.001426182 0 0.001426282 3.3 0.0014264219999999999 3.3 0.001426522 0 0.001426782 0 0.001426882 3.3 0.001427142 3.3 0.001427242 0 0.0014281019999999999 0 0.001428202 3.3 0.001429182 3.3 0.001429282 0 0.001429302 0 0.001429402 3.3 0.0014294619999999998 3.3 0.0014295619999999999 0 0.001431222 0 0.001431322 3.3 0.0014314619999999999 3.3 0.001431562 0 0.0014331419999999999 0 0.001433242 3.3 0.001433382 3.3 0.001433482 0 0.0014341019999999998 0 0.0014342019999999999 3.3 0.0014344619999999998 3.3 0.001434562 0 0.001434582 0 0.001434682 3.3 0.001434702 3.3 0.001434802 0 0.001435062 0 0.001435162 3.3 0.0014353019999999998 3.3 0.001435402 0 0.0014361419999999998 0 0.001436242 3.3 0.001436262 3.3 0.001436362 0 0.001437102 0 0.001437202 3.3 0.001437222 3.3 0.001437322 0 0.0014391419999999998 0 0.0014392419999999999 3.3 0.001439382 3.3 0.001439482 0 0.001441062 0 0.001441162 3.3 0.001441302 3.3 0.001441402 0 0.0014415419999999999 0 0.001441642 3.3 0.001441782 3.3 0.001441882 0 0.0014420219999999998 0 0.001442122 3.3 0.001442262 3.3 0.001442362 0 0.0014423819999999999 0 0.001442482 3.3 0.001442742 3.3 0.001442842 0 0.001442982 0 0.001443082 3.3 0.0014432219999999999 3.3 0.001443322 0 0.001443342 0 0.001443442 3.3 0.001443462 3.3 0.001443562 0 0.001443582 0 0.001443682 3.3 0.0014437019999999998 3.3 0.0014438019999999999 0 0.001443942 0 0.001444042 3.3 0.001444182 3.3 0.001444282 0 0.001445142 0 0.001445242 3.3 0.0014453019999999999 3.3 0.001445402 0 0.0014470619999999998 0 0.0014471619999999999 3.3 0.001447302 3.3 0.001447402 0 0.001448982 0 0.001449082 3.3 0.0014495819999999998 3.3 0.0014496819999999999 0 0.0014499419999999999 0 0.001450042 3.3 0.001450182 3.3 0.001450282 0 0.001450542 0 0.001450642 3.3 0.001450902 3.3 0.001451002 0 0.001451862 0 0.001451962 3.3 0.0014529419999999998 3.3 0.0014530419999999999 0 0.001453062 0 0.001453162 3.3 0.0014532219999999999 3.3 0.001453322 0 0.0014549819999999998 0 0.001455082 3.3 0.001455222 3.3 0.001455322 0 0.001456902 0 0.001457002 3.3 0.0014571419999999998 3.3 0.0014572419999999999 0 0.0014578619999999999 0 0.001457962 3.3 0.001458222 3.3 0.001458322 0 0.0014583419999999998 0 0.001458442 3.3 0.001458462 3.3 0.001458562 0 0.0014588219999999998 0 0.0014589219999999999 3.3 0.001459062 3.3 0.001459162 0 0.001459902 0 0.001460002 3.3 0.0014600219999999998 3.3 0.001460122 0 0.0014608619999999998 0 0.001460962 3.3 0.001460982 3.3 0.001461082 0 0.0014629019999999999 0 0.001463002 3.3 0.001463142 3.3 0.001463242 0 0.001464822 0 0.001464922 3.3 0.0014650619999999998 3.3 0.0014651619999999999 0 0.001465302 0 0.001465402 3.3 0.001465542 3.3 0.001465642 0 0.001465782 0 0.001465882 3.3 0.001466022 3.3 0.001466122 0 0.001466142 0 0.001466242 3.3 0.001466502 3.3 0.001466602 0 0.0014667419999999998 0 0.0014668419999999999 3.3 0.001466982 3.3 0.001467082 0 0.0014671019999999999 0 0.001467202 3.3 0.001467222 3.3 0.001467322 0 0.001467342 0 0.001467442 3.3 0.0014674619999999999 3.3 0.001467562 0 0.001467702 0 0.001467802 3.3 0.0014679419999999999 3.3 0.001468042 0 0.001468902 0 0.001469002 3.3 0.001469062 3.3 0.001469162 0 0.0014708219999999999 0 0.001470922 3.3 0.001471062 3.3 0.001471162 0 0.001472742 0 0.001472842 3.3 0.0014733419999999999 3.3 0.001473442 0 0.001473702 0 0.001473802 3.3 0.001473942 3.3 0.001474042 0 0.0014743019999999998 0 0.0014744019999999999 3.3 0.0014746619999999998 3.3 0.001474762 0 0.001475622 0 0.001475722 3.3 0.0014767019999999999 3.3 0.001476802 0 0.0014768219999999998 0 0.0014769219999999999 3.3 0.001476982 3.3 0.001477082 0 0.001478742 0 0.001478842 3.3 0.001478982 3.3 0.001479082 0 0.001480662 0 0.001480762 3.3 0.0014809019999999999 3.3 0.001481002 0 0.001481622 0 0.001481722 3.3 0.001481982 3.3 0.001482082 0 0.001482102 0 0.001482202 3.3 0.0014822219999999998 3.3 0.001482322 0 0.0014825819999999999 0 0.001482682 3.3 0.001482822 3.3 0.001482922 0 0.001483662 0 0.001483762 3.3 0.001483782 3.3 0.001483882 0 0.001484622 0 0.001484722 3.3 0.0014847419999999998 3.3 0.0014848419999999999 0 0.001486662 0 0.001486762 3.3 0.001486902 3.3 0.001487002 0 0.001488582 0 0.001488682 3.3 0.0014888219999999999 3.3 0.001488922 0 0.001489062 0 0.001489162 3.3 0.0014893019999999999 3.3 0.001489402 0 0.001489542 0 0.001489642 3.3 0.0014897819999999998 3.3 0.0014898819999999999 0 0.001489902 0 0.001490002 3.3 0.001490262 3.3 0.001490362 0 0.0014905019999999999 0 0.001490602 3.3 0.001490742 3.3 0.001490842 0 0.001490862 0 0.001490962 3.3 0.0014909819999999999 3.3 0.001491082 0 0.001491102 0 0.001491202 3.3 0.001491222 3.3 0.001491322 0 0.0014914619999999998 0 0.0014915619999999999 3.3 0.001491702 3.3 0.001491802 0 0.0014926619999999999 0 0.001492762 3.3 0.001492822 3.3 0.001492922 0 0.001494582 0 0.001494682 3.3 0.0014948219999999998 3.3 0.0014949219999999999 0 0.0014965019999999998 0 0.0014966019999999999 3.3 0.001497102 3.3 0.001497202 0 0.001497462 0 0.001497562 3.3 0.0014977019999999998 3.3 0.001497802 0 0.0014980619999999999 0 0.001498162 3.3 0.001498422 3.3 0.001498522 0 0.0014993819999999998 0 0.001499482 3.3 0.001500462 3.3 0.001500562 0 0.0015005819999999999 0 0.001500682 3.3 0.001500742 3.3 0.001500842 0 0.001502502 0 0.001502602 3.3 0.0015027419999999998 3.3 0.001502842 0 0.0015044219999999998 0 0.0015045219999999999 3.3 0.001504662 3.3 0.001504762 0 0.001505382 0 0.001505482 3.3 0.001505742 3.3 0.001505842 0 0.001505862 0 0.001505962 3.3 0.001505982 3.3 0.001506082 0 0.001506342 0 0.001506442 3.3 0.001506582 3.3 0.001506682 0 0.001507422 0 0.001507522 3.3 0.001507542 3.3 0.001507642 0 0.001508382 0 0.001508482 3.3 0.0015085019999999999 3.3 0.001508602 0 0.001510422 0 0.001510522 3.3 0.0015106619999999999 3.3 0.001510762 0 0.0015123419999999999 0 0.001512442 3.3 0.001512582 3.3 0.001512682 0 0.0015128219999999998 0 0.0015129219999999999 3.3 0.001513062 3.3 0.001513162 0 0.001513302 0 0.001513402 3.3 0.0015135419999999999 3.3 0.001513642 0 0.0015136619999999998 0 0.0015137619999999999 3.3 0.0015140219999999999 3.3 0.001514122 0 0.001514262 0 0.001514362 3.3 0.0015145019999999998 3.3 0.0015146019999999999 0 0.001514622 0 0.001514722 3.3 0.001514742 3.3 0.001514842 0 0.0015148619999999998 0 0.001514962 3.3 0.001514982 3.3 0.001515082 0 0.0015152219999999999 0 0.001515322 3.3 0.001515462 3.3 0.001515562 0 0.001516422 0 0.001516522 3.3 0.0015165819999999998 3.3 0.0015166819999999999 0 0.001518342 0 0.001518442 3.3 0.0015185819999999999 3.3 0.001518682 0 0.0015202619999999999 0 0.001520362 3.3 0.001520862 3.3 0.001520962 0 0.0015212219999999998 0 0.0015213219999999999 3.3 0.001521462 3.3 0.001521562 0 0.001521822 0 0.001521922 3.3 0.001522182 3.3 0.001522282 0 0.001523142 0 0.001523242 3.3 0.001524222 3.3 0.001524322 0 0.001524342 0 0.001524442 3.3 0.0015245019999999998 3.3 0.001524602 0 0.001526262 0 0.001526362 3.3 0.001526502 3.3 0.001526602 0 0.0015281819999999999 0 0.001528282 3.3 0.001528422 3.3 0.001528522 0 0.0015291419999999998 0 0.0015292419999999999 3.3 0.0015295019999999999 3.3 0.001529602 0 0.001529622 0 0.001529722 3.3 0.001529742 3.3 0.001529842 0 0.001530102 0 0.001530202 3.3 0.0015303419999999999 3.3 0.001530442 0 0.0015311819999999999 0 0.001531282 3.3 0.001531302 3.3 0.001531402 0 0.001532142 0 0.001532242 3.3 0.001532262 3.3 0.001532362 0 0.0015341819999999998 0 0.0015342819999999999 3.3 0.001534422 3.3 0.001534522 0 0.001536102 0 0.001536202 3.3 0.001536342 3.3 0.001536442 0 0.0015365819999999999 0 0.001536682 3.3 0.001536822 3.3 0.001536922 0 0.0015370619999999998 0 0.001537162 3.3 0.001537302 3.3 0.001537402 0 0.0015374219999999999 0 0.001537522 3.3 0.001537782 3.3 0.001537882 0 0.001538022 0 0.001538122 3.3 0.0015382619999999999 3.3 0.001538362 0 0.0015383819999999998 0 0.0015384819999999999 3.3 0.001538502 3.3 0.001538602 0 0.001538622 0 0.001538722 3.3 0.0015387419999999998 3.3 0.001538842 0 0.001538982 0 0.001539082 3.3 0.0015392219999999998 3.3 0.0015393219999999999 0 0.001540182 0 0.001540282 3.3 0.0015403419999999999 3.3 0.001540442 0 0.0015421019999999998 0 0.001542202 3.3 0.001542342 3.3 0.001542442 0 0.001544022 0 0.001544122 3.3 0.0015446219999999998 3.3 0.001544722 0 0.0015449819999999999 0 0.001545082 3.3 0.001545222 3.3 0.001545322 0 0.001545582 0 0.001545682 3.3 0.001545942 3.3 0.001546042 0 0.001546902 0 0.001547002 3.3 0.0015479819999999998 3.3 0.0015480819999999999 0 0.001548102 0 0.001548202 3.3 0.001548262 3.3 0.001548362 0 0.0015500219999999999 0 0.001550122 3.3 0.001550262 3.3 0.001550362 0 0.001551942 0 0.001552042 3.3 0.0015521819999999998 3.3 0.0015522819999999999 0 0.0015529019999999999 0 0.001553002 3.3 0.001553262 3.3 0.001553362 0 0.0015533819999999999 0 0.001553482 3.3 0.001553502 3.3 0.001553602 0 0.0015538619999999998 0 0.0015539619999999999 3.3 0.001554102 3.3 0.001554202 0 0.001554942 0 0.001555042 3.3 0.0015550619999999999 3.3 0.001555162 0 0.0015559019999999998 0 0.001556002 3.3 0.001556022 3.3 0.001556122 0 0.0015579419999999999 0 0.001558042 3.3 0.001558182 3.3 0.001558282 0 0.001559862 0 0.001559962 3.3 0.0015601019999999998 3.3 0.001560202 0 0.001560342 0 0.001560442 3.3 0.0015605819999999998 3.3 0.0015606819999999999 0 0.001560822 0 0.001560922 3.3 0.001561062 3.3 0.001561162 0 0.001561182 0 0.001561282 3.3 0.001561542 3.3 0.001561642 0 0.0015617819999999998 0 0.001561882 3.3 0.001562022 3.3 0.001562122 0 0.0015621419999999999 0 0.001562242 3.3 0.0015622619999999998 3.3 0.0015623619999999999 0 0.001562382 0 0.001562482 3.3 0.001562502 3.3 0.001562602 0 0.001562742 0 0.001562842 3.3 0.0015629819999999999 3.3 0.001563082 0 0.0015639419999999998 0 0.0015640419999999999 3.3 0.001564102 3.3 0.001564202 0 0.001565862 0 0.001565962 3.3 0.001566102 3.3 0.001566202 0 0.001567782 0 0.001567882 3.3 0.001568382 3.3 0.001568482 0 0.001568742 0 0.001568842 3.3 0.001568982 3.3 0.001569082 0 0.0015693419999999998 0 0.0015694419999999999 3.3 0.0015697019999999999 3.3 0.001569802 0 0.001570662 0 0.001570762 3.3 0.0015717419999999999 3.3 0.001571842 0 0.0015718619999999998 0 0.0015719619999999999 3.3 0.001572022 3.3 0.001572122 0 0.001573782 0 0.001573882 3.3 0.001574022 3.3 0.001574122 0 0.001575702 0 0.001575802 3.3 0.0015759419999999999 3.3 0.001576042 0 0.001576662 0 0.001576762 3.3 0.001577022 3.3 0.001577122 0 0.001577142 0 0.001577242 3.3 0.0015772619999999998 3.3 0.001577362 0 0.0015776219999999999 0 0.001577722 3.3 0.001577862 3.3 0.001577962 0 0.001578702 0 0.001578802 3.3 0.001578822 3.3 0.001578922 0 0.001579662 0 0.001579762 3.3 0.0015797819999999998 3.3 0.001579882 0 0.001581702 0 0.001581802 3.3 0.0015819419999999998 3.3 0.0015820419999999999 0 0.0015836219999999998 0 0.0015837219999999999 3.3 0.001583862 3.3 0.001583962 0 0.001584102 0 0.001584202 3.3 0.0015843419999999999 3.3 0.001584442 0 0.001584582 0 0.001584682 3.3 0.0015848219999999998 3.3 0.001584922 0 0.001584942 0 0.001585042 3.3 0.0015853019999999998 3.3 0.0015854019999999999 0 0.001585542 0 0.001585642 3.3 0.001585782 3.3 0.001585882 0 0.001585902 0 0.001586002 3.3 0.0015860219999999999 3.3 0.001586122 0 0.0015861419999999998 0 0.0015862419999999999 3.3 0.001586262 3.3 0.001586362 0 0.0015865019999999998 0 0.0015866019999999999 3.3 0.001586742 3.3 0.001586842 0 0.0015877019999999999 0 0.001587802 3.3 0.001587862 3.3 0.001587962 0 0.001589622 0 0.001589722 3.3 0.0015898619999999998 3.3 0.0015899619999999999 0 0.0015915419999999998 0 0.0015916419999999999 3.3 0.001592142 3.3 0.001592242 0 0.001592502 0 0.001592602 3.3 0.0015927419999999999 3.3 0.001592842 0 0.0015931019999999999 0 0.001593202 3.3 0.001593462 3.3 0.001593562 0 0.0015944219999999999 0 0.001594522 3.3 0.001595502 3.3 0.001595602 0 0.0015956219999999999 0 0.001595722 3.3 0.001595782 3.3 0.001595882 0 0.001597542 0 0.001597642 3.3 0.0015977819999999998 3.3 0.001597882 0 0.0015994619999999998 0 0.001599562 3.3 0.001599702 3.3 0.001599802 0 0.001600422 0 0.001600522 3.3 0.0016007819999999998 3.3 0.0016008819999999999 0 0.001600902 0 0.001601002 3.3 0.001601022 3.3 0.001601122 0 0.001601382 0 0.001601482 3.3 0.0016016219999999998 3.3 0.0016017219999999999 0 0.0016024619999999998 0 0.0016025619999999999 3.3 0.001602582 3.3 0.001602682 0 0.001603422 0 0.001603522 3.3 0.001603542 3.3 0.001603642 0 0.001605462 0 0.001605562 3.3 0.0016057019999999999 3.3 0.001605802 0 0.0016073819999999999 0 0.001607482 3.3 0.001607622 3.3 0.001607722 0 0.0016078619999999998 0 0.0016079619999999999 3.3 0.001608102 3.3 0.001608202 0 0.001608342 0 0.001608442 3.3 0.001608582 3.3 0.001608682 0 0.0016087019999999998 0 0.0016088019999999999 3.3 0.0016090619999999999 3.3 0.001609162 0 0.001609302 0 0.001609402 3.3 0.0016095419999999998 3.3 0.0016096419999999999 0 0.001609662 0 0.001609762 3.3 0.001609782 3.3 0.001609882 0 0.0016099019999999999 0 0.001610002 3.3 0.001610022 3.3 0.001610122 0 0.0016102619999999999 0 0.001610362 3.3 0.001610502 3.3 0.001610602 0 0.001611462 0 0.001611562 3.3 0.0016116219999999998 3.3 0.001611722 0 0.001613382 0 0.001613482 3.3 0.0016136219999999999 3.3 0.001613722 0 0.0016153019999999999 0 0.001615402 3.3 0.001615902 3.3 0.001616002 0 0.0016162619999999998 0 0.0016163619999999999 3.3 0.001616502 3.3 0.001616602 0 0.001616862 0 0.001616962 3.3 0.001617222 3.3 0.001617322 0 0.001618182 0 0.001618282 3.3 0.001619262 3.3 0.001619362 0 0.001619382 0 0.001619482 3.3 0.0016195419999999999 3.3 0.001619642 0 0.0016213019999999998 0 0.0016214019999999999 3.3 0.001621542 3.3 0.001621642 0 0.001623222 0 0.001623322 3.3 0.001623462 3.3 0.001623562 0 0.0016241819999999998 0 0.001624282 3.3 0.0016245419999999999 3.3 0.001624642 0 0.0016246619999999998 0 0.0016247619999999999 3.3 0.001624782 3.3 0.001624882 0 0.001625142 0 0.001625242 3.3 0.0016253819999999999 3.3 0.001625482 0 0.0016262219999999999 0 0.001626322 3.3 0.0016263419999999998 3.3 0.0016264419999999999 0 0.0016271819999999998 0 0.0016272819999999999 3.3 0.001627302 3.3 0.001627402 0 0.0016292219999999998 0 0.0016293219999999999 3.3 0.001629462 3.3 0.001629562 0 0.001631142 0 0.001631242 3.3 0.001631382 3.3 0.001631482 0 0.0016316219999999999 0 0.001631722 3.3 0.001631862 3.3 0.001631962 0 0.0016321019999999999 0 0.001632202 3.3 0.001632342 3.3 0.001632442 0 0.0016324619999999999 0 0.001632562 3.3 0.001632822 3.3 0.001632922 0 0.001633062 0 0.001633162 3.3 0.0016333019999999999 3.3 0.001633402 0 0.0016334219999999998 0 0.0016335219999999999 3.3 0.001633542 3.3 0.001633642 0 0.001633662 0 0.001633762 3.3 0.0016337819999999999 3.3 0.001633882 0 0.001634022 0 0.001634122 3.3 0.0016342619999999998 3.3 0.0016343619999999999 0 0.001635222 0 0.001635322 3.3 0.001635382 3.3 0.001635482 0 0.0016371419999999999 0 0.001637242 3.3 0.001637382 3.3 0.001637482 0 0.001639062 0 0.001639162 3.3 0.0016396619999999998 3.3 0.001639762 0 0.0016400219999999999 0 0.001640122 3.3 0.001640262 3.3 0.001640362 0 0.001640622 0 0.001640722 3.3 0.0016409819999999998 3.3 0.0016410819999999999 0 0.001641942 0 0.001642042 3.3 0.0016430219999999998 3.3 0.001643122 0 0.001643142 0 0.001643242 3.3 0.001643302 3.3 0.001643402 0 0.0016450619999999999 0 0.001645162 3.3 0.001645302 3.3 0.001645402 0 0.001646982 0 0.001647082 3.3 0.0016472219999999998 3.3 0.001647322 0 0.001647942 0 0.001648042 3.3 0.001648302 3.3 0.001648402 0 0.0016484219999999999 0 0.001648522 3.3 0.0016485419999999998 3.3 0.0016486419999999999 0 0.0016489019999999998 0 0.0016490019999999999 3.3 0.001649142 3.3 0.001649242 0 0.001649982 0 0.001650082 3.3 0.0016501019999999999 3.3 0.001650202 0 0.0016509419999999999 0 0.001651042 3.3 0.001651062 3.3 0.001651162 0 0.0016529819999999999 0 0.001653082 3.3 0.001653222 3.3 0.001653322 0 0.001654902 0 0.001655002 3.3 0.0016551419999999999 3.3 0.001655242 0 0.001655382 0 0.001655482 3.3 0.0016556219999999998 3.3 0.0016557219999999999 0 0.001655862 0 0.001655962 3.3 0.001656102 3.3 0.001656202 0 0.001656222 0 0.001656322 3.3 0.001656582 3.3 0.001656682 0 0.0016568219999999999 0 0.001656922 3.3 0.001657062 3.3 0.001657162 0 0.0016571819999999999 0 0.001657282 3.3 0.0016573019999999998 3.3 0.0016574019999999999 0 0.001657422 0 0.001657522 3.3 0.001657542 3.3 0.001657642 0 0.001657782 0 0.001657882 3.3 0.0016580219999999999 3.3 0.001658122 0 0.0016589819999999998 0 0.0016590819999999999 3.3 0.001659142 3.3 0.001659242 0 0.001660902 0 0.001661002 3.3 0.001661142 3.3 0.001661242 0 0.001662822 0 0.001662922 3.3 0.001663422 3.3 0.001663522 0 0.001663782 0 0.001663882 3.3 0.0016640219999999998 3.3 0.0016641219999999999 0 0.0016643819999999998 0 0.001664482 3.3 0.0016647419999999999 3.3 0.001664842 0 0.0016657019999999998 0 0.0016658019999999999 3.3 0.001666782 3.3 0.001666882 0 0.0016669019999999998 0 0.001667002 3.3 0.001667062 3.3 0.001667162 0 0.001668822 0 0.001668922 3.3 0.0016690619999999998 3.3 0.0016691619999999999 0 0.001670742 0 0.001670842 3.3 0.001670982 3.3 0.001671082 0 0.001671702 0 0.001671802 3.3 0.001672062 3.3 0.001672162 0 0.001672182 0 0.001672282 3.3 0.0016723019999999999 3.3 0.001672402 0 0.0016726619999999999 0 0.001672762 3.3 0.001672902 3.3 0.001673002 0 0.001673742 0 0.001673842 3.3 0.001673862 3.3 0.001673962 0 0.001674702 0 0.001674802 3.3 0.0016748219999999999 3.3 0.001674922 0 0.001676742 0 0.001676842 3.3 0.0016769819999999998 3.3 0.0016770819999999999 0 0.0016786619999999998 0 0.0016787619999999999 3.3 0.001678902 3.3 0.001679002 0 0.001679142 0 0.001679242 3.3 0.0016793819999999999 3.3 0.001679482 0 0.001679622 0 0.001679722 3.3 0.0016798619999999998 3.3 0.001679962 0 0.001679982 0 0.001680082 3.3 0.0016803419999999998 3.3 0.0016804419999999999 0 0.001680582 0 0.001680682 3.3 0.001680822 3.3 0.001680922 0 0.001680942 0 0.001681042 3.3 0.0016810619999999999 3.3 0.001681162 0 0.0016811819999999998 0 0.0016812819999999999 3.3 0.001681302 3.3 0.001681402 0 0.0016815419999999998 0 0.001681642 3.3 0.001681782 3.3 0.001681882 0 0.0016827419999999999 0 0.001682842 3.3 0.001682902 3.3 0.001683002 0 0.001684662 0 0.001684762 3.3 0.0016849019999999998 3.3 0.001685002 0 0.0016865819999999998 0 0.001686682 3.3 0.001687182 3.3 0.001687282 0 0.001687542 0 0.001687642 3.3 0.0016877819999999999 3.3 0.001687882 0 0.001688142 0 0.001688242 3.3 0.001688502 3.3 0.001688602 0 0.0016894619999999999 0 0.001689562 3.3 0.001690542 3.3 0.001690642 0 0.001690662 0 0.001690762 3.3 0.0016908219999999998 3.3 0.0016909219999999999 0 0.001692582 0 0.001692682 3.3 0.0016928219999999999 3.3 0.001692922 0 0.0016945019999999999 0 0.001694602 3.3 0.001694742 3.3 0.001694842 0 0.001695462 0 0.001695562 3.3 0.0016958219999999998 3.3 0.0016959219999999999 0 0.001695942 0 0.001696042 3.3 0.001696062 3.3 0.001696162 0 0.001696422 0 0.001696522 3.3 0.0016966619999999998 3.3 0.0016967619999999999 0 0.0016975019999999998 0 0.0016976019999999999 3.3 0.001697622 3.3 0.001697722 0 0.001698462 0 0.001698562 3.3 0.001698582 3.3 0.001698682 0 0.001700502 0 0.001700602 3.3 0.0017007419999999999 3.3 0.001700842 0 0.0017024219999999999 0 0.001702522 3.3 0.001702662 3.3 0.001702762 0 0.0017029019999999998 0 0.001703002 3.3 0.001703142 3.3 0.001703242 0 0.0017033819999999998 0 0.0017034819999999999 3.3 0.001703622 3.3 0.001703722 0 0.0017037419999999998 0 0.001703842 3.3 0.0017041019999999999 3.3 0.001704202 0 0.001704342 0 0.001704442 3.3 0.0017045819999999998 3.3 0.001704682 0 0.001704702 0 0.001704802 3.3 0.001704822 3.3 0.001704922 0 0.0017049419999999999 0 0.001705042 3.3 0.0017050619999999998 3.3 0.0017051619999999999 0 0.001705302 0 0.001705402 3.3 0.001705542 3.3 0.001705642 0 0.001706502 0 0.001706602 3.3 0.0017066619999999998 3.3 0.001706762 0 0.0017084219999999998 0 0.0017085219999999999 3.3 0.001708662 3.3 0.001708762 0 0.001710342 0 0.001710442 3.3 0.0017109419999999998 3.3 0.0017110419999999999 0 0.0017113019999999998 0 0.0017114019999999999 3.3 0.001711542 3.3 0.001711642 0 0.001711902 0 0.001712002 3.3 0.001712262 3.3 0.001712362 0 0.001713222 0 0.001713322 3.3 0.001714302 3.3 0.001714402 0 0.001714422 0 0.001714522 3.3 0.0017145819999999999 3.3 0.001714682 0 0.0017163419999999998 0 0.0017164419999999999 3.3 0.001716582 3.3 0.001716682 0 0.001718262 0 0.001718362 3.3 0.001718502 3.3 0.001718602 0 0.0017192219999999999 0 0.001719322 3.3 0.0017195819999999999 3.3 0.001719682 0 0.0017197019999999998 0 0.0017198019999999999 3.3 0.001719822 3.3 0.001719922 0 0.001720182 0 0.001720282 3.3 0.0017204219999999999 3.3 0.001720522 0 0.0017212619999999999 0 0.001721362 3.3 0.0017213819999999998 3.3 0.0017214819999999999 0 0.0017222219999999998 0 0.0017223219999999999 3.3 0.001722342 3.3 0.001722442 0 0.0017242619999999998 0 0.001724362 3.3 0.001724502 3.3 0.001724602 0 0.001726182 0 0.001726282 3.3 0.0017264219999999998 3.3 0.0017265219999999999 0 0.001726662 0 0.001726762 3.3 0.001726902 3.3 0.001727002 0 0.0017271419999999999 0 0.001727242 3.3 0.001727382 3.3 0.001727482 0 0.001727502 0 0.001727602 3.3 0.001727862 3.3 0.001727962 0 0.0017281019999999998 0 0.0017282019999999999 3.3 0.001728342 3.3 0.001728442 0 0.0017284619999999998 0 0.001728562 3.3 0.001728582 3.3 0.001728682 0 0.001728702 0 0.001728802 3.3 0.0017288219999999999 3.3 0.001728922 0 0.001729062 0 0.001729162 3.3 0.0017293019999999998 3.3 0.001729402 0 0.001730262 0 0.001730362 3.3 0.001730422 3.3 0.001730522 0 0.0017321819999999999 0 0.001732282 3.3 0.001732422 3.3 0.001732522 0 0.001734102 0 0.001734202 3.3 0.0017347019999999999 3.3 0.001734802 0 0.0017350619999999999 0 0.001735162 3.3 0.001735302 3.3 0.001735402 0 0.001735662 0 0.001735762 3.3 0.0017360219999999998 3.3 0.0017361219999999999 0 0.001736982 0 0.001737082 3.3 0.0017380619999999999 3.3 0.001738162 0 0.001738182 0 0.001738282 3.3 0.001738342 3.3 0.001738442 0 0.0017401019999999999 0 0.001740202 3.3 0.001740342 3.3 0.001740442 0 0.001742022 0 0.001742122 3.3 0.0017422619999999998 3.3 0.001742362 0 0.001742982 0 0.001743082 3.3 0.001743342 3.3 0.001743442 0 0.0017434619999999999 0 0.001743562 3.3 0.0017435819999999998 3.3 0.0017436819999999999 0 0.0017439419999999998 0 0.001744042 3.3 0.001744182 3.3 0.001744282 0 0.001745022 0 0.001745122 3.3 0.0017451419999999999 3.3 0.001745242 0 0.0017459819999999999 0 0.001746082 3.3 0.0017461019999999998 3.3 0.0017462019999999999 0 0.001748022 0 0.001748122 3.3 0.001748262 3.3 0.001748362 0 0.001749942 0 0.001750042 3.3 0.0017501819999999999 3.3 0.001750282 0 0.001750422 0 0.001750522 3.3 0.0017506619999999998 3.3 0.0017507619999999999 0 0.001750902 0 0.001751002 3.3 0.0017511419999999998 3.3 0.0017512419999999999 0 0.001751262 0 0.001751362 3.3 0.001751622 3.3 0.001751722 0 0.0017518619999999999 0 0.001751962 3.3 0.001752102 3.3 0.001752202 0 0.001752222 0 0.001752322 3.3 0.0017523419999999998 3.3 0.0017524419999999999 0 0.001752462 0 0.001752562 3.3 0.001752582 3.3 0.001752682 0 0.0017528219999999998 0 0.0017529219999999999 3.3 0.001753062 3.3 0.001753162 0 0.0017540219999999998 0 0.0017541219999999999 3.3 0.001754182 3.3 0.001754282 0 0.001755942 0 0.001756042 3.3 0.001756182 3.3 0.001756282 0 0.001757862 0 0.001757962 3.3 0.001758462 3.3 0.001758562 0 0.001758822 0 0.001758922 3.3 0.0017590619999999998 3.3 0.0017591619999999999 0 0.0017594219999999999 0 0.001759522 3.3 0.0017597819999999999 3.3 0.001759882 0 0.0017607419999999998 0 0.0017608419999999999 3.3 0.001761822 3.3 0.001761922 0 0.0017619419999999998 0 0.001762042 3.3 0.001762102 3.3 0.001762202 0 0.001763862 0 0.001763962 3.3 0.0017641019999999998 3.3 0.0017642019999999999 0 0.0017657819999999998 0 0.0017658819999999999 3.3 0.001766022 3.3 0.001766122 0 0.001766742 0 0.001766842 3.3 0.001767102 3.3 0.001767202 0 0.001767222 0 0.001767322 3.3 0.0017673419999999999 3.3 0.001767442 0 0.001767702 0 0.001767802 3.3 0.001767942 3.3 0.001768042 0 0.001768782 0 0.001768882 3.3 0.001768902 3.3 0.001769002 0 0.001769742 0 0.001769842 3.3 0.0017698619999999999 3.3 0.001769962 0 0.001771782 0 0.001771882 3.3 0.0017720219999999998 3.3 0.0017721219999999999 0 0.0017737019999999998 0 0.0017738019999999999 3.3 0.001773942 3.3 0.001774042 0 0.001774182 0 0.001774282 3.3 0.001774422 3.3 0.001774522 0 0.001774662 0 0.001774762 3.3 0.0017749019999999999 3.3 0.001775002 0 0.001775022 0 0.001775122 3.3 0.0017753819999999998 3.3 0.0017754819999999999 0 0.001775622 0 0.001775722 3.3 0.001775862 3.3 0.001775962 0 0.001775982 0 0.001776082 3.3 0.0017761019999999999 3.3 0.001776202 0 0.0017762219999999998 0 0.0017763219999999999 3.3 0.001776342 3.3 0.001776442 0 0.0017765819999999999 0 0.001776682 3.3 0.001776822 3.3 0.001776922 0 0.0017777819999999999 0 0.001777882 3.3 0.0017779419999999998 3.3 0.0017780419999999999 0 0.001779702 0 0.001779802 3.3 0.0017799419999999999 3.3 0.001780042 0 0.0017816219999999998 0 0.001781722 3.3 0.001782222 3.3 0.001782322 0 0.001782582 0 0.001782682 3.3 0.0017828219999999999 3.3 0.001782922 0 0.001783182 0 0.001783282 3.3 0.001783542 3.3 0.001783642 0 0.0017845019999999999 0 0.001784602 3.3 0.001785582 3.3 0.001785682 0 0.001785702 0 0.001785802 3.3 0.0017858619999999998 3.3 0.0017859619999999999 0)

* spi_miso_ram - 6 transitions
V_spi_miso_ram spi_miso_ram 0 PWL(0 3.3 6.3581e-05 3.3 6.3681e-05 0 6.7461e-05 0 6.7561e-05 3.3 0.000122741 3.3 0.000122841 0 0.000126621 0 0.000126721 3.3 0.000134621 3.3 0.000134721 0 0.000138501 0 0.000138601 3.3)

* Include circuit netlist
.include "./femto.spice"
.end
