* NGSPICE file created from femto.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_4 abstract view
.subckt sky130_fd_sc_hd__dlxtn_4 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt femto LEDS RXD TXD VGND VPWR clk resetn spi_clk spi_clk_ram spi_cs_n spi_cs_n_ram
+ spi_miso spi_miso_ram spi_mosi spi_mosi_ram
X_09671_ _05856_ _06013_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__nand2_1
X_18869_ net643 _02389_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18573__30 VGND VGND VPWR VPWR _18573__30/HI net30 sky130_fd_sc_hd__conb_1
XFILLER_0_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09105_ _05456_ _05323_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__or2_2
X_15959__695 clknet_1_0__leaf__03691_ VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__inv_2
XFILLER_0_115_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09036_ CPU.aluIn1\[24\] _05387_ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13937__97 clknet_1_1__leaf__08478_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__inv_2
XFILLER_0_32_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13655__1033 clknet_1_0__leaf__08450_ VGND VGND VPWR VPWR net1089 sky130_fd_sc_hd__inv_2
XFILLER_0_142_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15658__456 clknet_1_0__leaf__03644_ VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__inv_2
Xhold340 CPU.rs2\[11\] VGND VGND VPWR VPWR net1637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold351 mapped_spi_flash.rcv_data\[5\] VGND VGND VPWR VPWR net1648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold362 per_uart.rx_avail VGND VGND VPWR VPWR net1659 sky130_fd_sc_hd__dlygate4sd3_1
X_13607__990 clknet_1_1__leaf__08445_ VGND VGND VPWR VPWR net1046 sky130_fd_sc_hd__inv_2
Xhold373 per_uart.uart0.rxd_reg\[3\] VGND VGND VPWR VPWR net1670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 CPU.registerFile\[6\]\[2\] VGND VGND VPWR VPWR net1681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 CPU.registerFile\[28\]\[30\] VGND VGND VPWR VPWR net1692 sky130_fd_sc_hd__dlygate4sd3_1
X_09938_ _05313_ _05769_ _05770_ net1396 VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__a22o_1
X_09869_ _06175_ _06203_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__nor2_2
Xhold1040 CPU.registerFile\[18\]\[13\] VGND VGND VPWR VPWR net2337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 CPU.registerFile\[23\]\[21\] VGND VGND VPWR VPWR net2348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 CPU.registerFile\[8\]\[28\] VGND VGND VPWR VPWR net2359 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ _07579_ VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__clkbuf_1
Xhold1073 CPU.registerFile\[7\]\[11\] VGND VGND VPWR VPWR net2370 sky130_fd_sc_hd__dlygate4sd3_1
X_12880_ _06486_ net2264 _08131_ VGND VGND VPWR VPWR _08140_ sky130_fd_sc_hd__mux2_1
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1084 CPU.registerFile\[31\]\[25\] VGND VGND VPWR VPWR net2381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1095 CPU.registerFile\[9\]\[19\] VGND VGND VPWR VPWR net2392 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ net2444 _07343_ _07537_ VGND VGND VPWR VPWR _07543_ sky130_fd_sc_hd__mux2_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03645_ clknet_0__03645_ VGND VGND VPWR VPWR clknet_1_0__leaf__03645_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _08780_ _08790_ _08594_ VGND VGND VPWR VPWR _08791_ sky130_fd_sc_hd__o21a_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _07506_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__clkbuf_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10713_ _06829_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__clkbuf_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14481_ CPU.registerFile\[30\]\[4\] CPU.registerFile\[31\]\[4\] _08645_ VGND VGND
+ VPWR VPWR _08723_ sky130_fd_sc_hd__mux2_1
X_11693_ _07469_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16220_ _03940_ _03941_ _03720_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13432_ _08396_ VGND VGND VPWR VPWR _08397_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_125_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10644_ _06791_ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16151_ _03741_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__buf_4
X_10575_ net1875 _06124_ _06750_ VGND VGND VPWR VPWR _06754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15102_ CPU.registerFile\[22\]\[19\] CPU.registerFile\[23\]\[19\] _02998_ VGND VGND
+ VPWR VPWR _03165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12314_ _07836_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__clkbuf_1
X_16082_ _03806_ _03807_ _03763_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15033_ _06418_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12245_ net1523 _07785_ _07794_ _07755_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12176_ _07739_ _07746_ VGND VGND VPWR VPWR _07747_ sky130_fd_sc_hd__or2_1
X_11127_ net1356 _07135_ VGND VGND VPWR VPWR _07144_ sky130_fd_sc_hd__or2_1
X_16984_ _04479_ _04683_ _04687_ _04446_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18723_ net512 _02247_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[23\] sky130_fd_sc_hd__dfxtp_1
X_11058_ _05284_ CPU.Bimm\[5\] VGND VGND VPWR VPWR _07094_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10009_ _06338_ VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__clkbuf_1
X_18654_ clknet_leaf_11_clk _02178_ VGND VGND VPWR VPWR CPU.rs2\[26\] sky130_fd_sc_hd__dfxtp_1
X_15866_ clknet_1_1__leaf__03654_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__buf_1
X_14817_ _08409_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__buf_4
X_17605_ net1463 _05159_ _05160_ _07108_ VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__o22a_1
XFILLER_0_149_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18585_ net406 net42 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_15797_ net1582 _08348_ net1590 VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__o21ai_1
X_17536_ _08335_ _06042_ _05073_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14748_ _02818_ _02819_ _08695_ VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17467_ _08311_ _06329_ _08331_ VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__or3_1
XFILLER_0_156_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14679_ _06061_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13715__1087 clknet_1_1__leaf__08456_ VGND VGND VPWR VPWR net1143 sky130_fd_sc_hd__inv_2
XFILLER_0_156_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16418_ _03963_ _04133_ _04135_ _04006_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__a211o_1
XFILLER_0_104_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17398_ clknet_1_1__leaf__08340_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__buf_1
XFILLER_0_27_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19137_ clknet_leaf_15_clk _02657_ VGND VGND VPWR VPWR CPU.PC\[19\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_132_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16349_ _06148_ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__clkbuf_4
X_19068_ net60 _02588_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__08494_ clknet_0__08494_ VGND VGND VPWR VPWR clknet_1_1__leaf__08494_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14258__386 clknet_1_1__leaf__08510_ VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__inv_2
XFILLER_0_11_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18019_ net1030 _01547_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__03639_ _03639_ VGND VGND VPWR VPWR clknet_0__03639_ sky130_fd_sc_hd__clkbuf_16
X_09723_ _06063_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__buf_4
X_09654_ CPU.PC\[20\] _05996_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09585_ _05927_ _05928_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__nor2_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_829 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13944__103 clknet_1_1__leaf__08479_ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__inv_2
XFILLER_0_64_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10360_ _06631_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__clkbuf_1
X_15892__635 clknet_1_1__leaf__03684_ VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__inv_2
XFILLER_0_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09019_ CPU.rs2\[23\] _05247_ _05251_ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__o21a_1
X_13732__1102 clknet_1_1__leaf__08458_ VGND VGND VPWR VPWR net1158 sky130_fd_sc_hd__inv_2
XFILLER_0_131_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10291_ net1728 _06413_ _06580_ VGND VGND VPWR VPWR _06586_ sky130_fd_sc_hd__mux2_1
X_12030_ CPU.registerFile\[24\]\[19\] _07337_ _07646_ VGND VGND VPWR VPWR _07649_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold170 mapped_spi_ram.cmd_addr\[8\] VGND VGND VPWR VPWR net1467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 per_uart.uart0.txd_reg\[6\] VGND VGND VPWR VPWR net1478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 mapped_spi_ram.rcv_data\[13\] VGND VGND VPWR VPWR net1489 sky130_fd_sc_hd__dlygate4sd3_1
X_13540__930 clknet_1_1__leaf__08438_ VGND VGND VPWR VPWR net986 sky130_fd_sc_hd__inv_2
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13990__145 clknet_1_0__leaf__08483_ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__inv_2
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ _06292_ net1940 _08167_ VGND VGND VPWR VPWR _08168_ sky130_fd_sc_hd__mux2_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _08108_ VGND VGND VPWR VPWR _08131_ sky130_fd_sc_hd__buf_4
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14602_ _06036_ VGND VGND VPWR VPWR _08841_ sky130_fd_sc_hd__clkbuf_4
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ net2019 _07326_ _07526_ VGND VGND VPWR VPWR _07534_ sky130_fd_sc_hd__mux2_1
X_18370_ net191 _01898_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ CPU.registerFile\[0\]\[31\] _08411_ _03632_ _06036_ VGND VGND VPWR VPWR _03633_
+ sky130_fd_sc_hd__o211a_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _08093_ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__clkbuf_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14533_ _08772_ _08773_ _08695_ VGND VGND VPWR VPWR _08774_ sky130_fd_sc_hd__mux2_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _07497_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17252_ CPU.registerFile\[15\]\[31\] CPU.registerFile\[14\]\[31\] _03698_ VGND VGND
+ VPWR VPWR _04948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14464_ _08585_ _08586_ CPU.registerFile\[1\]\[3\] VGND VGND VPWR VPWR _08707_ sky130_fd_sc_hd__a21o_1
X_11676_ _07460_ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16203_ CPU.registerFile\[16\]\[4\] _03848_ _03769_ _03925_ VGND VGND VPWR VPWR _03926_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13415_ _08386_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__clkbuf_1
X_17183_ _03766_ _04878_ _04880_ _03716_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__a211o_1
X_10627_ _06782_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14395_ CPU.registerFile\[16\]\[2\] _08412_ _08638_ _06037_ VGND VGND VPWR VPWR _08639_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16134_ CPU.registerFile\[8\]\[3\] _08394_ _06150_ _03857_ VGND VGND VPWR VPWR _03858_
+ sky130_fd_sc_hd__o211a_1
X_10558_ net2146 _05839_ _06739_ VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16065_ _03726_ _03727_ CPU.registerFile\[1\]\[1\] VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__a21o_1
X_13916__78 clknet_1_0__leaf__08476_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__inv_2
X_13277_ net1598 _08357_ VGND VGND VPWR VPWR _08358_ sky130_fd_sc_hd__or2_1
X_10489_ net1954 _05839_ _06702_ VGND VGND VPWR VPWR _06708_ sky130_fd_sc_hd__mux2_1
X_15016_ CPU.registerFile\[21\]\[17\] _02960_ VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__or2_1
X_12228_ _07783_ VGND VGND VPWR VPWR _07784_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12159_ net1466 _07714_ _07734_ _07713_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16967_ _04419_ _04668_ _04670_ _04383_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__a211o_1
X_18706_ net495 _02230_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[6\] sky130_fd_sc_hd__dfxtp_1
X_16898_ _04502_ _04591_ _04595_ _04603_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__a31o_2
X_18637_ clknet_leaf_17_clk _02161_ VGND VGND VPWR VPWR CPU.rs2\[9\] sky130_fd_sc_hd__dfxtp_1
X_13654__1032 clknet_1_0__leaf__08450_ VGND VGND VPWR VPWR net1088 sky130_fd_sc_hd__inv_2
X_15687__482 clknet_1_1__leaf__03647_ VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__inv_2
X_09370_ _05659_ _05678_ _05721_ _05683_ VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__a211o_1
X_18568_ net389 net25 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17519_ _05055_ _06111_ _05061_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__or3_1
X_18499_ net320 _02023_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_812 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13255__775 clknet_1_0__leaf__08344_ VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__inv_2
XFILLER_0_74_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15841__589 clknet_1_1__leaf__03679_ VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__inv_2
XFILLER_0_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14191__326 clknet_1_1__leaf__08503_ VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__08477_ clknet_0__08477_ VGND VGND VPWR VPWR clknet_1_1__leaf__08477_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17416__38 clknet_1_0__leaf__05014_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__inv_2
X_09706_ _05881_ _06039_ _06047_ _05744_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_69_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09637_ CPU.PC\[14\] _05980_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__nand2_1
X_14011__163 clknet_1_1__leaf__08486_ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__inv_2
X_14085__231 clknet_1_0__leaf__08492_ VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__inv_2
X_09568_ _05911_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_139_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13570__956 clknet_1_0__leaf__08442_ VGND VGND VPWR VPWR net1012 sky130_fd_sc_hd__inv_2
XFILLER_0_93_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09499_ _05831_ _05813_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11530_ _07382_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15900__642 clknet_1_0__leaf__03685_ VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__inv_2
X_11461_ _07336_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13200_ _05286_ _05290_ _06519_ _05296_ VGND VGND VPWR VPWR _08314_ sky130_fd_sc_hd__or4bb_1
X_10412_ _06599_ net2484 _06665_ VGND VGND VPWR VPWR _06667_ sky130_fd_sc_hd__mux2_1
X_11392_ _07293_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__05014_ clknet_0__05014_ VGND VGND VPWR VPWR clknet_1_0__leaf__05014_
+ sky130_fd_sc_hd__clkbuf_16
X_13131_ net1604 _08271_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__xor2_1
X_10343_ _06082_ VGND VGND VPWR VPWR _06620_ sky130_fd_sc_hd__buf_4
XFILLER_0_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13062_ net1418 VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__clkbuf_1
X_10274_ net1754 _06224_ _06569_ VGND VGND VPWR VPWR _06577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12013_ net2518 _07320_ _07635_ VGND VGND VPWR VPWR _07640_ sky130_fd_sc_hd__mux2_1
X_17870_ clknet_leaf_24_clk _00019_ VGND VGND VPWR VPWR CPU.cycles\[13\] sky130_fd_sc_hd__dfxtp_1
X_13714__1086 clknet_1_0__leaf__08456_ VGND VGND VPWR VPWR net1142 sky130_fd_sc_hd__inv_2
X_16821_ CPU.registerFile\[27\]\[19\] CPU.registerFile\[26\]\[19\] _04242_ VGND VGND
+ VPWR VPWR _04529_ sky130_fd_sc_hd__mux2_1
X_13321__821 clknet_1_1__leaf__08363_ VGND VGND VPWR VPWR net877 sky130_fd_sc_hd__inv_2
XFILLER_0_45_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16752_ CPU.registerFile\[9\]\[18\] _04460_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__or2_1
X_13964_ clknet_1_0__leaf__08473_ VGND VGND VPWR VPWR _08481_ sky130_fd_sc_hd__buf_1
X_12915_ _06106_ net1564 _08156_ VGND VGND VPWR VPWR _08159_ sky130_fd_sc_hd__mux2_1
X_16683_ _04305_ _04387_ _04393_ _04072_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_0__f__08497_ clknet_0__08497_ VGND VGND VPWR VPWR clknet_1_0__leaf__08497_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_158_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18422_ net243 _01950_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ _08122_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__clkbuf_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18353_ net174 _01881_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ CPU.registerFile\[24\]\[31\] _08582_ _03615_ _08540_ VGND VGND VPWR VPWR
+ _03616_ sky130_fd_sc_hd__o211a_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _08084_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__clkbuf_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14516_ CPU.registerFile\[22\]\[5\] CPU.registerFile\[23\]\[5\] _08756_ VGND VGND
+ VPWR VPWR _08757_ sky130_fd_sc_hd__mux2_1
X_11728_ _07487_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__clkbuf_1
X_18284_ net1295 _01812_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_15496_ CPU.registerFile\[13\]\[29\] CPU.registerFile\[12\]\[29\] _08794_ VGND VGND
+ VPWR VPWR _03549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17235_ _03722_ _04929_ _04931_ _04612_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__a211o_1
X_14447_ _08535_ _08684_ _08689_ _08554_ VGND VGND VPWR VPWR _08690_ sky130_fd_sc_hd__o211a_1
X_11659_ _07450_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__08500_ _08500_ VGND VGND VPWR VPWR clknet_0__08500_ sky130_fd_sc_hd__clkbuf_16
X_13547__936 clknet_1_1__leaf__08439_ VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__inv_2
XFILLER_0_80_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17166_ CPU.registerFile\[20\]\[28\] CPU.registerFile\[21\]\[28\] _03737_ VGND VGND
+ VPWR VPWR _04865_ sky130_fd_sc_hd__mux2_1
X_14378_ CPU.registerFile\[8\]\[1\] _08526_ _08621_ _08622_ VGND VGND VPWR VPWR _08623_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold906 CPU.registerFile\[11\]\[27\] VGND VGND VPWR VPWR net2203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16117_ _03735_ _03836_ _03841_ _03755_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__o211a_1
Xhold917 CPU.registerFile\[17\]\[18\] VGND VGND VPWR VPWR net2214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold928 CPU.registerFile\[23\]\[13\] VGND VGND VPWR VPWR net2225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold939 CPU.registerFile\[7\]\[17\] VGND VGND VPWR VPWR net2236 sky130_fd_sc_hd__dlygate4sd3_1
X_17097_ _04579_ _04580_ CPU.registerFile\[17\]\[26\] VGND VGND VPWR VPWR _04798_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__08362_ _08362_ VGND VGND VPWR VPWR clknet_0__08362_ sky130_fd_sc_hd__clkbuf_16
X_16048_ _06109_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__clkbuf_4
X_17999_ net1010 _01527_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09422_ _05410_ _05506_ _05507_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__a21oi_1
X_09353_ _05585_ _05589_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09284_ CPU.state\[3\] CPU.state\[2\] VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__nor2_2
XFILLER_0_129_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08999_ _05349_ _05350_ VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__or2_2
X_10961_ mapped_spi_flash.cmd_addr\[19\] _05641_ _07009_ VGND VGND VPWR VPWR _07012_
+ sky130_fd_sc_hd__mux2_1
X_12700_ _06624_ net2623 _08040_ VGND VGND VPWR VPWR _08044_ sky130_fd_sc_hd__mux2_1
X_10892_ CPU.aluIn1\[4\] _06958_ _06880_ VGND VGND VPWR VPWR _06959_ sky130_fd_sc_hd__mux2_1
X_12631_ _08007_ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15350_ _03202_ _03394_ _03398_ _03406_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__a31o_1
X_12562_ net2419 _07337_ _07968_ VGND VGND VPWR VPWR _07971_ sky130_fd_sc_hd__mux2_1
X_15824__573 clknet_1_0__leaf__03678_ VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__inv_2
X_13351__847 clknet_1_1__leaf__08367_ VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__inv_2
XFILLER_0_108_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15898__641 clknet_1_0__leaf__03684_ VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__inv_2
X_14301_ _06059_ VGND VGND VPWR VPWR _08547_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11513_ _07371_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__clkbuf_1
X_15281_ CPU.registerFile\[10\]\[23\] CPU.registerFile\[11\]\[23\] _03183_ VGND VGND
+ VPWR VPWR _03340_ sky130_fd_sc_hd__mux2_1
X_12493_ net2059 _07337_ _07931_ VGND VGND VPWR VPWR _07934_ sky130_fd_sc_hd__mux2_1
X_17020_ _04479_ _04718_ _04722_ _04446_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11444_ net2150 _07324_ _07312_ VGND VGND VPWR VPWR _07325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11375_ _07284_ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13996__151 clknet_1_1__leaf__08483_ VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__inv_2
X_13114_ net1448 VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__inv_2
X_10326_ _06608_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__clkbuf_1
X_18971_ net745 _02491_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ net1601 VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__clkbuf_1
X_17922_ clknet_leaf_26_clk _01450_ VGND VGND VPWR VPWR CPU.Bimm\[9\] sky130_fd_sc_hd__dfxtp_4
X_10257_ net2157 _06032_ _06558_ VGND VGND VPWR VPWR _06568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10188_ _05841_ _06333_ _05693_ VGND VGND VPWR VPWR _06510_ sky130_fd_sc_hd__mux2_1
X_17853_ net933 _01415_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_16804_ CPU.registerFile\[13\]\[19\] _04380_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__or2_1
X_14996_ _08857_ _03059_ _03061_ _02903_ VGND VGND VPWR VPWR _03062_ sky130_fd_sc_hd__a211o_1
X_17784_ net864 _01346_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_16735_ _04441_ _04442_ _04444_ _04208_ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__a211o_1
X_16666_ CPU.registerFile\[8\]\[16\] _04101_ _04102_ _04376_ VGND VGND VPWR VPWR _04377_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18405_ net226 _01933_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_12829_ _08113_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__clkbuf_1
X_16597_ _03985_ _03986_ CPU.registerFile\[1\]\[14\] VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18336_ net157 _01864_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_15548_ _03591_ _03599_ _05861_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18267_ net1278 _01795_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15479_ CPU.registerFile\[17\]\[29\] _08528_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17218_ CPU.registerFile\[12\]\[30\] _03694_ _03763_ _04914_ VGND VGND VPWR VPWR
+ _04915_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18198_ net1209 net1309 VGND VGND VPWR VPWR mapped_spi_ram.snd_bitcount\[5\] sky130_fd_sc_hd__dfxtp_1
X_13829__1190 clknet_1_0__leaf__08467_ VGND VGND VPWR VPWR net1246 sky130_fd_sc_hd__inv_2
Xhold703 CPU.registerFile\[7\]\[21\] VGND VGND VPWR VPWR net2000 sky130_fd_sc_hd__dlygate4sd3_1
X_17149_ CPU.registerFile\[5\]\[28\] CPU.registerFile\[4\]\[28\] _03697_ VGND VGND
+ VPWR VPWR _04848_ sky130_fd_sc_hd__mux2_1
Xhold714 CPU.registerFile\[21\]\[30\] VGND VGND VPWR VPWR net2011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold725 CPU.registerFile\[30\]\[8\] VGND VGND VPWR VPWR net2022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold736 CPU.registerFile\[30\]\[9\] VGND VGND VPWR VPWR net2033 sky130_fd_sc_hd__dlygate4sd3_1
X_13328__827 clknet_1_1__leaf__08364_ VGND VGND VPWR VPWR net883 sky130_fd_sc_hd__inv_2
Xhold747 CPU.registerFile\[18\]\[15\] VGND VGND VPWR VPWR net2044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 CPU.registerFile\[24\]\[0\] VGND VGND VPWR VPWR net2055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold769 CPU.registerFile\[20\]\[12\] VGND VGND VPWR VPWR net2066 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ _05309_ _05749_ VGND VGND VPWR VPWR _06302_ sky130_fd_sc_hd__nor2_1
Xclkbuf_0__08345_ _08345_ VGND VGND VPWR VPWR clknet_0__08345_ sky130_fd_sc_hd__clkbuf_16
X_08922_ CPU.Iimm\[1\] _05244_ _05273_ CPU.aluIn1\[1\] VGND VGND VPWR VPWR _05274_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09405_ _05413_ _05523_ _05755_ _05517_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_94_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09336_ net1540 VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13713__1085 clknet_1_0__leaf__08456_ VGND VGND VPWR VPWR net1141 sky130_fd_sc_hd__inv_2
XFILLER_0_7_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09267_ CPU.aluIn1\[9\] CPU.Bimm\[9\] CPU.Bimm\[8\] CPU.aluIn1\[8\] VGND VGND VPWR
+ VPWR _05619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14123__264 clknet_1_1__leaf__08497_ VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__inv_2
XFILLER_0_35_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09198_ _05549_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11160_ _06854_ VGND VGND VPWR VPWR _07163_ sky130_fd_sc_hd__buf_4
XFILLER_0_31_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10111_ _05284_ _05285_ _05528_ _06436_ VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__o22a_1
X_11091_ mapped_spi_flash.snd_bitcount\[2\] _07118_ VGND VGND VPWR VPWR _07119_ sky130_fd_sc_hd__nor2_1
X_10042_ _05884_ _06369_ VGND VGND VPWR VPWR _06370_ sky130_fd_sc_hd__nor2_1
Xhold30 mapped_spi_flash.rcv_data\[11\] VGND VGND VPWR VPWR net1327 sky130_fd_sc_hd__clkbuf_2
X_15711__504 clknet_1_0__leaf__03649_ VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__inv_2
Xhold41 mapped_spi_flash.rcv_data\[3\] VGND VGND VPWR VPWR net1338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 mapped_spi_ram.cmd_addr\[6\] VGND VGND VPWR VPWR net1349 sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ _02751_ _02916_ _02918_ _02759_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__a211o_1
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold63 mapped_spi_ram.cmd_addr\[5\] VGND VGND VPWR VPWR net1360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 mapped_spi_ram.cmd_addr\[28\] VGND VGND VPWR VPWR net1371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 _05785_ VGND VGND VPWR VPWR net1382 sky130_fd_sc_hd__buf_1
Xhold96 mapped_spi_flash.clk_div VGND VGND VPWR VPWR net1393 sky130_fd_sc_hd__dlygate4sd3_1
X_14781_ _02849_ _02850_ _02851_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__mux2_1
X_11993_ _07628_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__clkbuf_1
X_16520_ CPU.registerFile\[0\]\[12\] _04233_ _04068_ _04234_ VGND VGND VPWR VPWR _04235_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10944_ _06985_ VGND VGND VPWR VPWR _07000_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16451_ _04037_ _04164_ _04167_ _03803_ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__a211o_1
XFILLER_0_128_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10875_ CPU.aluReg\[9\] CPU.aluReg\[7\] _06939_ VGND VGND VPWR VPWR _06946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15402_ _03230_ _03453_ _03457_ _03151_ VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__o211a_1
X_12614_ _07998_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__clkbuf_1
X_19170_ clknet_leaf_5_clk net2625 VGND VGND VPWR VPWR per_uart.uart0.rx_busy sky130_fd_sc_hd__dfxtp_1
X_16382_ CPU.registerFile\[10\]\[9\] CPU.registerFile\[11\]\[9\] _03931_ VGND VGND
+ VPWR VPWR _04100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18121_ net1132 _01649_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15333_ net1580 _03201_ _03389_ _03390_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__o211a_1
X_12545_ net2512 _07320_ _07957_ VGND VGND VPWR VPWR _07962_ sky130_fd_sc_hd__mux2_1
X_18052_ net1063 _01580_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15264_ _03156_ _03320_ _03322_ _03163_ VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__a211o_1
XFILLER_0_151_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12476_ net2203 _07320_ _07920_ VGND VGND VPWR VPWR _07925_ sky130_fd_sc_hd__mux2_1
X_17003_ _04419_ _04703_ _04705_ _04383_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_667 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11427_ _07313_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__03641_ clknet_0__03641_ VGND VGND VPWR VPWR clknet_1_1__leaf__03641_
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_5 CPU.mem_wdata\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15195_ _03253_ _03254_ _03255_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11358_ net1692 _05767_ _07274_ VGND VGND VPWR VPWR _07276_ sky130_fd_sc_hd__mux2_1
X_10309_ _06596_ VGND VGND VPWR VPWR _06597_ sky130_fd_sc_hd__buf_4
X_18954_ net728 _02474_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11289_ _07239_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__clkbuf_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ CPU.registerFile\[4\]\[30\] net1347 _08217_ VGND VGND VPWR VPWR _08219_ sky130_fd_sc_hd__mux2_1
X_17905_ clknet_leaf_24_clk _01433_ VGND VGND VPWR VPWR CPU.Jimm\[12\] sky130_fd_sc_hd__dfxtp_4
X_18885_ net659 _02405_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_15651__451 clknet_1_1__leaf__03642_ VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__inv_2
X_17836_ net916 _01398_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_17767_ net847 _01329_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14979_ CPU.registerFile\[30\]\[16\] CPU.registerFile\[31\]\[16\] _02887_ VGND VGND
+ VPWR VPWR _03045_ sky130_fd_sc_hd__mux2_1
X_16718_ _03744_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__buf_4
XFILLER_0_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17698_ CPU.mem_wdata\[2\] per_uart.d_in_uart\[2\] _05218_ VGND VGND VPWR VPWR _05223_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16649_ _04075_ _04356_ _04360_ _04042_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09121_ _05328_ _05471_ _05472_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__a21o_1
XFILLER_0_162_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18319_ net140 _01847_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_919 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09052_ _05385_ _05388_ _05403_ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold500 CPU.registerFile\[28\]\[27\] VGND VGND VPWR VPWR net1797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 CPU.registerFile\[5\]\[15\] VGND VGND VPWR VPWR net1808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 CPU.registerFile\[30\]\[21\] VGND VGND VPWR VPWR net1819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold533 CPU.registerFile\[22\]\[3\] VGND VGND VPWR VPWR net1830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold544 CPU.registerFile\[22\]\[19\] VGND VGND VPWR VPWR net1841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 CPU.registerFile\[9\]\[6\] VGND VGND VPWR VPWR net1852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 CPU.registerFile\[5\]\[12\] VGND VGND VPWR VPWR net1863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 CPU.registerFile\[10\]\[21\] VGND VGND VPWR VPWR net1874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 CPU.registerFile\[30\]\[3\] VGND VGND VPWR VPWR net1885 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ _05912_ _06282_ _06285_ VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold599 CPU.registerFile\[15\]\[10\] VGND VGND VPWR VPWR net1896 sky130_fd_sc_hd__dlygate4sd3_1
X_13380__873 clknet_1_1__leaf__08370_ VGND VGND VPWR VPWR net929 sky130_fd_sc_hd__inv_2
X_08905_ CPU.rs2\[28\] _05247_ _05251_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ CPU.PC\[14\] _05888_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__nor2_1
Xhold1200 CPU.registerFile\[4\]\[21\] VGND VGND VPWR VPWR net2497 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1211 CPU.registerFile\[8\]\[13\] VGND VGND VPWR VPWR net2508 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1222 CPU.registerFile\[1\]\[31\] VGND VGND VPWR VPWR net2519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1233 CPU.registerFile\[25\]\[21\] VGND VGND VPWR VPWR net2530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 CPU.registerFile\[12\]\[6\] VGND VGND VPWR VPWR net2541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1255 CPU.registerFile\[25\]\[17\] VGND VGND VPWR VPWR net2552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 CPU.registerFile\[24\]\[31\] VGND VGND VPWR VPWR net2563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1277 _05177_ VGND VGND VPWR VPWR net2574 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1288 CPU.registerFile\[9\]\[10\] VGND VGND VPWR VPWR net2585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 CPU.registerFile\[1\]\[24\] VGND VGND VPWR VPWR net2596 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10660_ net2488 _06292_ _06799_ VGND VGND VPWR VPWR _06800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09319_ CPU.PC\[17\] _05636_ _05669_ _05670_ _05235_ VGND VGND VPWR VPWR _05671_
+ sky130_fd_sc_hd__o221a_1
X_10591_ _06762_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12330_ _06594_ _07488_ VGND VGND VPWR VPWR _07847_ sky130_fd_sc_hd__nand2_4
X_12261_ net1556 _07800_ VGND VGND VPWR VPWR _07804_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11212_ _07197_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__clkbuf_1
X_15936__674 clknet_1_1__leaf__03689_ VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__inv_2
Xoutput7 net7 VGND VGND VPWR VPWR spi_clk sky130_fd_sc_hd__clkbuf_4
X_12192_ mapped_spi_ram.cmd_addr\[0\] _07749_ _07706_ CPU.mem_wdata\[1\] _07695_ VGND
+ VGND VPWR VPWR _07756_ sky130_fd_sc_hd__a221o_1
X_11143_ net1599 _07147_ _07153_ _07151_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__o211a_1
X_13795__1159 clknet_1_1__leaf__08464_ VGND VGND VPWR VPWR net1215 sky130_fd_sc_hd__inv_2
XFILLER_0_102_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11074_ mapped_spi_flash.cmd_addr\[1\] _06983_ _06984_ mapped_spi_flash.cmd_addr\[0\]
+ VGND VGND VPWR VPWR _07106_ sky130_fd_sc_hd__a22o_1
X_14902_ CPU.registerFile\[24\]\[14\] _02928_ _02969_ _02771_ VGND VGND VPWR VPWR
+ _02970_ sky130_fd_sc_hd__o211a_1
X_10025_ _05970_ _05946_ VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__and2b_1
X_18670_ net459 _02194_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_17621_ _05169_ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14833_ _08418_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__clkbuf_4
X_14764_ _02826_ _02829_ _02835_ _02746_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__o211a_1
X_17552_ per_uart.uart0.tx_count16\[3\] _03658_ _05119_ VGND VGND VPWR VPWR _05120_
+ sky130_fd_sc_hd__or3_2
X_11976_ _07619_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16503_ _04210_ _04218_ _04138_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__o21a_1
XFILLER_0_156_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17483_ _05022_ _06277_ _08256_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__o21ai_1
X_10927_ mapped_spi_flash.cmd_addr\[30\] _06983_ _06985_ mapped_spi_flash.cmd_addr\[29\]
+ VGND VGND VPWR VPWR _06988_ sky130_fd_sc_hd__a22o_1
X_14695_ _06062_ VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__buf_4
XFILLER_0_39_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16434_ CPU.registerFile\[6\]\[10\] CPU.registerFile\[7\]\[10\] _04022_ VGND VGND
+ VPWR VPWR _04151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10858_ CPU.aluReg\[13\] CPU.aluReg\[11\] _06906_ VGND VGND VPWR VPWR _06933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15681__477 clknet_1_1__leaf__03646_ VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__inv_2
XFILLER_0_128_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17323__736 clknet_1_1__leaf__04982_ VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__inv_2
XFILLER_0_156_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16365_ _04037_ _04079_ _04083_ _03803_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__a211o_1
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19153_ clknet_leaf_4_clk net1452 VGND VGND VPWR VPWR per_uart.uart0.txd_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10789_ _06860_ VGND VGND VPWR VPWR _06880_ sky130_fd_sc_hd__buf_4
XFILLER_0_143_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15316_ _03372_ _03373_ _08541_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__mux2_1
X_18104_ net1115 _01632_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_12528_ net1993 _07372_ _07942_ VGND VGND VPWR VPWR _07952_ sky130_fd_sc_hd__mux2_1
X_16296_ CPU.registerFile\[15\]\[7\] CPU.registerFile\[14\]\[7\] _03705_ VGND VGND
+ VPWR VPWR _04016_ sky130_fd_sc_hd__mux2_1
X_19084_ clknet_leaf_0_clk _02604_ VGND VGND VPWR VPWR per_uart.uart0.rxd_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15247_ _08418_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__clkbuf_4
X_18035_ net1046 _01563_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12459_ _07915_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__clkbuf_1
X_15178_ _03230_ _03233_ _03239_ _03151_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0__03655_ _03655_ VGND VGND VPWR VPWR clknet_0__03655_ sky130_fd_sc_hd__clkbuf_16
X_18937_ net711 _02457_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_09670_ _06012_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__buf_4
X_18868_ net642 _02388_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13712__1084 clknet_1_0__leaf__08456_ VGND VGND VPWR VPWR net1140 sky130_fd_sc_hd__inv_2
X_17819_ net899 _01381_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_18799_ net588 _02323_ VGND VGND VPWR VPWR CPU.aluReg\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17298__713 clknet_1_0__leaf__04980_ VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__inv_2
XFILLER_0_116_943 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09104_ CPU.aluIn1\[13\] _05322_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09035_ CPU.rs2\[24\] _05247_ _05251_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold330 CPU.rs2\[19\] VGND VGND VPWR VPWR net1627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 CPU.rs2\[20\] VGND VGND VPWR VPWR net1638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 net7 VGND VGND VPWR VPWR net1649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 _05181_ VGND VGND VPWR VPWR net1660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold374 _05173_ VGND VGND VPWR VPWR net1671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 CPU.registerFile\[5\]\[19\] VGND VGND VPWR VPWR net1682 sky130_fd_sc_hd__dlygate4sd3_1
X_14235__365 clknet_1_1__leaf__08508_ VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__inv_2
Xhold396 CPU.registerFile\[6\]\[3\] VGND VGND VPWR VPWR net1693 sky130_fd_sc_hd__dlygate4sd3_1
X_09937_ _05313_ _05523_ _05749_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__o21ai_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _05693_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__clkbuf_4
Xhold1030 CPU.registerFile\[14\]\[8\] VGND VGND VPWR VPWR net2327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 CPU.registerFile\[2\]\[27\] VGND VGND VPWR VPWR net2338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1052 CPU.registerFile\[3\]\[6\] VGND VGND VPWR VPWR net2349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1063 CPU.registerFile\[12\]\[30\] VGND VGND VPWR VPWR net2360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 CPU.registerFile\[27\]\[26\] VGND VGND VPWR VPWR net2371 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ _05891_ _06136_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__or2_1
Xhold1085 CPU.registerFile\[2\]\[24\] VGND VGND VPWR VPWR net2382 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _07542_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__clkbuf_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1096 per_uart.uart0.tx_count16\[0\] VGND VGND VPWR VPWR net2393 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03644_ clknet_0__03644_ VGND VGND VPWR VPWR clknet_1_0__leaf__03644_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _06626_ net2174 _07501_ VGND VGND VPWR VPWR _07506_ sky130_fd_sc_hd__mux2_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14129__270 clknet_1_0__leaf__08497_ VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__inv_2
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ net2401 _06083_ _06827_ VGND VGND VPWR VPWR _06829_ sky130_fd_sc_hd__mux2_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _08532_ VGND VGND VPWR VPWR _08722_ sky130_fd_sc_hd__clkbuf_4
X_11692_ net2177 _07341_ _07464_ VGND VGND VPWR VPWR _07469_ sky130_fd_sc_hd__mux2_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13431_ mapped_spi_flash.rcv_data\[8\] _05859_ _06147_ VGND VGND VPWR VPWR _08396_
+ sky130_fd_sc_hd__a21o_4
XFILLER_0_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10643_ net2364 _06106_ _06788_ VGND VGND VPWR VPWR _06791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16150_ CPU.registerFile\[28\]\[3\] CPU.registerFile\[29\]\[3\] _03739_ VGND VGND
+ VPWR VPWR _03874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10574_ _06753_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__clkbuf_1
X_15101_ _03156_ _03158_ _03162_ _03163_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12313_ _07833_ net1311 net1303 VGND VGND VPWR VPWR _07836_ sky130_fd_sc_hd__mux2_1
X_16081_ CPU.registerFile\[20\]\[1\] CPU.registerFile\[21\]\[1\] _03761_ VGND VGND
+ VPWR VPWR _03807_ sky130_fd_sc_hd__mux2_1
X_15032_ _03095_ _03096_ _02937_ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__mux2_1
X_12244_ net1373 _07787_ VGND VGND VPWR VPWR _07794_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15717__510 clknet_1_1__leaf__03649_ VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__inv_2
X_12175_ mapped_spi_ram.cmd_addr\[7\] _05714_ _07724_ VGND VGND VPWR VPWR _07746_
+ sky130_fd_sc_hd__mux2_1
X_11126_ net1356 _07133_ _07143_ _07138_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16983_ _04441_ _04684_ _04686_ _04612_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__a211o_1
X_18722_ net511 _02246_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[22\] sky130_fd_sc_hd__dfxtp_1
X_11057_ net1534 _07054_ _07093_ _07069_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10008_ net2564 _06337_ _06293_ VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__mux2_1
X_18653_ clknet_leaf_11_clk _02177_ VGND VGND VPWR VPWR CPU.rs2\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17604_ per_uart.d_in_uart\[1\] _05134_ _05157_ per_uart.uart0.txd_reg\[2\] VGND
+ VGND VPWR VPWR _05160_ sky130_fd_sc_hd__o22a_1
X_14816_ _08837_ _02883_ _02885_ _08802_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__a211o_1
X_18584_ net405 net41 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15796_ _08349_ _03666_ _03661_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17535_ _05104_ _05105_ _05058_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14747_ CPU.registerFile\[13\]\[10\] CPU.registerFile\[12\]\[10\] _08693_ VGND VGND
+ VPWR VPWR _02819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11959_ _06620_ net2440 _07609_ VGND VGND VPWR VPWR _07611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17466_ _08379_ _05017_ _06328_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__o21bai_1
X_14678_ _08414_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16417_ CPU.registerFile\[16\]\[9\] _03848_ _04090_ _04134_ VGND VGND VPWR VPWR _04135_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19136_ clknet_leaf_15_clk _02656_ VGND VGND VPWR VPWR CPU.PC\[18\] sky130_fd_sc_hd__dfxtp_2
X_16348_ CPU.registerFile\[2\]\[8\] CPU.registerFile\[3\]\[8\] _04027_ VGND VGND VPWR
+ VPWR _04067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16279_ CPU.registerFile\[22\]\[6\] CPU.registerFile\[23\]\[6\] _03958_ VGND VGND
+ VPWR VPWR _04000_ sky130_fd_sc_hd__mux2_1
X_19067_ net59 _02587_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08493_ clknet_0__08493_ VGND VGND VPWR VPWR clknet_1_1__leaf__08493_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18018_ net1029 _01546_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__03638_ _03638_ VGND VGND VPWR VPWR clknet_0__03638_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09722_ _06062_ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__clkbuf_4
X_18235__19 VGND VGND VPWR VPWR _18235__19/HI net19 sky130_fd_sc_hd__conb_1
X_09653_ CPU.PC\[20\] _05996_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09584_ CPU.PC\[18\] _05926_ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__nor2_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17349__10 clknet_1_0__leaf__04984_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__inv_2
XFILLER_0_93_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13794__1158 clknet_1_1__leaf__08464_ VGND VGND VPWR VPWR net1214 sky130_fd_sc_hd__inv_2
XFILLER_0_147_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13232__754 clknet_1_1__leaf__08342_ VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__inv_2
XFILLER_0_162_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09018_ _05363_ _05369_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__nor2_1
X_10290_ _06585_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold160 _02259_ VGND VGND VPWR VPWR net1457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 mapped_spi_ram.rcv_data\[3\] VGND VGND VPWR VPWR net1468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _02679_ VGND VGND VPWR VPWR net1479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 mapped_spi_ram.cmd_addr\[10\] VGND VGND VPWR VPWR net1490 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12931_ _08144_ VGND VGND VPWR VPWR _08167_ sky130_fd_sc_hd__buf_4
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ _08130_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__clkbuf_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _07533_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__clkbuf_1
X_14601_ CPU.registerFile\[21\]\[7\] _08718_ VGND VGND VPWR VPWR _08840_ sky130_fd_sc_hd__or2_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _08567_ _08569_ CPU.registerFile\[1\]\[31\] VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__a21o_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _06649_ net2216 _08087_ VGND VGND VPWR VPWR _08093_ sky130_fd_sc_hd__mux2_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ CPU.registerFile\[13\]\[5\] CPU.registerFile\[12\]\[5\] _08693_ VGND VGND
+ VPWR VPWR _08773_ sky130_fd_sc_hd__mux2_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _06609_ net2350 _07490_ VGND VGND VPWR VPWR _07497_ sky130_fd_sc_hd__mux2_1
X_14062__210 clknet_1_1__leaf__08490_ VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__inv_2
XFILLER_0_139_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17251_ _03703_ _04944_ _04946_ _06142_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__a211o_1
X_14463_ _08410_ VGND VGND VPWR VPWR _08706_ sky130_fd_sc_hd__clkbuf_4
X_11675_ net2259 _07324_ _07453_ VGND VGND VPWR VPWR _07460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13414_ _05738_ _06333_ _00000_ VGND VGND VPWR VPWR _08386_ sky130_fd_sc_hd__mux2_1
X_16202_ _03770_ _03771_ CPU.registerFile\[17\]\[4\] VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__a21o_1
X_17182_ CPU.registerFile\[12\]\[29\] _03694_ _03763_ _04879_ VGND VGND VPWR VPWR
+ _04880_ sky130_fd_sc_hd__o211a_1
X_10626_ net2384 _05825_ _06777_ VGND VGND VPWR VPWR _06782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14394_ CPU.registerFile\[17\]\[2\] _06456_ VGND VGND VPWR VPWR _08638_ sky130_fd_sc_hd__or2_1
X_13711__1083 clknet_1_0__leaf__08456_ VGND VGND VPWR VPWR net1139 sky130_fd_sc_hd__inv_2
X_16133_ CPU.registerFile\[9\]\[3\] _03698_ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__or2_1
X_13345_ clknet_1_1__leaf__08366_ VGND VGND VPWR VPWR _08367_ sky130_fd_sc_hd__buf_1
X_10557_ _06744_ VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16064_ CPU.registerFile\[2\]\[1\] CPU.registerFile\[3\]\[1\] _03693_ VGND VGND VPWR
+ VPWR _03790_ sky130_fd_sc_hd__mux2_1
X_13276_ per_uart.uart0.enable16_counter\[12\] _08356_ VGND VGND VPWR VPWR _08357_
+ sky130_fd_sc_hd__or2_1
X_10488_ _06707_ VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__clkbuf_1
X_15015_ _08526_ VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__clkbuf_4
X_12227_ _07687_ _07779_ _07782_ VGND VGND VPWR VPWR _07783_ sky130_fd_sc_hd__or3b_1
XFILLER_0_121_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12158_ _07715_ _07733_ VGND VGND VPWR VPWR _07734_ sky130_fd_sc_hd__or2_1
X_11109_ _07132_ VGND VGND VPWR VPWR _07133_ sky130_fd_sc_hd__clkbuf_4
X_16966_ CPU.registerFile\[12\]\[23\] _04421_ _04422_ _04669_ VGND VGND VPWR VPWR
+ _04670_ sky130_fd_sc_hd__o211a_1
X_12089_ _07001_ net2649 _07198_ VGND VGND VPWR VPWR _07685_ sky130_fd_sc_hd__and3_1
X_18705_ net494 _02229_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[5\] sky130_fd_sc_hd__dfxtp_1
X_16897_ _04305_ _04598_ _04602_ _04476_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__o211a_1
X_18636_ clknet_leaf_17_clk _02160_ VGND VGND VPWR VPWR CPU.rs2\[8\] sky130_fd_sc_hd__dfxtp_1
X_18567_ net388 net24 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17518_ _05075_ _05025_ _06121_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__o21bai_1
X_18498_ net319 _02022_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17449_ _08334_ _06432_ _08255_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19119_ net102 _02639_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__08476_ clknet_0__08476_ VGND VGND VPWR VPWR clknet_1_1__leaf__08476_
+ sky130_fd_sc_hd__clkbuf_16
X_13524__915 clknet_1_1__leaf__08437_ VGND VGND VPWR VPWR net971 sky130_fd_sc_hd__inv_2
XFILLER_0_112_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09705_ _05369_ _05532_ _05535_ CPU.aluReg\[21\] _06046_ VGND VGND VPWR VPWR _06047_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09636_ CPU.Jimm\[14\] _05921_ _05923_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__a21o_1
X_09567_ _05910_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09498_ _05385_ _05532_ _05535_ CPU.aluReg\[25\] VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11460_ net1737 _07335_ _07333_ VGND VGND VPWR VPWR _07336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10411_ _06666_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11391_ net1821 _06224_ _07285_ VGND VGND VPWR VPWR _07293_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__05013_ clknet_0__05013_ VGND VGND VPWR VPWR clknet_1_0__leaf__05013_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_162_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13130_ _08271_ _08272_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__nor2_1
X_10342_ _06619_ VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_696 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13061_ CPU.registerFile\[4\]\[14\] net1417 _08228_ VGND VGND VPWR VPWR _08236_ sky130_fd_sc_hd__mux2_1
X_10273_ _06576_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__clkbuf_1
X_12012_ _07639_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__clkbuf_1
X_13921__82 clknet_1_0__leaf__08477_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__inv_2
X_16820_ _04525_ _04527_ _04279_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__mux2_1
X_16751_ _03697_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__buf_2
XFILLER_0_45_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12914_ _08158_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__clkbuf_1
X_16682_ _04347_ _04388_ _04392_ _04117_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_0__f__08496_ clknet_0__08496_ VGND VGND VPWR VPWR clknet_1_0__leaf__08496_
+ sky130_fd_sc_hd__clkbuf_16
X_18421_ net242 _01949_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12845_ _06083_ net2358 _08120_ VGND VGND VPWR VPWR _08122_ sky130_fd_sc_hd__mux2_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ net173 _01880_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _08566_ _08568_ CPU.registerFile\[25\]\[31\] VGND VGND VPWR VPWR _03615_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _06632_ net2210 _08076_ VGND VGND VPWR VPWR _08084_ sky130_fd_sc_hd__mux2_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11727_ net2270 _07376_ _07452_ VGND VGND VPWR VPWR _07487_ sky130_fd_sc_hd__mux2_1
X_14515_ _08522_ VGND VGND VPWR VPWR _08756_ sky130_fd_sc_hd__buf_4
X_15495_ CPU.registerFile\[15\]\[29\] CPU.registerFile\[14\]\[29\] _08560_ VGND VGND
+ VPWR VPWR _03548_ sky130_fd_sc_hd__mux2_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18283_ net1294 _01811_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17234_ CPU.registerFile\[24\]\[30\] _03724_ _03725_ _04930_ VGND VGND VPWR VPWR
+ _04931_ sky130_fd_sc_hd__o211a_1
X_11658_ net2292 _07376_ _07415_ VGND VGND VPWR VPWR _07450_ sky130_fd_sc_hd__mux2_1
X_14446_ _08543_ _08685_ _08688_ _08552_ VGND VGND VPWR VPWR _08689_ sky130_fd_sc_hd__a211o_1
XFILLER_0_37_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10609_ _06771_ VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__clkbuf_1
X_14377_ _08549_ VGND VGND VPWR VPWR _08622_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17165_ CPU.registerFile\[22\]\[28\] CPU.registerFile\[23\]\[28\] _03761_ VGND VGND
+ VPWR VPWR _04864_ sky130_fd_sc_hd__mux2_1
X_15875__620 clknet_1_1__leaf__03682_ VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__inv_2
X_11589_ net1702 _07376_ _07378_ VGND VGND VPWR VPWR _07413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold907 CPU.registerFile\[17\]\[9\] VGND VGND VPWR VPWR net2204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold918 CPU.registerFile\[12\]\[11\] VGND VGND VPWR VPWR net2215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16116_ _03702_ _03838_ _03840_ _03803_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__a211o_1
X_17096_ CPU.registerFile\[19\]\[26\] CPU.registerFile\[18\]\[26\] _03745_ VGND VGND
+ VPWR VPWR _04797_ sky130_fd_sc_hd__mux2_1
Xhold929 CPU.registerFile\[21\]\[22\] VGND VGND VPWR VPWR net2226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08361_ _08361_ VGND VGND VPWR VPWR clknet_0__08361_ sky130_fd_sc_hd__clkbuf_16
X_16047_ _03766_ _03768_ _03773_ _06142_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__a211o_1
X_13973__130 clknet_1_0__leaf__08481_ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__inv_2
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13793__1157 clknet_1_1__leaf__08464_ VGND VGND VPWR VPWR net1213 sky130_fd_sc_hd__inv_2
X_17998_ net1009 _01526_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_16949_ _04652_ _04653_ _04365_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__mux2_1
X_14069__216 clknet_1_0__leaf__08491_ VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__inv_2
XFILLER_0_79_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09421_ _05255_ _05522_ _05749_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__o21a_1
X_18619_ net440 _02143_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17421__42 clknet_1_1__leaf__05015_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__inv_2
X_09352_ _05558_ _05701_ _05702_ _05703_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09283_ _05559_ _05560_ _05633_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15776__562 clknet_1_1__leaf__03656_ VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__inv_2
XFILLER_0_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__08459_ clknet_0__08459_ VGND VGND VPWR VPWR clknet_1_1__leaf__08459_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13305__806 clknet_1_1__leaf__08362_ VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__inv_2
X_15930__669 clknet_1_0__leaf__03688_ VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__inv_2
X_08998_ CPU.aluIn1\[19\] _05348_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13710__1082 clknet_1_0__leaf__08456_ VGND VGND VPWR VPWR net1138 sky130_fd_sc_hd__inv_2
X_10960_ net1546 _07007_ _07011_ _06856_ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13494__888 clknet_1_1__leaf__08434_ VGND VGND VPWR VPWR net944 sky130_fd_sc_hd__inv_2
X_09619_ _05951_ _05961_ _05962_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__a21o_1
X_10891_ CPU.aluReg\[5\] CPU.aluReg\[3\] _06939_ VGND VGND VPWR VPWR _06958_ sky130_fd_sc_hd__mux2_1
X_12630_ _06622_ net1781 _08004_ VGND VGND VPWR VPWR _08007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13238__760 clknet_1_0__leaf__08342_ VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__inv_2
X_12561_ _07970_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14300_ _06058_ VGND VGND VPWR VPWR _08546_ sky130_fd_sc_hd__buf_4
X_11512_ net1898 _07370_ _07354_ VGND VGND VPWR VPWR _07371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15280_ _03337_ _03338_ _08541_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12492_ _07933_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14231_ clknet_1_0__leaf__08506_ VGND VGND VPWR VPWR _08508_ sky130_fd_sc_hd__buf_1
X_11443_ _05852_ VGND VGND VPWR VPWR _07324_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11374_ net1747 _06032_ _07274_ VGND VGND VPWR VPWR _07284_ sky130_fd_sc_hd__mux2_1
X_14174__311 clknet_1_1__leaf__08501_ VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__inv_2
X_13113_ _08263_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__clkbuf_1
X_10325_ _06607_ net1771 _06597_ VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__mux2_1
X_18970_ net744 _02490_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ CPU.registerFile\[4\]\[22\] _06031_ _08217_ VGND VGND VPWR VPWR _08227_ sky130_fd_sc_hd__mux2_1
X_17921_ clknet_leaf_26_clk _01449_ VGND VGND VPWR VPWR CPU.Bimm\[8\] sky130_fd_sc_hd__dfxtp_4
X_10256_ _06567_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__clkbuf_1
X_17852_ net932 _01414_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_10187_ _06509_ VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__clkbuf_1
X_16803_ CPU.registerFile\[15\]\[19\] CPU.registerFile\[14\]\[19\] _04146_ VGND VGND
+ VPWR VPWR _04511_ sky130_fd_sc_hd__mux2_1
X_17783_ net863 _01345_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_14995_ CPU.registerFile\[8\]\[16\] _03018_ _03060_ _02864_ VGND VGND VPWR VPWR _03061_
+ sky130_fd_sc_hd__o211a_1
X_16734_ CPU.registerFile\[24\]\[17\] _04319_ _04165_ _04443_ VGND VGND VPWR VPWR
+ _04444_ sky130_fd_sc_hd__o211a_1
X_16665_ CPU.registerFile\[9\]\[16\] _04056_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__or2_1
X_15907__649 clknet_1_1__leaf__03685_ VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__inv_2
XFILLER_0_29_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18404_ net225 _01932_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[4\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__08479_ clknet_0__08479_ VGND VGND VPWR VPWR clknet_1_0__leaf__08479_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_158_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12828_ _05805_ net2241 _08109_ VGND VGND VPWR VPWR _08113_ sky130_fd_sc_hd__mux2_1
X_16596_ CPU.registerFile\[2\]\[14\] CPU.registerFile\[3\]\[14\] _04027_ VGND VGND
+ VPWR VPWR _04309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18335_ net156 _01863_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15547_ _08557_ _03594_ _03598_ _05876_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__o211a_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _06615_ net2293 _08065_ VGND VGND VPWR VPWR _08075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18266_ net1277 _01794_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_15478_ CPU.registerFile\[19\]\[29\] CPU.registerFile\[18\]\[29\] _06456_ VGND VGND
+ VPWR VPWR _03531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17217_ CPU.registerFile\[13\]\[30\] _03767_ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14429_ _08425_ _08654_ _08672_ _08597_ VGND VGND VPWR VPWR _08673_ sky130_fd_sc_hd__a211o_1
X_18197_ net1208 _01725_ VGND VGND VPWR VPWR mapped_spi_ram.snd_bitcount\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold704 CPU.registerFile\[5\]\[17\] VGND VGND VPWR VPWR net2001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17148_ CPU.registerFile\[6\]\[28\] CPU.registerFile\[7\]\[28\] _03847_ VGND VGND
+ VPWR VPWR _04847_ sky130_fd_sc_hd__mux2_1
X_14040__190 clknet_1_1__leaf__08488_ VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__inv_2
Xhold715 CPU.registerFile\[27\]\[20\] VGND VGND VPWR VPWR net2012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 CPU.registerFile\[31\]\[31\] VGND VGND VPWR VPWR net2023 sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 CPU.registerFile\[7\]\[8\] VGND VGND VPWR VPWR net2034 sky130_fd_sc_hd__dlygate4sd3_1
X_17292__708 clknet_1_0__leaf__04979_ VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__inv_2
XFILLER_0_110_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold748 CPU.registerFile\[13\]\[14\] VGND VGND VPWR VPWR net2045 sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ _06126_ _06296_ _06300_ _05818_ VGND VGND VPWR VPWR _06301_ sky130_fd_sc_hd__o211a_1
X_17079_ CPU.registerFile\[2\]\[26\] CPU.registerFile\[3\]\[26\] _04431_ VGND VGND
+ VPWR VPWR _04780_ sky130_fd_sc_hd__mux2_1
Xhold759 CPU.registerFile\[26\]\[31\] VGND VGND VPWR VPWR net2056 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__08344_ _08344_ VGND VGND VPWR VPWR clknet_0__08344_ sky130_fd_sc_hd__clkbuf_16
X_08921_ _05240_ _05241_ _05272_ _05243_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_110_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13900__63 clknet_1_1__leaf__08475_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__inv_2
XFILLER_0_79_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09404_ _05752_ _05754_ _05424_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09335_ _05684_ _05686_ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09266_ _05600_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09197_ _05546_ _05548_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10110_ _05284_ _05285_ _05523_ VGND VGND VPWR VPWR _06436_ sky130_fd_sc_hd__a21oi_1
X_11090_ mapped_spi_flash.snd_bitcount\[1\] mapped_spi_flash.snd_bitcount\[0\] _07114_
+ VGND VGND VPWR VPWR _07118_ sky130_fd_sc_hd__or3_1
XFILLER_0_101_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10041_ CPU.PC\[6\] _05883_ CPU.PC\[7\] VGND VGND VPWR VPWR _06369_ sky130_fd_sc_hd__a21oi_1
Xhold20 _01752_ VGND VGND VPWR VPWR net1317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 _06105_ VGND VGND VPWR VPWR net1328 sky130_fd_sc_hd__buf_1
Xhold42 _05824_ VGND VGND VPWR VPWR net1339 sky130_fd_sc_hd__clkbuf_2
Xhold53 _01733_ VGND VGND VPWR VPWR net1350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 CPU.aluReg\[1\] VGND VGND VPWR VPWR net1361 sky130_fd_sc_hd__dlygate4sd3_1
X_13502__895 clknet_1_0__leaf__08435_ VGND VGND VPWR VPWR net951 sky130_fd_sc_hd__inv_2
Xhold75 mapped_spi_ram.cmd_addr\[29\] VGND VGND VPWR VPWR net1372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 _08220_ VGND VGND VPWR VPWR net1383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 _07183_ VGND VGND VPWR VPWR net1394 sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ _06653_ net2187 _07620_ VGND VGND VPWR VPWR _07628_ sky130_fd_sc_hd__mux2_1
X_14780_ _08549_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__buf_4
X_13731_ clknet_1_0__leaf__08451_ VGND VGND VPWR VPWR _08458_ sky130_fd_sc_hd__buf_1
XFILLER_0_58_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10943_ mapped_spi_flash.state\[2\] mapped_spi_flash.state\[1\] _06981_ VGND VGND
+ VPWR VPWR _06999_ sky130_fd_sc_hd__o21a_2
X_16450_ CPU.registerFile\[24\]\[10\] _03915_ _04165_ _04166_ VGND VGND VPWR VPWR
+ _04167_ sky130_fd_sc_hd__o211a_1
X_10874_ _06945_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18594__51 VGND VGND VPWR VPWR _18594__51/HI net51 sky130_fd_sc_hd__conb_1
X_15401_ _08414_ _03454_ _03456_ _03111_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__a211o_1
XFILLER_0_156_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12613_ _06605_ net2330 _07993_ VGND VGND VPWR VPWR _07998_ sky130_fd_sc_hd__mux2_1
X_17400__23 clknet_1_0__leaf__05013_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__inv_2
X_16381_ _08397_ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18120_ net1131 _01648_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_12544_ _07961_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__clkbuf_1
X_13792__1156 clknet_1_1__leaf__08464_ VGND VGND VPWR VPWR net1212 sky130_fd_sc_hd__inv_2
X_15332_ _06855_ VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18051_ net1062 _01579_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12475_ _07924_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__clkbuf_1
X_15263_ CPU.registerFile\[16\]\[23\] _03159_ _03321_ _03161_ VGND VGND VPWR VPWR
+ _03322_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14098__242 clknet_1_0__leaf__08494_ VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__inv_2
XFILLER_0_34_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17002_ CPU.registerFile\[12\]\[24\] _04421_ _04422_ _04704_ VGND VGND VPWR VPWR
+ _04705_ sky130_fd_sc_hd__o211a_1
X_11426_ net1680 _07309_ _07312_ VGND VGND VPWR VPWR _07313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__03640_ clknet_0__03640_ VGND VGND VPWR VPWR clknet_1_1__leaf__03640_
+ sky130_fd_sc_hd__clkbuf_16
X_15194_ _08549_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__buf_4
XANTENNA_6 CPU.mem_wdata\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11357_ _07275_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13730__1101 clknet_1_1__leaf__08457_ VGND VGND VPWR VPWR net1157 sky130_fd_sc_hd__inv_2
XFILLER_0_21_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10308_ _06594_ _06595_ VGND VGND VPWR VPWR _06596_ sky130_fd_sc_hd__nand2_4
X_18953_ net727 _02473_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11288_ net2014 _05734_ _07238_ VGND VGND VPWR VPWR _07239_ sky130_fd_sc_hd__mux2_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ net1411 VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__clkbuf_1
X_17904_ clknet_leaf_25_clk _01432_ VGND VGND VPWR VPWR CPU.Bimm\[4\] sky130_fd_sc_hd__dfxtp_1
X_15913__653 clknet_1_1__leaf__03687_ VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__inv_2
X_10239_ net1697 _05734_ _06558_ VGND VGND VPWR VPWR _06559_ sky130_fd_sc_hd__mux2_1
X_18884_ net658 _02404_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17835_ net915 _01397_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_17766_ net846 _01328_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_14978_ _08837_ _03040_ _03042_ _03043_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16717_ CPU.registerFile\[6\]\[17\] CPU.registerFile\[7\]\[17\] _04426_ VGND VGND
+ VPWR VPWR _04427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17697_ _05222_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16648_ _04037_ _04357_ _04359_ _04208_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13334__832 clknet_1_0__leaf__08365_ VGND VGND VPWR VPWR net888 sky130_fd_sc_hd__inv_2
XFILLER_0_146_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16579_ _03963_ _04290_ _04292_ _04006_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__a211o_1
X_09120_ _05325_ CPU.aluIn1\[15\] VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__and2b_1
X_18318_ net139 _01846_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09051_ CPU.aluIn1\[25\] _05383_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__or2_1
X_18249_ net1260 _01777_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17300__715 clknet_1_0__leaf__04980_ VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__inv_2
XFILLER_0_114_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold501 CPU.registerFile\[28\]\[11\] VGND VGND VPWR VPWR net1798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold512 CPU.registerFile\[10\]\[7\] VGND VGND VPWR VPWR net1809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold523 CPU.registerFile\[22\]\[22\] VGND VGND VPWR VPWR net1820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 CPU.registerFile\[20\]\[19\] VGND VGND VPWR VPWR net1831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold545 CPU.registerFile\[28\]\[26\] VGND VGND VPWR VPWR net1842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold556 CPU.registerFile\[22\]\[24\] VGND VGND VPWR VPWR net1853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold567 CPU.registerFile\[10\]\[17\] VGND VGND VPWR VPWR net1864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 CPU.registerFile\[18\]\[18\] VGND VGND VPWR VPWR net1875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold589 CPU.registerFile\[10\]\[25\] VGND VGND VPWR VPWR net1886 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ CPU.cycles\[11\] _05553_ _06197_ _06284_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__o2bb2a_1
X_08904_ CPU.aluIn1\[29\] _05254_ VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__nor2_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _06218_ _05983_ VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__xnor2_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1201 _08229_ VGND VGND VPWR VPWR net2498 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1212 CPU.registerFile\[8\]\[24\] VGND VGND VPWR VPWR net2509 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1223 CPU.registerFile\[25\]\[13\] VGND VGND VPWR VPWR net2520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1234 CPU.registerFile\[7\]\[15\] VGND VGND VPWR VPWR net2531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1245 CPU.registerFile\[12\]\[10\] VGND VGND VPWR VPWR net2542 sky130_fd_sc_hd__dlygate4sd3_1
X_17348__9 clknet_1_0__leaf__04984_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__inv_2
Xhold1256 CPU.registerFile\[1\]\[25\] VGND VGND VPWR VPWR net2553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 CPU.registerFile\[16\]\[9\] VGND VGND VPWR VPWR net2564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1278 CPU.aluReg\[6\] VGND VGND VPWR VPWR net2575 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1289 mapped_spi_flash.cmd_addr\[30\] VGND VGND VPWR VPWR net2586 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13652__1031 clknet_1_1__leaf__08449_ VGND VGND VPWR VPWR net1087 sky130_fd_sc_hd__inv_2
XFILLER_0_48_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14047__196 clknet_1_1__leaf__08489_ VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__inv_2
X_09318_ _05624_ _05668_ _05558_ VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__a21o_1
X_10590_ net2352 _06292_ _06761_ VGND VGND VPWR VPWR _06762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09249_ CPU.aluIn1\[8\] CPU.Bimm\[8\] VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12260_ net1556 _07799_ _07803_ _07796_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11211_ _07195_ _07196_ net2634 VGND VGND VPWR VPWR _07197_ sky130_fd_sc_hd__mux2_1
X_12191_ net1345 _07738_ _07754_ _07755_ VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput8 net8 VGND VGND VPWR VPWR spi_clk_ram sky130_fd_sc_hd__clkbuf_4
Xoutput10 net10 VGND VGND VPWR VPWR spi_cs_n_ram sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11142_ net1351 _07149_ VGND VGND VPWR VPWR _07153_ sky130_fd_sc_hd__or2_1
X_15635__436 clknet_1_0__leaf__03641_ VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__inv_2
X_11073_ net1545 _07054_ _07105_ _07069_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__o211a_1
X_14901_ _08808_ _08809_ CPU.registerFile\[25\]\[14\] VGND VGND VPWR VPWR _02969_
+ sky130_fd_sc_hd__a21o_1
X_10024_ _06349_ _06351_ _06352_ _05541_ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__o31a_1
X_17620_ _06853_ per_uart.uart0.uart_rxd2 _05168_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__and3_1
X_14832_ CPU.registerFile\[8\]\[12\] _08776_ _02901_ _02864_ VGND VGND VPWR VPWR _02902_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17551_ _05118_ per_uart.uart0.tx_count16\[2\] per_uart.tx_busy VGND VGND VPWR VPWR
+ _05119_ sky130_fd_sc_hd__or3b_1
X_14763_ _08785_ _02830_ _02834_ _08870_ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__a211o_1
X_11975_ _06636_ net2430 _07609_ VGND VGND VPWR VPWR _07619_ sky130_fd_sc_hd__mux2_1
X_16502_ _04170_ _04213_ _04217_ _04180_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17482_ _05060_ _05062_ _05020_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__a21oi_1
X_10926_ _06987_ VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__clkbuf_1
X_14694_ _02765_ _02766_ _08609_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16433_ _04015_ _04147_ _04149_ _03979_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__a211o_1
X_10857_ _06932_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19152_ clknet_leaf_7_clk _02672_ VGND VGND VPWR VPWR per_uart.uart0.tx_bitcount\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16364_ CPU.registerFile\[24\]\[8\] _03915_ _03747_ _04082_ VGND VGND VPWR VPWR _04083_
+ sky130_fd_sc_hd__o211a_1
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10788_ CPU.aluReg\[29\] CPU.aluReg\[27\] _06872_ VGND VGND VPWR VPWR _06879_ sky130_fd_sc_hd__mux2_1
X_13576_ clknet_1_1__leaf__08440_ VGND VGND VPWR VPWR _08443_ sky130_fd_sc_hd__buf_1
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18103_ net1114 _01631_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_15315_ CPU.registerFile\[13\]\[24\] CPU.registerFile\[12\]\[24\] _08794_ VGND VGND
+ VPWR VPWR _03373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12527_ _07951_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19083_ clknet_leaf_0_clk _02603_ VGND VGND VPWR VPWR per_uart.uart0.rxd_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16295_ _03702_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__clkbuf_4
X_18034_ net1045 _01562_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_15246_ CPU.registerFile\[8\]\[22\] _03018_ _03305_ _03268_ VGND VGND VPWR VPWR _03306_
+ sky130_fd_sc_hd__o211a_1
X_12458_ net1724 _07370_ _07906_ VGND VGND VPWR VPWR _07915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11409_ _07302_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__clkbuf_1
X_12389_ _07878_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15177_ _03027_ _03234_ _03238_ _03111_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__a211o_1
XFILLER_0_50_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__03654_ _03654_ VGND VGND VPWR VPWR clknet_0__03654_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_120_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18936_ net710 _02456_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_18867_ net641 _02387_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14152__291 clknet_1_1__leaf__08499_ VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__inv_2
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17818_ net898 _01380_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_18798_ net587 _02322_ VGND VGND VPWR VPWR CPU.aluReg\[28\] sky130_fd_sc_hd__dfxtp_1
X_17749_ net834 _01315_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15740__531 clknet_1_1__leaf__03651_ VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__inv_2
XFILLER_0_17_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09103_ _05428_ _05448_ _05454_ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09034_ _05384_ _05385_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_914 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold320 CPU.aluReg\[0\] VGND VGND VPWR VPWR net1617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold331 CPU.registerFile\[31\]\[17\] VGND VGND VPWR VPWR net1628 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold342 per_uart.uart0.rx_bitcount\[3\] VGND VGND VPWR VPWR net1639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold353 CPU.rs2\[18\] VGND VGND VPWR VPWR net1650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 mapped_spi_flash.snd_bitcount\[1\] VGND VGND VPWR VPWR net1661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 CPU.registerFile\[10\]\[30\] VGND VGND VPWR VPWR net1672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold386 CPU.registerFile\[10\]\[0\] VGND VGND VPWR VPWR net1683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 CPU.registerFile\[15\]\[21\] VGND VGND VPWR VPWR net1694 sky130_fd_sc_hd__dlygate4sd3_1
X_09936_ _06268_ VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__clkbuf_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13791__1155 clknet_1_0__leaf__08464_ VGND VGND VPWR VPWR net1211 sky130_fd_sc_hd__inv_2
X_09867_ _05520_ VGND VGND VPWR VPWR _06202_ sky130_fd_sc_hd__buf_4
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1020 CPU.registerFile\[26\]\[9\] VGND VGND VPWR VPWR net2317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 CPU.registerFile\[16\]\[19\] VGND VGND VPWR VPWR net2328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 CPU.registerFile\[3\]\[3\] VGND VGND VPWR VPWR net2339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1053 CPU.registerFile\[21\]\[25\] VGND VGND VPWR VPWR net2350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1064 CPU.aluIn1\[24\] VGND VGND VPWR VPWR net2361 sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ CPU.PC\[17\] _05890_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__nor2_1
Xhold1075 CPU.registerFile\[23\]\[3\] VGND VGND VPWR VPWR net2372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 CPU.registerFile\[22\]\[18\] VGND VGND VPWR VPWR net2383 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 CPU.registerFile\[21\]\[24\] VGND VGND VPWR VPWR net2394 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03643_ clknet_0__03643_ VGND VGND VPWR VPWR clknet_1_0__leaf__03643_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _07505_ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__clkbuf_1
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _06828_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__clkbuf_1
X_11691_ _07468_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__clkbuf_1
X_18564__21 VGND VGND VPWR VPWR _18564__21/HI net21 sky130_fd_sc_hd__conb_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13614__996 clknet_1_0__leaf__08446_ VGND VGND VPWR VPWR net1052 sky130_fd_sc_hd__inv_2
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10642_ _06790_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__clkbuf_1
X_13430_ _08395_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10573_ net1927 _06106_ _06750_ VGND VGND VPWR VPWR _06753_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15100_ _08419_ VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__clkbuf_4
X_12312_ _07784_ _07834_ _05236_ _07675_ VGND VGND VPWR VPWR _07835_ sky130_fd_sc_hd__a211o_1
XFILLER_0_133_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16080_ CPU.registerFile\[22\]\[1\] CPU.registerFile\[23\]\[1\] _03759_ VGND VGND
+ VPWR VPWR _03806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15031_ CPU.registerFile\[13\]\[17\] CPU.registerFile\[12\]\[17\] _02935_ VGND VGND
+ VPWR VPWR _03096_ sky130_fd_sc_hd__mux2_1
X_12243_ net1373 _07785_ _07793_ _07755_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12174_ net1462 _07738_ _07745_ _07737_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__o211a_1
X_11125_ net1578 _07135_ VGND VGND VPWR VPWR _07143_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16982_ CPU.registerFile\[24\]\[23\] _04319_ _04569_ _04685_ VGND VGND VPWR VPWR
+ _04686_ sky130_fd_sc_hd__o211a_1
X_13872__1229 clknet_1_0__leaf__08471_ VGND VGND VPWR VPWR net1285 sky130_fd_sc_hd__inv_2
X_18721_ net510 _02245_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[21\] sky130_fd_sc_hd__dfxtp_1
X_15933_ clknet_1_0__leaf__03686_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__buf_1
X_11056_ _07048_ _07092_ VGND VGND VPWR VPWR _07093_ sky130_fd_sc_hd__or2_1
X_10007_ net1332 VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__buf_4
X_18652_ clknet_leaf_11_clk _02176_ VGND VGND VPWR VPWR CPU.rs2\[24\] sky130_fd_sc_hd__dfxtp_1
X_17603_ _05237_ _05158_ _05159_ net1451 VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__o22a_1
X_14815_ CPU.registerFile\[20\]\[12\] _08839_ _02884_ _08841_ VGND VGND VPWR VPWR
+ _02885_ sky130_fd_sc_hd__o211a_1
X_18583_ net404 net40 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_15795_ net1582 _08348_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17534_ _08310_ _06039_ _05061_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__or3_1
X_14746_ CPU.registerFile\[15\]\[10\] CPU.registerFile\[14\]\[10\] _08771_ VGND VGND
+ VPWR VPWR _02818_ sky130_fd_sc_hd__mux2_1
X_11958_ _07610_ VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17465_ _05016_ CPU.PC\[8\] _05047_ _05048_ _07002_ VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__o221a_1
X_10909_ net1617 _06971_ _06868_ VGND VGND VPWR VPWR _06972_ sky130_fd_sc_hd__mux2_1
X_14677_ _06339_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__clkbuf_4
X_11889_ _06617_ net1934 _07573_ VGND VGND VPWR VPWR _07574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16416_ _03770_ _03771_ CPU.registerFile\[17\]\[9\] VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13589__973 clknet_1_1__leaf__08444_ VGND VGND VPWR VPWR net1029 sky130_fd_sc_hd__inv_2
XFILLER_0_55_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19135_ clknet_leaf_16_clk _02655_ VGND VGND VPWR VPWR CPU.PC\[17\] sky130_fd_sc_hd__dfxtp_2
X_16347_ _04064_ _04065_ _03720_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19066_ net58 _02586_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[19\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__08492_ clknet_0__08492_ VGND VGND VPWR VPWR clknet_1_1__leaf__08492_
+ sky130_fd_sc_hd__clkbuf_16
X_16278_ _03735_ _03994_ _03998_ _03755_ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__o211a_1
X_18017_ net1028 _01545_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_15229_ CPU.registerFile\[20\]\[22\] _03080_ _03288_ _03082_ VGND VGND VPWR VPWR
+ _03289_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13651__1030 clknet_1_1__leaf__08449_ VGND VGND VPWR VPWR net1086 sky130_fd_sc_hd__inv_2
X_15770__557 clknet_1_1__leaf__03655_ VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__inv_2
X_09721_ _06061_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18919_ net693 _02439_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09652_ CPU.Iimm\[0\] _05545_ _05914_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__mux2_1
X_09583_ CPU.PC\[18\] _05926_ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17306__721 clknet_1_1__leaf__04980_ VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__inv_2
XFILLER_0_9_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09017_ CPU.aluIn1\[21\] _05368_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14159__297 clknet_1_1__leaf__08500_ VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__inv_2
Xhold150 _02221_ VGND VGND VPWR VPWR net1447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold161 mapped_spi_ram.rcv_data\[6\] VGND VGND VPWR VPWR net1458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 mapped_spi_ram.rcv_data\[1\] VGND VGND VPWR VPWR net1469 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold183 mapped_spi_ram.div_counter\[1\] VGND VGND VPWR VPWR net1480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 mapped_spi_flash.cmd_addr\[8\] VGND VGND VPWR VPWR net1491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09919_ _06181_ _06251_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__and2_1
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12930_ _08166_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__clkbuf_1
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _06267_ net2212 _08120_ VGND VGND VPWR VPWR _08130_ sky130_fd_sc_hd__mux2_1
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15747__537 clknet_1_1__leaf__03652_ VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__inv_2
X_14600_ _08526_ VGND VGND VPWR VPWR _08839_ sky130_fd_sc_hd__clkbuf_4
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ net2099 _07324_ _07526_ VGND VGND VPWR VPWR _07533_ sky130_fd_sc_hd__mux2_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ CPU.registerFile\[2\]\[31\] CPU.registerFile\[3\]\[31\] _08564_ VGND VGND
+ VPWR VPWR _03631_ sky130_fd_sc_hd__mux2_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _08092_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__clkbuf_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ CPU.registerFile\[15\]\[5\] CPU.registerFile\[14\]\[5\] _08771_ VGND VGND
+ VPWR VPWR _08772_ sky130_fd_sc_hd__mux2_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _07496_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__clkbuf_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17250_ CPU.registerFile\[8\]\[31\] _03707_ _03708_ _04945_ VGND VGND VPWR VPWR _04946_
+ sky130_fd_sc_hd__o211a_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14462_ CPU.registerFile\[2\]\[3\] CPU.registerFile\[3\]\[3\] _08629_ VGND VGND VPWR
+ VPWR _08705_ sky130_fd_sc_hd__mux2_1
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _07459_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16201_ CPU.registerFile\[19\]\[4\] CPU.registerFile\[18\]\[4\] _03923_ VGND VGND
+ VPWR VPWR _03924_ sky130_fd_sc_hd__mux2_1
X_13413_ _08385_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17181_ CPU.registerFile\[13\]\[29\] _03767_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__or2_1
X_10625_ _06781_ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14393_ CPU.registerFile\[19\]\[2\] CPU.registerFile\[18\]\[2\] _06064_ VGND VGND
+ VPWR VPWR _08637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16132_ CPU.registerFile\[10\]\[3\] CPU.registerFile\[11\]\[3\] _03694_ VGND VGND
+ VPWR VPWR _03856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13344_ clknet_1_0__leaf__08340_ VGND VGND VPWR VPWR _08366_ sky130_fd_sc_hd__buf_1
X_10556_ net2068 _05825_ _06739_ VGND VGND VPWR VPWR _06744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16063_ _03787_ _03788_ _03720_ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10487_ net2015 _05825_ _06702_ VGND VGND VPWR VPWR _06707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13275_ net1624 _08355_ VGND VGND VPWR VPWR _08356_ sky130_fd_sc_hd__or2_1
X_15014_ CPU.registerFile\[22\]\[17\] CPU.registerFile\[23\]\[17\] _02998_ VGND VGND
+ VPWR VPWR _03079_ sky130_fd_sc_hd__mux2_1
X_12226_ mapped_spi_ram.rcv_bitcount\[5\] mapped_spi_ram.rcv_bitcount\[4\] _07781_
+ VGND VGND VPWR VPWR _07782_ sky130_fd_sc_hd__or3_2
X_12157_ mapped_spi_ram.cmd_addr\[12\] _07086_ _07724_ VGND VGND VPWR VPWR _07733_
+ sky130_fd_sc_hd__mux2_1
X_11108_ _07129_ _07131_ VGND VGND VPWR VPWR _07132_ sky130_fd_sc_hd__nand2_4
X_16965_ CPU.registerFile\[13\]\[23\] _04380_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__or2_1
X_12088_ _06856_ _07684_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__nand2_1
X_18704_ net493 _02228_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[4\] sky130_fd_sc_hd__dfxtp_1
X_11039_ CPU.PC\[8\] _05643_ VGND VGND VPWR VPWR _07078_ sky130_fd_sc_hd__or2_1
X_16896_ _04347_ _04599_ _04601_ _04521_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__a211o_1
X_18635_ clknet_leaf_17_clk _02159_ VGND VGND VPWR VPWR CPU.mem_wdata\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_59_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18566_ net387 net23 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17517_ _05069_ net2548 _05090_ _05091_ _05053_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14729_ CPU.registerFile\[16\]\[10\] _02755_ _02800_ _02757_ VGND VGND VPWR VPWR
+ _02801_ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18497_ net318 _02021_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17448_ _06424_ _05024_ _05034_ _05880_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__a211o_1
XFILLER_0_157_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13669__1045 clknet_1_1__leaf__08452_ VGND VGND VPWR VPWR net1101 sky130_fd_sc_hd__inv_2
X_17379_ per_uart.uart0.rxd_reg\[7\] _04992_ _04993_ per_uart.uart0.rxd_reg\[6\] VGND
+ VGND VPWR VPWR _05005_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13790__1154 clknet_1_0__leaf__08464_ VGND VGND VPWR VPWR net1210 sky130_fd_sc_hd__inv_2
X_19118_ net101 _02638_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19049_ net791 _02569_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[2\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__08475_ clknet_0__08475_ VGND VGND VPWR VPWR clknet_1_1__leaf__08475_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09704_ _05380_ _06040_ _06045_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09635_ _05941_ _05977_ _05978_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__a21o_1
X_09566_ _05548_ _05422_ _05538_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__or3b_4
XFILLER_0_66_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15588__393 clknet_1_0__leaf__08511_ VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__inv_2
X_09497_ _05385_ _05522_ _05749_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__o21ai_1
X_13871__1228 clknet_1_0__leaf__08471_ VGND VGND VPWR VPWR net1284 sky130_fd_sc_hd__inv_2
XFILLER_0_19_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10410_ _06593_ net2318 _06665_ VGND VGND VPWR VPWR _06666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11390_ _07292_ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10341_ _06617_ net1694 _06618_ VGND VGND VPWR VPWR _06619_ sky130_fd_sc_hd__mux2_1
X_13060_ net1415 VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__clkbuf_1
X_10272_ net1805 _06200_ _06569_ VGND VGND VPWR VPWR _06576_ sky130_fd_sc_hd__mux2_1
X_14092__237 clknet_1_1__leaf__08493_ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__inv_2
X_12011_ net2320 _07318_ _07635_ VGND VGND VPWR VPWR _07639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16750_ CPU.registerFile\[10\]\[18\] CPU.registerFile\[11\]\[18\] _04335_ VGND VGND
+ VPWR VPWR _04459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12913_ _06083_ net2158 _08156_ VGND VGND VPWR VPWR _08158_ sky130_fd_sc_hd__mux2_1
X_16681_ CPU.registerFile\[0\]\[16\] _04233_ _04068_ _04391_ VGND VGND VPWR VPWR _04392_
+ sky130_fd_sc_hd__o211a_1
X_18420_ net241 _01948_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[20\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__08495_ clknet_0__08495_ VGND VGND VPWR VPWR clknet_1_0__leaf__08495_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _08121_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ net172 _01879_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ CPU.registerFile\[27\]\[31\] CPU.registerFile\[26\]\[31\] _08576_ VGND VGND
+ VPWR VPWR _03614_ sky130_fd_sc_hd__mux2_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _08083_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__clkbuf_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14514_ _08415_ _08752_ _08754_ _08420_ VGND VGND VPWR VPWR _08755_ sky130_fd_sc_hd__a211o_1
X_11726_ _07486_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__clkbuf_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ net1293 _01810_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _03202_ _03534_ _03538_ _03546_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17233_ _03726_ _03727_ CPU.registerFile\[25\]\[30\] VGND VGND VPWR VPWR _04930_
+ sky130_fd_sc_hd__a21o_1
X_14445_ CPU.registerFile\[24\]\[3\] _08686_ _08687_ _08550_ VGND VGND VPWR VPWR _08688_
+ sky130_fd_sc_hd__o211a_1
X_11657_ _07449_ VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17164_ _03714_ _04858_ _04862_ _08403_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__o211a_1
X_10608_ net2296 _06508_ _06761_ VGND VGND VPWR VPWR _06771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14376_ _08567_ _08569_ CPU.registerFile\[9\]\[1\] VGND VGND VPWR VPWR _08621_ sky130_fd_sc_hd__a21o_1
X_11588_ _07412_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16115_ CPU.registerFile\[24\]\[2\] _08393_ _03747_ _03839_ VGND VGND VPWR VPWR _03840_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold908 CPU.registerFile\[21\]\[15\] VGND VGND VPWR VPWR net2205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold919 CPU.registerFile\[26\]\[6\] VGND VGND VPWR VPWR net2216 sky130_fd_sc_hd__dlygate4sd3_1
X_17095_ _04794_ _04795_ _03742_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__mux2_1
X_10539_ net1951 _06508_ _06724_ VGND VGND VPWR VPWR _06734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16046_ CPU.registerFile\[16\]\[0\] _06173_ _03769_ _03772_ VGND VGND VPWR VPWR _03773_
+ sky130_fd_sc_hd__o211a_1
X_12209_ _07769_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13189_ CPU.cycles\[28\] _08303_ net1549 VGND VGND VPWR VPWR _08306_ sky130_fd_sc_hd__a21oi_1
X_17997_ net1008 _01525_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_16948_ CPU.registerFile\[20\]\[22\] CPU.registerFile\[21\]\[22\] _04287_ VGND VGND
+ VPWR VPWR _04653_ sky130_fd_sc_hd__mux2_1
X_13261__781 clknet_1_0__leaf__08344_ VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__inv_2
XFILLER_0_79_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16879_ _04573_ _04585_ _04542_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09420_ _05535_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__buf_4
X_18618_ net439 _02142_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09351_ _05235_ VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__buf_4
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18549_ net370 _02073_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09282_ _05559_ _05560_ _05633_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__08458_ clknet_0__08458_ VGND VGND VPWR VPWR clknet_1_1__leaf__08458_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__08489_ _08489_ VGND VGND VPWR VPWR clknet_0__08489_ sky130_fd_sc_hd__clkbuf_16
X_08997_ CPU.aluIn1\[19\] _05348_ VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__and2_1
X_09618_ CPU.PC\[4\] _05950_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__and2_1
X_10890_ _06957_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__clkbuf_1
X_09549_ CPU.PC\[20\] _05892_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12560_ net2375 _07335_ _07968_ VGND VGND VPWR VPWR _07970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11511_ _06485_ VGND VGND VPWR VPWR _07370_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15859__605 clknet_1_1__leaf__03681_ VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__inv_2
X_12491_ net2111 _07335_ _07931_ VGND VGND VPWR VPWR _07933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11442_ _07323_ VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11373_ _07283_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14100__244 clknet_1_0__leaf__08494_ VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__inv_2
X_13507__900 clknet_1_1__leaf__08435_ VGND VGND VPWR VPWR net956 sky130_fd_sc_hd__inv_2
XFILLER_0_33_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10324_ _05838_ VGND VGND VPWR VPWR _06607_ sky130_fd_sc_hd__clkbuf_4
X_13112_ _06992_ _08262_ VGND VGND VPWR VPWR _08263_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13957__115 clknet_1_0__leaf__08480_ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__inv_2
XFILLER_0_131_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13043_ _08226_ VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__clkbuf_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17920_ clknet_leaf_26_clk _01448_ VGND VGND VPWR VPWR CPU.Bimm\[7\] sky130_fd_sc_hd__dfxtp_2
X_10255_ net1844 _06010_ _06558_ VGND VGND VPWR VPWR _06567_ sky130_fd_sc_hd__mux2_1
X_17851_ net931 _01413_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_10186_ net2297 _06508_ _06293_ VGND VGND VPWR VPWR _06509_ sky130_fd_sc_hd__mux2_1
X_16802_ _04503_ _04504_ _04508_ _04509_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__a211o_1
X_17782_ net862 _01344_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_13668__1044 clknet_1_1__leaf__08452_ VGND VGND VPWR VPWR net1100 sky130_fd_sc_hd__inv_2
X_14994_ _02733_ _02734_ CPU.registerFile\[9\]\[16\] VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__a21o_1
X_16733_ _04080_ _04081_ CPU.registerFile\[25\]\[17\] VGND VGND VPWR VPWR _04443_
+ sky130_fd_sc_hd__a21o_1
X_16664_ CPU.registerFile\[10\]\[16\] CPU.registerFile\[11\]\[16\] _04335_ VGND VGND
+ VPWR VPWR _04375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__08478_ clknet_0__08478_ VGND VGND VPWR VPWR clknet_1_0__leaf__08478_
+ sky130_fd_sc_hd__clkbuf_16
X_18403_ net224 _01931_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_12827_ _08112_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16595_ _04306_ _04307_ _04153_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18334_ net155 _01862_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15546_ _08414_ _03595_ _03597_ _08419_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__a211o_1
X_12758_ _08074_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__clkbuf_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11709_ net2411 _07358_ _07475_ VGND VGND VPWR VPWR _07478_ sky130_fd_sc_hd__mux2_1
X_18265_ net1276 _01793_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15477_ net1584 _03201_ _03530_ _03390_ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__o211a_1
X_12689_ _06613_ net2431 _08029_ VGND VGND VPWR VPWR _08038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17216_ CPU.registerFile\[15\]\[30\] CPU.registerFile\[14\]\[30\] _03698_ VGND VGND
+ VPWR VPWR _04913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14428_ _08663_ _08671_ _08594_ VGND VGND VPWR VPWR _08672_ sky130_fd_sc_hd__o21a_1
XFILLER_0_71_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18196_ net1207 _01724_ VGND VGND VPWR VPWR mapped_spi_ram.snd_bitcount\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17147_ _03766_ _04843_ _04845_ _03716_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__a211o_1
XFILLER_0_80_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold705 CPU.registerFile\[14\]\[7\] VGND VGND VPWR VPWR net2002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14359_ CPU.registerFile\[21\]\[1\] _08528_ VGND VGND VPWR VPWR _08604_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold716 CPU.registerFile\[17\]\[3\] VGND VGND VPWR VPWR net2013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 CPU.registerFile\[21\]\[4\] VGND VGND VPWR VPWR net2024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 CPU.registerFile\[18\]\[28\] VGND VGND VPWR VPWR net2035 sky130_fd_sc_hd__dlygate4sd3_1
X_17078_ _04777_ _04778_ _04557_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__mux2_1
Xhold749 CPU.registerFile\[27\]\[10\] VGND VGND VPWR VPWR net2046 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__08343_ _08343_ VGND VGND VPWR VPWR clknet_0__08343_ sky130_fd_sc_hd__clkbuf_16
X_16029_ _03735_ _03743_ _03754_ _03755_ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__o211a_1
X_08920_ CPU.mem_wdata\[1\] VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13749__1118 clknet_1_1__leaf__08459_ VGND VGND VPWR VPWR net1174 sky130_fd_sc_hd__inv_2
X_13870__1227 clknet_1_0__leaf__08471_ VGND VGND VPWR VPWR net1283 sky130_fd_sc_hd__inv_2
X_15964__700 clknet_1_0__leaf__03691_ VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__inv_2
XFILLER_0_79_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09403_ _05415_ _05753_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__and2b_1
XFILLER_0_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09334_ mapped_spi_ram.rcv_data\[7\] _05685_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09265_ _05567_ _05569_ _05594_ _05605_ _05616_ VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__a311o_1
XFILLER_0_16_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09196_ _05547_ CPU.instr\[6\] CPU.instr\[2\] VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__or3b_1
XFILLER_0_161_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10040_ _05547_ _05880_ VGND VGND VPWR VPWR _06368_ sky130_fd_sc_hd__or2_2
Xhold10 mapped_spi_ram.state\[2\] VGND VGND VPWR VPWR net1307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 mapped_spi_ram.cmd_addr\[0\] VGND VGND VPWR VPWR net1318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 _08231_ VGND VGND VPWR VPWR net1329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 _08222_ VGND VGND VPWR VPWR net1340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 mapped_spi_flash.rcv_data\[18\] VGND VGND VPWR VPWR net1351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 _06529_ VGND VGND VPWR VPWR net1362 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold76 mapped_spi_ram.rcv_data\[25\] VGND VGND VPWR VPWR net1373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 mapped_spi_flash.rcv_data\[16\] VGND VGND VPWR VPWR net1384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 _07187_ VGND VGND VPWR VPWR net1395 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ _07627_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10942_ _06998_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10873_ net1331 _06944_ _06922_ VGND VGND VPWR VPWR _06945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15400_ CPU.registerFile\[0\]\[26\] _08411_ _03455_ _03195_ VGND VGND VPWR VPWR _03456_
+ sky130_fd_sc_hd__o211a_1
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12612_ _07997_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__clkbuf_1
X_16380_ _08403_ VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_149_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15331_ _03155_ _03371_ _03388_ _03243_ VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__a211o_2
XFILLER_0_137_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12543_ net2549 _07318_ _07957_ VGND VGND VPWR VPWR _07961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18050_ net1061 _01578_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_15262_ CPU.registerFile\[17\]\[23\] _03036_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__or2_1
X_12474_ net1869 _07318_ _07920_ VGND VGND VPWR VPWR _07924_ sky130_fd_sc_hd__mux2_1
X_14024__175 clknet_1_0__leaf__08487_ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__inv_2
X_17001_ CPU.registerFile\[13\]\[24\] _04380_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__or2_1
X_11425_ _07311_ VGND VGND VPWR VPWR _07312_ sky130_fd_sc_hd__buf_4
XFILLER_0_50_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15193_ CPU.registerFile\[28\]\[21\] CPU.registerFile\[29\]\[21\] _03212_ VGND VGND
+ VPWR VPWR _03254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13583__968 clknet_1_1__leaf__08443_ VGND VGND VPWR VPWR net1024 sky130_fd_sc_hd__inv_2
XANTENNA_7 _02838_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11356_ net1851 _05734_ _07274_ VGND VGND VPWR VPWR _07275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10307_ _05735_ _05736_ CPU.writeBack VGND VGND VPWR VPWR _06595_ sky130_fd_sc_hd__and3_4
X_18952_ net726 _02472_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_14075_ clknet_1_0__leaf__08484_ VGND VGND VPWR VPWR _08492_ sky130_fd_sc_hd__buf_1
X_11287_ _07237_ VGND VGND VPWR VPWR _07238_ sky130_fd_sc_hd__buf_4
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ CPU.registerFile\[4\]\[31\] net1410 _08217_ VGND VGND VPWR VPWR _08218_ sky130_fd_sc_hd__mux2_1
X_17903_ clknet_leaf_25_clk _01431_ VGND VGND VPWR VPWR CPU.Bimm\[3\] sky130_fd_sc_hd__dfxtp_1
X_10238_ _06557_ VGND VGND VPWR VPWR _06558_ sky130_fd_sc_hd__buf_4
X_18883_ net657 _02403_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_10169_ mapped_spi_ram.rcv_data\[26\] _05857_ VGND VGND VPWR VPWR _06492_ sky130_fd_sc_hd__and2_1
X_17834_ net914 _01396_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15612__415 clknet_1_1__leaf__03639_ VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__inv_2
XFILLER_0_107_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17765_ net845 _01327_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_14977_ _08532_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__buf_4
X_16716_ _06171_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__buf_4
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17696_ _05207_ _05221_ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16647_ CPU.registerFile\[24\]\[15\] _04319_ _04165_ _04358_ VGND VGND VPWR VPWR
+ _04359_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16578_ CPU.registerFile\[16\]\[13\] _04252_ _04090_ _04291_ VGND VGND VPWR VPWR
+ _04292_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15529_ _08580_ _03578_ _03580_ _08418_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__a211o_1
X_18317_ net138 _01845_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09050_ _05381_ _05382_ _05401_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__a21o_1
X_18248_ net1259 _01776_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18179_ net1190 _01707_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold502 CPU.registerFile\[7\]\[24\] VGND VGND VPWR VPWR net1799 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold513 CPU.registerFile\[20\]\[26\] VGND VGND VPWR VPWR net1810 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold524 CPU.registerFile\[28\]\[14\] VGND VGND VPWR VPWR net1821 sky130_fd_sc_hd__dlygate4sd3_1
Xhold535 CPU.registerFile\[27\]\[29\] VGND VGND VPWR VPWR net1832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 CPU.registerFile\[13\]\[31\] VGND VGND VPWR VPWR net1843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 CPU.registerFile\[22\]\[15\] VGND VGND VPWR VPWR net1854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold568 CPU.registerFile\[30\]\[26\] VGND VGND VPWR VPWR net1865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold579 CPU.registerFile\[20\]\[23\] VGND VGND VPWR VPWR net1876 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ _05887_ _06283_ VGND VGND VPWR VPWR _06284_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08903_ CPU.aluIn1\[29\] _05254_ VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__and2_2
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _05939_ _05979_ _05984_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__a21bo_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1202 CPU.registerFile\[1\]\[20\] VGND VGND VPWR VPWR net2499 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1213 CPU.registerFile\[23\]\[28\] VGND VGND VPWR VPWR net2510 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 CPU.registerFile\[1\]\[30\] VGND VGND VPWR VPWR net2521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 CPU.registerFile\[18\]\[22\] VGND VGND VPWR VPWR net2532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 CPU.registerFile\[25\]\[20\] VGND VGND VPWR VPWR net2543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 CPU.registerFile\[30\]\[2\] VGND VGND VPWR VPWR net2554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1268 CPU.registerFile\[1\]\[14\] VGND VGND VPWR VPWR net2565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 CPU.registerFile\[8\]\[6\] VGND VGND VPWR VPWR net2576 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09317_ _05624_ _05668_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09248_ _05595_ _05596_ _05599_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13667__1043 clknet_1_1__leaf__08452_ VGND VGND VPWR VPWR net1099 sky130_fd_sc_hd__inv_2
XFILLER_0_16_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09179_ _05530_ _05527_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__nor2_2
XFILLER_0_133_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11210_ mapped_spi_flash.rcv_bitcount\[0\] mapped_spi_flash.state\[3\] _07188_ VGND
+ VGND VPWR VPWR _07196_ sky130_fd_sc_hd__a21o_1
X_12190_ _07163_ VGND VGND VPWR VPWR _07755_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput11 net11 VGND VGND VPWR VPWR spi_mosi sky130_fd_sc_hd__clkbuf_4
Xoutput9 net9 VGND VGND VPWR VPWR spi_cs_n sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11141_ net1351 _07147_ _07152_ _07151_ VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11072_ _06983_ _07104_ VGND VGND VPWR VPWR _07105_ sky130_fd_sc_hd__or2_1
X_14900_ CPU.registerFile\[27\]\[14\] CPU.registerFile\[26\]\[14\] _02768_ VGND VGND
+ VPWR VPWR _02968_ sky130_fd_sc_hd__mux2_1
X_10023_ _05267_ _05523_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__nor2_1
X_13281__784 clknet_1_1__leaf__08345_ VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__inv_2
X_14212__345 clknet_1_0__leaf__08505_ VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__inv_2
X_14831_ _02733_ _02734_ CPU.registerFile\[9\]\[12\] VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17550_ per_uart.uart0.tx_count16\[1\] per_uart.uart0.tx_count16\[0\] VGND VGND VPWR
+ VPWR _05118_ sky130_fd_sc_hd__or2_1
X_14762_ CPU.registerFile\[0\]\[10\] _08706_ _02833_ _02791_ VGND VGND VPWR VPWR _02834_
+ sky130_fd_sc_hd__o211a_1
X_13891__55 clknet_1_0__leaf__08474_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__inv_2
X_11974_ _07618_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__clkbuf_1
X_16501_ _03963_ _04214_ _04216_ _04006_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__a211o_1
X_17481_ _05055_ _06284_ _05061_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__or3_1
X_10925_ _06973_ _06986_ VGND VGND VPWR VPWR _06987_ sky130_fd_sc_hd__and2_1
X_14693_ CPU.registerFile\[28\]\[9\] CPU.registerFile\[29\]\[9\] _08538_ VGND VGND
+ VPWR VPWR _02766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16432_ CPU.registerFile\[12\]\[10\] _04017_ _04018_ _04148_ VGND VGND VPWR VPWR
+ _04149_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10856_ net2672 _06931_ _06922_ VGND VGND VPWR VPWR _06932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19151_ clknet_leaf_4_clk _02671_ VGND VGND VPWR VPWR per_uart.uart0.tx_bitcount\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16363_ _04080_ _04081_ CPU.registerFile\[25\]\[8\] VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__a21o_1
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14106__250 clknet_1_1__leaf__08494_ VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__inv_2
X_10787_ _06878_ VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__clkbuf_1
X_18102_ net1113 _01630_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_13748__1117 clknet_1_1__leaf__08459_ VGND VGND VPWR VPWR net1173 sky130_fd_sc_hd__inv_2
XFILLER_0_82_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15314_ CPU.registerFile\[15\]\[24\] CPU.registerFile\[14\]\[24\] _03013_ VGND VGND
+ VPWR VPWR _03372_ sky130_fd_sc_hd__mux2_1
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12526_ net2162 _07370_ _07942_ VGND VGND VPWR VPWR _07951_ sky130_fd_sc_hd__mux2_1
X_19082_ clknet_leaf_27_clk _02602_ VGND VGND VPWR VPWR per_uart.uart0.rxd_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16294_ _08398_ _04011_ _04013_ _08401_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__a211o_1
XFILLER_0_82_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18033_ net1044 _01561_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_15245_ _03138_ _03139_ CPU.registerFile\[9\]\[22\] VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__a21o_1
X_12457_ _07914_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11408_ net2071 _06413_ _07296_ VGND VGND VPWR VPWR _07302_ sky130_fd_sc_hd__mux2_1
X_15176_ CPU.registerFile\[0\]\[20\] _02948_ _03237_ _03195_ VGND VGND VPWR VPWR _03238_
+ sky130_fd_sc_hd__o211a_1
X_12388_ _06653_ net1827 _07870_ VGND VGND VPWR VPWR _07878_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__03653_ _03653_ VGND VGND VPWR VPWR clknet_0__03653_ sky130_fd_sc_hd__clkbuf_16
X_15837__585 clknet_1_1__leaf__03679_ VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__inv_2
X_11339_ _07265_ VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__clkbuf_1
X_13364__859 clknet_1_1__leaf__08368_ VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__inv_2
XFILLER_0_120_672 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18935_ net709 _02455_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_13009_ _08208_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18866_ net640 _02386_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_14187__322 clknet_1_1__leaf__08503_ VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__inv_2
X_17817_ net897 _01379_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_18797_ net586 _02321_ VGND VGND VPWR VPWR CPU.aluReg\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17748_ net833 _01314_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_17679_ _05680_ _05659_ _05208_ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09102_ _05310_ _05449_ _05451_ _05453_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__or4b_1
XFILLER_0_150_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17391__15 clknet_1_1__leaf__04985_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__inv_2
XFILLER_0_150_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09033_ CPU.aluIn1\[25\] _05383_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__and2_2
X_13566__952 clknet_1_0__leaf__08442_ VGND VGND VPWR VPWR net1008 sky130_fd_sc_hd__inv_2
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_926 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold310 _08302_ VGND VGND VPWR VPWR net1607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 _08179_ VGND VGND VPWR VPWR net1618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 CPU.cycles\[19\] VGND VGND VPWR VPWR net1629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold343 mapped_spi_flash.rcv_data\[1\] VGND VGND VPWR VPWR net1640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold354 CPU.rs2\[8\] VGND VGND VPWR VPWR net1651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 per_uart.uart0.rxd_reg\[4\] VGND VGND VPWR VPWR net1662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 CPU.registerFile\[3\]\[19\] VGND VGND VPWR VPWR net1673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 CPU.registerFile\[19\]\[21\] VGND VGND VPWR VPWR net1684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 CPU.registerFile\[19\]\[29\] VGND VGND VPWR VPWR net1695 sky130_fd_sc_hd__dlygate4sd3_1
X_09935_ net2290 _06267_ _06055_ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ _06201_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__clkbuf_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1010 CPU.registerFile\[8\]\[26\] VGND VGND VPWR VPWR net2307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 CPU.registerFile\[14\]\[31\] VGND VGND VPWR VPWR net2318 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 CPU.registerFile\[21\]\[21\] VGND VGND VPWR VPWR net2329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 CPU.registerFile\[20\]\[16\] VGND VGND VPWR VPWR net2340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1054 CPU.registerFile\[22\]\[23\] VGND VGND VPWR VPWR net2351 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ _05933_ _05993_ VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__xnor2_1
Xhold1065 CPU.registerFile\[12\]\[26\] VGND VGND VPWR VPWR net2362 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1076 CPU.registerFile\[14\]\[29\] VGND VGND VPWR VPWR net2373 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 CPU.registerFile\[1\]\[27\] VGND VGND VPWR VPWR net2384 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1098 CPU.registerFile\[7\]\[3\] VGND VGND VPWR VPWR net2395 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03642_ clknet_0__03642_ VGND VGND VPWR VPWR clknet_1_0__leaf__03642_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ net2176 _06054_ _06827_ VGND VGND VPWR VPWR _06828_ sky130_fd_sc_hd__mux2_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ net2439 _07339_ _07464_ VGND VGND VPWR VPWR _07468_ sky130_fd_sc_hd__mux2_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15942__680 clknet_1_0__leaf__03689_ VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__inv_2
XFILLER_0_64_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10641_ net2499 _06083_ _06788_ VGND VGND VPWR VPWR _06790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10572_ _06752_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12311_ net1298 net1302 VGND VGND VPWR VPWR _07834_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13928__89 clknet_1_1__leaf__08477_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__inv_2
XFILLER_0_106_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15030_ CPU.registerFile\[15\]\[17\] CPU.registerFile\[14\]\[17\] _03013_ VGND VGND
+ VPWR VPWR _03095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_948 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12242_ mapped_spi_ram.rcv_data\[26\] _07787_ VGND VGND VPWR VPWR _07793_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12173_ _07739_ _07744_ VGND VGND VPWR VPWR _07745_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11124_ net1578 _07133_ _07142_ _07138_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__o211a_1
X_14136__276 clknet_1_0__leaf__08498_ VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__inv_2
X_16981_ _04484_ _04485_ CPU.registerFile\[25\]\[23\] VGND VGND VPWR VPWR _04685_
+ sky130_fd_sc_hd__a21o_1
X_18720_ net509 _02244_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[20\] sky130_fd_sc_hd__dfxtp_1
X_11055_ mapped_spi_flash.cmd_addr\[5\] _07091_ _07039_ VGND VGND VPWR VPWR _07092_
+ sky130_fd_sc_hd__mux2_1
X_10006_ _05745_ _06326_ _06331_ _06335_ VGND VGND VPWR VPWR _06336_ sky130_fd_sc_hd__a211o_1
X_18651_ clknet_leaf_11_clk _02175_ VGND VGND VPWR VPWR CPU.rs2\[23\] sky130_fd_sc_hd__dfxtp_1
X_14814_ CPU.registerFile\[21\]\[12\] _08718_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__or2_1
X_17602_ _05134_ _05157_ _05236_ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__a21oi_4
X_15794_ _03665_ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__clkbuf_1
X_18582_ net403 net39 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_17533_ _05075_ _05025_ _06051_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__o21bai_1
X_14745_ _02798_ _02802_ _02806_ _02816_ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__a31o_1
X_11957_ _06617_ net2348 _07609_ VGND VGND VPWR VPWR _07610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17464_ _05022_ _06347_ _08256_ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10908_ CPU.aluReg\[1\] _06861_ _06862_ _06970_ VGND VGND VPWR VPWR _06971_ sky130_fd_sc_hd__a31o_1
X_14676_ net1651 _08514_ _02749_ _08751_ VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__o211a_1
X_11888_ _07561_ VGND VGND VPWR VPWR _07573_ sky130_fd_sc_hd__buf_4
X_15724__516 clknet_1_0__leaf__03650_ VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__inv_2
XFILLER_0_39_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16415_ CPU.registerFile\[19\]\[9\] CPU.registerFile\[18\]\[9\] _03923_ VGND VGND
+ VPWR VPWR _04133_ sky130_fd_sc_hd__mux2_1
X_10839_ net2668 _06918_ _06889_ VGND VGND VPWR VPWR _06919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16346_ CPU.registerFile\[5\]\[8\] CPU.registerFile\[4\]\[8\] _04024_ VGND VGND VPWR
+ VPWR _04065_ sky130_fd_sc_hd__mux2_1
X_19134_ clknet_leaf_16_clk _02654_ VGND VGND VPWR VPWR CPU.PC\[16\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_82_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12509_ _07919_ VGND VGND VPWR VPWR _07942_ sky130_fd_sc_hd__buf_4
XFILLER_0_120_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19065_ net807 _02585_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_16277_ _03702_ _03995_ _03997_ _03803_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__a211o_1
XFILLER_0_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__08491_ clknet_0__08491_ VGND VGND VPWR VPWR clknet_1_1__leaf__08491_
+ sky130_fd_sc_hd__clkbuf_16
X_18016_ net1027 _01544_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_15228_ CPU.registerFile\[21\]\[22\] _02960_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15159_ _03202_ _03206_ _03210_ _03220_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__a31o_1
X_15618__421 clknet_1_0__leaf__03639_ VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__inv_2
X_09720_ _06060_ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__buf_4
X_18918_ net692 _02438_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_09651_ _05929_ _05994_ _05927_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__a21o_1
X_18849_ clknet_leaf_7_clk _02373_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_13666__1042 clknet_1_1__leaf__08452_ VGND VGND VPWR VPWR net1098 sky130_fd_sc_hd__inv_2
X_09582_ CPU.Jimm\[18\] _05921_ _05923_ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14241__371 clknet_1_0__leaf__08508_ VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__inv_2
XFILLER_0_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09016_ CPU.rs2\[21\] _05246_ _05250_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__o21a_1
X_13347__843 clknet_1_1__leaf__08367_ VGND VGND VPWR VPWR net899 sky130_fd_sc_hd__inv_2
Xhold140 mapped_spi_ram.rcv_data\[29\] VGND VGND VPWR VPWR net1437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 CPU.cycles\[0\] VGND VGND VPWR VPWR net1448 sky130_fd_sc_hd__buf_1
Xhold162 mapped_spi_ram.rcv_data\[5\] VGND VGND VPWR VPWR net1459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold173 _01691_ VGND VGND VPWR VPWR net1470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _02712_ VGND VGND VPWR VPWR net1481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold195 mapped_spi_flash.cmd_addr\[3\] VGND VGND VPWR VPWR net1492 sky130_fd_sc_hd__dlygate4sd3_1
X_09918_ _05319_ _06180_ _05455_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__or3_1
X_13747__1116 clknet_1_1__leaf__08459_ VGND VGND VPWR VPWR net1172 sky130_fd_sc_hd__inv_2
X_09849_ _05470_ _06184_ _05328_ VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__a21oi_1
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ _08129_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__clkbuf_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _07532_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__clkbuf_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _06647_ net2357 _08087_ VGND VGND VPWR VPWR _08092_ sky130_fd_sc_hd__mux2_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _06061_ VGND VGND VPWR VPWR _08771_ sky130_fd_sc_hd__buf_4
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _06607_ net2052 _07490_ VGND VGND VPWR VPWR _07496_ sky130_fd_sc_hd__mux2_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _08702_ _08703_ _08578_ VGND VGND VPWR VPWR _08704_ sky130_fd_sc_hd__mux2_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11673_ net2307 _07322_ _07453_ VGND VGND VPWR VPWR _07459_ sky130_fd_sc_hd__mux2_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16200_ _03744_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__buf_4
X_13412_ _05735_ _06341_ _00000_ VGND VGND VPWR VPWR _08385_ sky130_fd_sc_hd__mux2_1
X_17180_ CPU.registerFile\[15\]\[29\] CPU.registerFile\[14\]\[29\] _04550_ VGND VGND
+ VPWR VPWR _04878_ sky130_fd_sc_hd__mux2_1
X_10624_ net2557 _05805_ _06777_ VGND VGND VPWR VPWR _06781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14392_ CPU.mem_wdata\[1\] _08514_ _08636_ _07822_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16131_ CPU.aluIn1\[2\] _03566_ _03854_ _03855_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__o211a_1
X_10555_ _06743_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16062_ CPU.registerFile\[5\]\[1\] CPU.registerFile\[4\]\[1\] _03704_ VGND VGND VPWR
+ VPWR _03788_ sky130_fd_sc_hd__mux2_1
X_13274_ net1587 _08354_ VGND VGND VPWR VPWR _08355_ sky130_fd_sc_hd__or2_1
X_10486_ _06706_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15013_ _08520_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__clkbuf_4
X_12225_ mapped_spi_ram.rcv_bitcount\[3\] _07780_ VGND VGND VPWR VPWR _07781_ sky130_fd_sc_hd__or2_2
X_13287__790 clknet_1_0__leaf__08345_ VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__inv_2
X_14218__351 clknet_1_1__leaf__08505_ VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__inv_2
X_12156_ net1519 _07714_ _07732_ _07713_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__o211a_1
X_11107_ _06974_ _07130_ VGND VGND VPWR VPWR _07131_ sky130_fd_sc_hd__nor2_1
X_16964_ CPU.registerFile\[15\]\[23\] CPU.registerFile\[14\]\[23\] _04550_ VGND VGND
+ VPWR VPWR _04668_ sky130_fd_sc_hd__mux2_1
X_12087_ _07670_ _07674_ _07677_ _07683_ VGND VGND VPWR VPWR _07684_ sky130_fd_sc_hd__a22o_1
X_18703_ net492 _02227_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[3\] sky130_fd_sc_hd__dfxtp_1
X_11038_ _07055_ _07076_ VGND VGND VPWR VPWR _07077_ sky130_fd_sc_hd__nor2_1
X_16895_ CPU.registerFile\[0\]\[21\] _04233_ _04472_ _04600_ VGND VGND VPWR VPWR _04601_
+ sky130_fd_sc_hd__o211a_1
X_18634_ clknet_leaf_17_clk _02158_ VGND VGND VPWR VPWR CPU.mem_wdata\[6\] sky130_fd_sc_hd__dfxtp_2
X_15949__686 clknet_1_1__leaf__03690_ VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__inv_2
XFILLER_0_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18565_ net386 net22 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_12989_ net2131 _07343_ _08192_ VGND VGND VPWR VPWR _08198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17516_ _08335_ _06128_ _05073_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14728_ CPU.registerFile\[17\]\[10\] _08795_ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__or2_1
X_18496_ net317 _02020_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14659_ _06058_ VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__clkbuf_4
X_17447_ _08311_ _06422_ _08331_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__nor3_1
XFILLER_0_157_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17378_ _05004_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19117_ net100 _02637_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_16329_ CPU.registerFile\[16\]\[7\] _03848_ _03769_ _04048_ VGND VGND VPWR VPWR _04049_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19048_ net790 _02568_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[1\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__08474_ clknet_0__08474_ VGND VGND VPWR VPWR clknet_1_1__leaf__08474_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17336__748 clknet_1_1__leaf__04983_ VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__inv_2
X_15694__489 clknet_1_1__leaf__03647_ VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__inv_2
XFILLER_0_11_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09703_ _06017_ _06042_ _06044_ _05800_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09634_ _05923_ _05940_ CPU.PC\[12\] VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__o21a_1
X_09565_ CPU.Iimm\[3\] _05758_ _05790_ CPU.cycles\[23\] _05908_ VGND VGND VPWR VPWR
+ _05909_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09496_ _05555_ _05841_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10340_ _06596_ VGND VGND VPWR VPWR _06618_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10271_ _06575_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__clkbuf_1
X_12010_ _07638_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__clkbuf_1
X_15753__542 clknet_1_0__leaf__03653_ VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__inv_2
X_12912_ _08157_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__clkbuf_1
X_16680_ _04389_ _04390_ CPU.registerFile\[1\]\[16\] VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__a21o_1
Xclkbuf_1_0__f__08494_ clknet_0__08494_ VGND VGND VPWR VPWR clknet_1_0__leaf__08494_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12843_ _06054_ net2379 _08120_ VGND VGND VPWR VPWR _08121_ sky130_fd_sc_hd__mux2_1
X_14248__377 clknet_1_0__leaf__08509_ VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__inv_2
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18350_ net171 _01878_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_15562_ _03611_ _03612_ _08588_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__mux2_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _06630_ net2517 _08076_ VGND VGND VPWR VPWR _08083_ sky130_fd_sc_hd__mux2_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ CPU.registerFile\[16\]\[5\] _08412_ _08753_ _06037_ VGND VGND VPWR VPWR _08754_
+ sky130_fd_sc_hd__o211a_1
X_11725_ net2273 _07374_ _07452_ VGND VGND VPWR VPWR _07486_ sky130_fd_sc_hd__mux2_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15493_ _06013_ _03541_ _03545_ _08422_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__o211a_1
X_18281_ net1292 _01809_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17232_ CPU.registerFile\[27\]\[30\] CPU.registerFile\[26\]\[30\] _04646_ VGND VGND
+ VPWR VPWR _04929_ sky130_fd_sc_hd__mux2_1
X_14444_ _08546_ _08547_ CPU.registerFile\[25\]\[3\] VGND VGND VPWR VPWR _08687_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11656_ net2100 _07374_ _07415_ VGND VGND VPWR VPWR _07449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17163_ _03722_ _04859_ _04861_ _04612_ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__a211o_1
X_10607_ _06770_ VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14375_ CPU.registerFile\[10\]\[1\] CPU.registerFile\[11\]\[1\] _08564_ VGND VGND
+ VPWR VPWR _08620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_870 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11587_ net1836 _07374_ _07378_ VGND VGND VPWR VPWR _07412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16114_ _03749_ _03751_ CPU.registerFile\[25\]\[2\] VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17094_ CPU.registerFile\[20\]\[26\] CPU.registerFile\[21\]\[26\] _03737_ VGND VGND
+ VPWR VPWR _04795_ sky130_fd_sc_hd__mux2_1
Xhold909 CPU.registerFile\[29\]\[24\] VGND VGND VPWR VPWR net2206 sky130_fd_sc_hd__dlygate4sd3_1
X_10538_ _06733_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16045_ _03770_ _03771_ CPU.registerFile\[17\]\[0\] VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10469_ _06696_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__clkbuf_1
X_12208_ _07768_ net1330 _07764_ VGND VGND VPWR VPWR _07769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13188_ CPU.cycles\[28\] CPU.cycles\[29\] _08303_ VGND VGND VPWR VPWR _08305_ sky130_fd_sc_hd__and3_1
X_12139_ _07715_ _07720_ VGND VGND VPWR VPWR _07721_ sky130_fd_sc_hd__or2_1
X_17996_ net1007 _01524_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16947_ CPU.registerFile\[22\]\[22\] CPU.registerFile\[23\]\[22\] _04362_ VGND VGND
+ VPWR VPWR _04652_ sky130_fd_sc_hd__mux2_1
X_16878_ _04574_ _04577_ _04583_ _04584_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__o211a_1
X_18617_ net438 _02141_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_15882__626 clknet_1_1__leaf__03683_ VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__inv_2
XFILLER_0_149_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09350_ CPU.PC\[3\] _05643_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__or2_1
X_18548_ net369 _02072_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13530__921 clknet_1_0__leaf__08437_ VGND VGND VPWR VPWR net977 sky130_fd_sc_hd__inv_2
X_09281_ _05629_ _05632_ _05630_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__a21oi_1
X_18479_ net300 _02003_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13980__136 clknet_1_1__leaf__08482_ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__inv_2
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13746__1115 clknet_1_0__leaf__08459_ VGND VGND VPWR VPWR net1171 sky130_fd_sc_hd__inv_2
XFILLER_0_132_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15702__496 clknet_1_0__leaf__03648_ VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__08457_ clknet_0__08457_ VGND VGND VPWR VPWR clknet_1_1__leaf__08457_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08488_ _08488_ VGND VGND VPWR VPWR clknet_0__08488_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08996_ CPU.rs2\[19\] _05246_ _05250_ VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__o21a_1
X_09617_ _05957_ _05959_ _05960_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09548_ CPU.PC\[19\] CPU.PC\[18\] _05891_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09479_ _05826_ VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11510_ _07369_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12490_ _07932_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11441_ net1800 _07322_ _07312_ VGND VGND VPWR VPWR _07323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11372_ net1706 _06010_ _07274_ VGND VGND VPWR VPWR _07283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13111_ _07670_ _07674_ _07761_ _07749_ VGND VGND VPWR VPWR _08262_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10323_ _06606_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__clkbuf_1
X_17319__732 clknet_1_0__leaf__04982_ VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__inv_2
X_15677__473 clknet_1_0__leaf__03646_ VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__inv_2
X_13042_ net2179 _06009_ _08217_ VGND VGND VPWR VPWR _08226_ sky130_fd_sc_hd__mux2_1
X_10254_ _06566_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__clkbuf_1
X_17850_ net930 _01412_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_13245__766 clknet_1_0__leaf__08343_ VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__inv_2
X_10185_ _06507_ VGND VGND VPWR VPWR _06508_ sky130_fd_sc_hd__clkbuf_4
X_16801_ _08400_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__clkbuf_4
X_17781_ net861 _01343_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_14993_ CPU.registerFile\[10\]\[16\] CPU.registerFile\[11\]\[16\] _02779_ VGND VGND
+ VPWR VPWR _03059_ sky130_fd_sc_hd__mux2_1
X_16732_ CPU.registerFile\[27\]\[17\] CPU.registerFile\[26\]\[17\] _04242_ VGND VGND
+ VPWR VPWR _04442_ sky130_fd_sc_hd__mux2_1
X_13875_ clknet_1_1__leaf__08462_ VGND VGND VPWR VPWR _08472_ sky130_fd_sc_hd__buf_1
X_16663_ CPU.aluIn1\[15\] _04054_ _04374_ _04259_ VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__08477_ clknet_0__08477_ VGND VGND VPWR VPWR clknet_1_0__leaf__08477_
+ sky130_fd_sc_hd__clkbuf_16
X_18402_ net223 _01930_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_12826_ _05786_ net2284 _08109_ VGND VGND VPWR VPWR _08112_ sky130_fd_sc_hd__mux2_1
X_14181__317 clknet_1_1__leaf__08502_ VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__inv_2
X_16594_ CPU.registerFile\[5\]\[14\] CPU.registerFile\[4\]\[14\] _04024_ VGND VGND
+ VPWR VPWR _04307_ sky130_fd_sc_hd__mux2_1
X_13806__1169 clknet_1_0__leaf__08465_ VGND VGND VPWR VPWR net1225 sky130_fd_sc_hd__inv_2
XFILLER_0_158_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18333_ net154 _01861_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15545_ CPU.registerFile\[0\]\[30\] _08411_ _03596_ _06036_ VGND VGND VPWR VPWR _03597_
+ sky130_fd_sc_hd__o211a_1
X_12757_ _06613_ net2266 _08065_ VGND VGND VPWR VPWR _08074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _07477_ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18264_ net1275 _01792_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_15476_ _03155_ _03512_ _03529_ _03243_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__a211o_2
X_12688_ _08037_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17215_ _03703_ _04909_ _04911_ _06142_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__a211o_1
X_14427_ _08574_ _08666_ _08670_ _08592_ VGND VGND VPWR VPWR _08671_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11639_ _07440_ VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__clkbuf_1
X_18195_ net1206 net1313 VGND VGND VPWR VPWR mapped_spi_ram.snd_bitcount\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17146_ CPU.registerFile\[12\]\[28\] _03694_ _03763_ _04844_ VGND VGND VPWR VPWR
+ _04845_ sky130_fd_sc_hd__o211a_1
X_14358_ CPU.registerFile\[22\]\[1\] CPU.registerFile\[23\]\[1\] _08523_ VGND VGND
+ VPWR VPWR _08603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold706 CPU.registerFile\[18\]\[23\] VGND VGND VPWR VPWR net2003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 CPU.registerFile\[2\]\[31\] VGND VGND VPWR VPWR net2014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold728 CPU.registerFile\[15\]\[31\] VGND VGND VPWR VPWR net2025 sky130_fd_sc_hd__dlygate4sd3_1
X_17077_ CPU.registerFile\[5\]\[26\] CPU.registerFile\[4\]\[26\] _04428_ VGND VGND
+ VPWR VPWR _04778_ sky130_fd_sc_hd__mux2_1
X_14001__154 clknet_1_1__leaf__08485_ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__inv_2
XFILLER_0_0_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold739 CPU.registerFile\[27\]\[31\] VGND VGND VPWR VPWR net2036 sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ _08532_ VGND VGND VPWR VPWR _08535_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__08342_ _08342_ VGND VGND VPWR VPWR clknet_0__08342_ sky130_fd_sc_hd__clkbuf_16
X_13560__947 clknet_1_1__leaf__08441_ VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__inv_2
X_16028_ _08403_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__buf_4
XFILLER_0_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13897__61 clknet_1_1__leaf__08474_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__inv_2
XFILLER_0_137_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17979_ net990 _01507_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09402_ _05414_ _05255_ _05259_ _05411_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__or4_1
XFILLER_0_149_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09333_ _05683_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09264_ _05608_ _05610_ _05612_ _05615_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__or4_1
XFILLER_0_118_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09195_ CPU.instr\[3\] VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__buf_2
XFILLER_0_117_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__08509_ clknet_0__08509_ VGND VGND VPWR VPWR clknet_1_1__leaf__08509_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13728__1099 clknet_1_1__leaf__08457_ VGND VGND VPWR VPWR net1155 sky130_fd_sc_hd__inv_2
XFILLER_0_12_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold11 _07760_ VGND VGND VPWR VPWR net1308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 mapped_spi_ram.rcv_data\[0\] VGND VGND VPWR VPWR net1319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 mapped_spi_ram.snd_bitcount\[4\] VGND VGND VPWR VPWR net1330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 mapped_spi_ram.cmd_addr\[7\] VGND VGND VPWR VPWR net1341 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ CPU.aluIn1\[14\] _05330_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__and2_1
Xhold55 _06313_ VGND VGND VPWR VPWR net1352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 _08250_ VGND VGND VPWR VPWR net1363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 _01715_ VGND VGND VPWR VPWR net1374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 _06360_ VGND VGND VPWR VPWR net1385 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _06651_ net2589 _07620_ VGND VGND VPWR VPWR _07627_ sky130_fd_sc_hd__mux2_1
X_13537__927 clknet_1_0__leaf__08438_ VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__inv_2
Xhold99 CPU.aluReg\[11\] VGND VGND VPWR VPWR net1396 sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ _06992_ _06997_ VGND VGND VPWR VPWR _06998_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_871 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17397__21 clknet_1_1__leaf__04985_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__inv_2
X_10872_ CPU.aluIn1\[9\] _06943_ _06914_ VGND VGND VPWR VPWR _06944_ sky130_fd_sc_hd__mux2_1
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12611_ _06603_ net1703 _07993_ VGND VGND VPWR VPWR _07997_ sky130_fd_sc_hd__mux2_1
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15330_ _03379_ _03387_ _03241_ VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__o21a_1
X_12542_ _07960_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15261_ CPU.registerFile\[19\]\[23\] CPU.registerFile\[18\]\[23\] _03157_ VGND VGND
+ VPWR VPWR _03320_ sky130_fd_sc_hd__mux2_1
X_12473_ _07923_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__clkbuf_1
X_17000_ CPU.registerFile\[15\]\[24\] CPU.registerFile\[14\]\[24\] _04550_ VGND VGND
+ VPWR VPWR _04703_ sky130_fd_sc_hd__mux2_1
X_11424_ _06774_ _07310_ VGND VGND VPWR VPWR _07311_ sky130_fd_sc_hd__nor2_4
X_15192_ CPU.registerFile\[30\]\[21\] CPU.registerFile\[31\]\[21\] _02887_ VGND VGND
+ VPWR VPWR _03253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_8 _03242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11355_ _07273_ VGND VGND VPWR VPWR _07274_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10306_ _05739_ _05737_ _05738_ VGND VGND VPWR VPWR _06594_ sky130_fd_sc_hd__and3b_4
XFILLER_0_104_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18951_ net725 _02471_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11286_ _07236_ _06775_ VGND VGND VPWR VPWR _07237_ sky130_fd_sc_hd__nor2_2
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13025_ _08216_ VGND VGND VPWR VPWR _08217_ sky130_fd_sc_hd__buf_4
X_17902_ clknet_leaf_26_clk _01430_ VGND VGND VPWR VPWR CPU.Bimm\[2\] sky130_fd_sc_hd__dfxtp_1
X_10237_ _05735_ _05736_ _05740_ VGND VGND VPWR VPWR _06557_ sky130_fd_sc_hd__and3_4
X_18882_ net656 _02402_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_17833_ net913 _01395_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_10168_ CPU.PC\[2\] _06197_ _05911_ _06490_ VGND VGND VPWR VPWR _06491_ sky130_fd_sc_hd__o22ai_2
X_17764_ net844 _01326_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_13745__1114 clknet_1_0__leaf__08459_ VGND VGND VPWR VPWR net1170 sky130_fd_sc_hd__inv_2
X_10099_ _05911_ _06424_ VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__nor2_1
X_14976_ CPU.registerFile\[20\]\[16\] _08839_ _03041_ _08841_ VGND VGND VPWR VPWR
+ _03042_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16715_ _04419_ _04420_ _04424_ _04383_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__a211o_1
X_17695_ CPU.mem_wdata\[1\] per_uart.d_in_uart\[1\] _05218_ VGND VGND VPWR VPWR _05221_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16646_ _04080_ _04081_ CPU.registerFile\[25\]\[15\] VGND VGND VPWR VPWR _04358_
+ sky130_fd_sc_hd__a21o_1
X_18585__42 VGND VGND VPWR VPWR _18585__42/HI net42 sky130_fd_sc_hd__conb_1
XFILLER_0_69_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12809_ _08100_ _08101_ _06869_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__o21a_1
X_16577_ _04175_ _04176_ CPU.registerFile\[17\]\[13\] VGND VGND VPWR VPWR _04291_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18316_ net137 _01844_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15528_ CPU.registerFile\[24\]\[30\] _08582_ _03579_ _08540_ VGND VGND VPWR VPWR
+ _03580_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18247_ net1258 _01775_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_15459_ CPU.registerFile\[15\]\[28\] CPU.registerFile\[14\]\[28\] _08560_ VGND VGND
+ VPWR VPWR _03513_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__04985_ _04985_ VGND VGND VPWR VPWR clknet_0__04985_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_115_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18178_ net1189 net1567 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold503 CPU.registerFile\[5\]\[26\] VGND VGND VPWR VPWR net1800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 CPU.registerFile\[11\]\[29\] VGND VGND VPWR VPWR net1811 sky130_fd_sc_hd__dlygate4sd3_1
X_17129_ CPU.registerFile\[22\]\[27\] CPU.registerFile\[23\]\[27\] _03761_ VGND VGND
+ VPWR VPWR _04829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold525 CPU.registerFile\[13\]\[8\] VGND VGND VPWR VPWR net1822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 CPU.registerFile\[7\]\[22\] VGND VGND VPWR VPWR net1833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold547 CPU.registerFile\[19\]\[23\] VGND VGND VPWR VPWR net1844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 CPU.registerFile\[18\]\[29\] VGND VGND VPWR VPWR net1855 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ CPU.PC\[11\] _05886_ VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__nor2_1
Xhold569 CPU.registerFile\[3\]\[0\] VGND VGND VPWR VPWR net1866 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08902_ CPU.rs2\[29\] _05247_ _05251_ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _06211_ _06216_ _05744_ VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1203 CPU.registerFile\[2\]\[17\] VGND VGND VPWR VPWR net2500 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1214 CPU.registerFile\[16\]\[13\] VGND VGND VPWR VPWR net2511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 CPU.registerFile\[12\]\[23\] VGND VGND VPWR VPWR net2522 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1236 CPU.registerFile\[1\]\[9\] VGND VGND VPWR VPWR net2533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 CPU.registerFile\[12\]\[31\] VGND VGND VPWR VPWR net2544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1258 CPU.registerFile\[14\]\[15\] VGND VGND VPWR VPWR net2555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 CPU.registerFile\[26\]\[12\] VGND VGND VPWR VPWR net2566 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09316_ CPU.aluIn1\[16\] _05544_ _05664_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09247_ _05597_ _05598_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09178_ CPU.Jimm\[12\] VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_16_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput12 net12 VGND VGND VPWR VPWR spi_mosi_ram sky130_fd_sc_hd__clkbuf_4
X_11140_ net1370 _07149_ VGND VGND VPWR VPWR _07152_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13805__1168 clknet_1_0__leaf__08465_ VGND VGND VPWR VPWR net1224 sky130_fd_sc_hd__inv_2
X_11071_ mapped_spi_flash.cmd_addr\[1\] _05714_ _06976_ VGND VGND VPWR VPWR _07104_
+ sky130_fd_sc_hd__mux2_1
X_10022_ _05263_ _05533_ _05536_ CPU.aluReg\[8\] _06350_ VGND VGND VPWR VPWR _06351_
+ sky130_fd_sc_hd__a221o_1
X_14830_ CPU.registerFile\[10\]\[12\] CPU.registerFile\[11\]\[12\] _02779_ VGND VGND
+ VPWR VPWR _02900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14761_ _02831_ _02832_ CPU.registerFile\[1\]\[10\] VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__a21o_1
X_11973_ _06634_ net2225 _07609_ VGND VGND VPWR VPWR _07618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16500_ CPU.registerFile\[16\]\[11\] _03848_ _04090_ _04215_ VGND VGND VPWR VPWR
+ _04216_ sky130_fd_sc_hd__o211a_1
X_10924_ net11 _06983_ _06985_ net2586 VGND VGND VPWR VPWR _06986_ sky130_fd_sc_hd__a22o_1
X_17480_ net13 VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__clkbuf_2
X_14692_ CPU.registerFile\[30\]\[9\] CPU.registerFile\[31\]\[9\] _08645_ VGND VGND
+ VPWR VPWR _02765_ sky130_fd_sc_hd__mux2_1
X_13318__818 clknet_1_1__leaf__08363_ VGND VGND VPWR VPWR net874 sky130_fd_sc_hd__inv_2
X_16431_ CPU.registerFile\[13\]\[10\] _03976_ VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10855_ CPU.aluIn1\[13\] _06930_ _06914_ VGND VGND VPWR VPWR _06931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19150_ clknet_leaf_5_clk net2200 VGND VGND VPWR VPWR per_uart.uart0.tx_bitcount\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16362_ _05690_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__clkbuf_4
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10786_ CPU.aluReg\[29\] _06877_ _06869_ VGND VGND VPWR VPWR _06878_ sky130_fd_sc_hd__mux2_1
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18101_ net1112 _01629_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[11\] sky130_fd_sc_hd__dfxtp_1
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12525_ _07950_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__clkbuf_1
X_15313_ _03202_ _03358_ _03362_ _03370_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__a31o_1
X_16293_ CPU.registerFile\[8\]\[7\] _08394_ _06150_ _04012_ VGND VGND VPWR VPWR _04013_
+ sky130_fd_sc_hd__o211a_1
X_19081_ clknet_leaf_27_clk _02601_ VGND VGND VPWR VPWR per_uart.uart0.rxd_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18032_ net1043 _01560_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_12456_ net1699 _07368_ _07906_ VGND VGND VPWR VPWR _07914_ sky130_fd_sc_hd__mux2_1
X_15244_ CPU.registerFile\[10\]\[22\] CPU.registerFile\[11\]\[22\] _03183_ VGND VGND
+ VPWR VPWR _03304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11407_ _07301_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15175_ _03235_ _03236_ CPU.registerFile\[1\]\[20\] VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12387_ _07877_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__03652_ _03652_ VGND VGND VPWR VPWR clknet_0__03652_ sky130_fd_sc_hd__clkbuf_16
X_11338_ CPU.registerFile\[2\]\[7\] _06386_ _07260_ VGND VGND VPWR VPWR _07265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18934_ net708 _02454_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_11269_ _06647_ net2124 _07223_ VGND VGND VPWR VPWR _07228_ sky130_fd_sc_hd__mux2_1
X_13008_ net1911 _07362_ _08203_ VGND VGND VPWR VPWR _08208_ sky130_fd_sc_hd__mux2_1
X_18865_ net639 _02385_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_14113__255 clknet_1_1__leaf__08496_ VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__inv_2
X_17816_ net896 _01378_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_18796_ net585 _02320_ VGND VGND VPWR VPWR CPU.aluReg\[26\] sky130_fd_sc_hd__dfxtp_1
X_17747_ net832 _01313_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_14959_ _03023_ _03024_ _03025_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17678_ _05672_ VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13727__1098 clknet_1_1__leaf__08457_ VGND VGND VPWR VPWR net1154 sky130_fd_sc_hd__inv_2
X_16629_ CPU.registerFile\[13\]\[15\] _03976_ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__or2_1
XFILLER_0_159_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09101_ _05452_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_162_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14007__160 clknet_1_0__leaf__08485_ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__inv_2
XFILLER_0_26_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09032_ CPU.aluIn1\[25\] _05383_ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold300 CPU.registerFile\[13\]\[27\] VGND VGND VPWR VPWR net1597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold311 CPU.cycles\[18\] VGND VGND VPWR VPWR net1608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold322 mapped_spi_flash.rcv_data\[12\] VGND VGND VPWR VPWR net1619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 mapped_spi_flash.rcv_bitcount\[0\] VGND VGND VPWR VPWR net1630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold344 _05851_ VGND VGND VPWR VPWR net1641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 mapped_spi_flash.state\[0\] VGND VGND VPWR VPWR net1652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 _05174_ VGND VGND VPWR VPWR net1663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 CPU.registerFile\[6\]\[7\] VGND VGND VPWR VPWR net1674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold388 CPU.registerFile\[19\]\[25\] VGND VGND VPWR VPWR net1685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 CPU.registerFile\[10\]\[31\] VGND VGND VPWR VPWR net1696 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09934_ _06266_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__buf_4
XFILLER_0_110_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09865_ net2365 _06200_ _06055_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__mux2_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1000 CPU.registerFile\[16\]\[2\] VGND VGND VPWR VPWR net2297 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 CPU.registerFile\[16\]\[7\] VGND VGND VPWR VPWR net2308 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1022 CPU.registerFile\[29\]\[26\] VGND VGND VPWR VPWR net2319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 CPU.registerFile\[27\]\[27\] VGND VGND VPWR VPWR net2330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 CPU.registerFile\[16\]\[27\] VGND VGND VPWR VPWR net2341 sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ _05346_ _05769_ _05770_ net1335 _06133_ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__a221o_2
Xhold1055 CPU.registerFile\[18\]\[11\] VGND VGND VPWR VPWR net2352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 CPU.registerFile\[16\]\[11\] VGND VGND VPWR VPWR net2363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1077 CPU.registerFile\[2\]\[11\] VGND VGND VPWR VPWR net2374 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1088 CPU.registerFile\[16\]\[21\] VGND VGND VPWR VPWR net2385 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03641_ clknet_0__03641_ VGND VGND VPWR VPWR clknet_1_0__leaf__03641_
+ sky130_fd_sc_hd__clkbuf_16
Xhold1099 CPU.registerFile\[16\]\[30\] VGND VGND VPWR VPWR net2396 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10640_ _06789_ VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10571_ net1813 _06083_ _06750_ VGND VGND VPWR VPWR _06752_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12310_ _07670_ _07671_ _07832_ net1298 VGND VGND VPWR VPWR _07833_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13744__1113 clknet_1_0__leaf__08459_ VGND VGND VPWR VPWR net1169 sky130_fd_sc_hd__inv_2
XFILLER_0_161_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12241_ net1429 _07785_ _07792_ _07755_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12172_ mapped_spi_ram.cmd_addr\[8\] _05704_ _07724_ VGND VGND VPWR VPWR _07744_
+ sky130_fd_sc_hd__mux2_1
X_11123_ mapped_spi_flash.rcv_data\[26\] _07135_ VGND VGND VPWR VPWR _07142_ sky130_fd_sc_hd__or2_1
X_16980_ CPU.registerFile\[27\]\[23\] CPU.registerFile\[26\]\[23\] _04646_ VGND VGND
+ VPWR VPWR _04684_ sky130_fd_sc_hd__mux2_1
X_11054_ CPU.PC\[6\] _07031_ _07090_ _06853_ VGND VGND VPWR VPWR _07091_ sky130_fd_sc_hd__o211a_1
X_10005_ _06202_ _06334_ _06177_ VGND VGND VPWR VPWR _06335_ sky130_fd_sc_hd__o21a_1
X_18650_ clknet_leaf_11_clk _02174_ VGND VGND VPWR VPWR CPU.rs2\[22\] sky130_fd_sc_hd__dfxtp_1
X_17601_ per_uart.d_in_uart\[0\] _05134_ _05157_ per_uart.uart0.txd_reg\[1\] VGND
+ VGND VPWR VPWR _05158_ sky130_fd_sc_hd__o22a_1
X_14813_ CPU.registerFile\[22\]\[12\] CPU.registerFile\[23\]\[12\] _08756_ VGND VGND
+ VPWR VPWR _02883_ sky130_fd_sc_hd__mux2_1
X_18581_ net402 net38 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_15793_ _03660_ _03664_ _08348_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__or3b_1
XFILLER_0_99_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17532_ _05069_ net2642 _05102_ _05103_ _06858_ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__o221a_1
XFILLER_0_98_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14744_ _08722_ _02810_ _02815_ _08851_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__o211a_1
X_11956_ _07597_ VGND VGND VPWR VPWR _07609_ sky130_fd_sc_hd__buf_4
X_17463_ _05045_ _05046_ _05020_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__a21oi_1
X_10907_ _05437_ _06861_ VGND VGND VPWR VPWR _06970_ sky130_fd_sc_hd__nor2_1
X_14675_ _08425_ _02727_ _02748_ _08597_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__a211o_1
X_11887_ _07572_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16414_ _04130_ _04131_ _03961_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10838_ CPU.aluIn1\[17\] _06917_ _06914_ VGND VGND VPWR VPWR _06918_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13370__864 clknet_1_0__leaf__08369_ VGND VGND VPWR VPWR net920 sky130_fd_sc_hd__inv_2
X_19133_ clknet_leaf_15_clk _02653_ VGND VGND VPWR VPWR CPU.PC\[15\] sky130_fd_sc_hd__dfxtp_2
X_16345_ CPU.registerFile\[6\]\[8\] CPU.registerFile\[7\]\[8\] _04022_ VGND VGND VPWR
+ VPWR _04064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10769_ CPU.aluReg\[31\] CPU.Bimm\[10\] _06862_ VGND VGND VPWR VPWR _06863_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12508_ _07941_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__clkbuf_1
X_19064_ net806 _02584_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[17\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__08490_ clknet_0__08490_ VGND VGND VPWR VPWR clknet_1_1__leaf__08490_
+ sky130_fd_sc_hd__clkbuf_16
X_16276_ CPU.registerFile\[24\]\[6\] _03915_ _03747_ _03996_ VGND VGND VPWR VPWR _03997_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18015_ net1026 _01543_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12439_ net1793 _07351_ _07895_ VGND VGND VPWR VPWR _07905_ sky130_fd_sc_hd__mux2_1
X_15227_ CPU.registerFile\[22\]\[22\] CPU.registerFile\[23\]\[22\] _02998_ VGND VGND
+ VPWR VPWR _03287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15158_ _02964_ _03214_ _03219_ _03092_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14109_ clknet_1_0__leaf__08495_ VGND VGND VPWR VPWR _08496_ sky130_fd_sc_hd__buf_1
X_15089_ _03143_ _03152_ _02837_ VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__o21a_2
XFILLER_0_129_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18917_ net691 _02437_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09650_ _05933_ _05993_ _05931_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__a21o_1
X_18848_ clknet_leaf_7_clk _02372_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_09581_ CPU.PC\[19\] _05924_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__xor2_2
XFILLER_0_54_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18779_ net568 _02303_ VGND VGND VPWR VPWR CPU.aluReg\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15926__665 clknet_1_1__leaf__03688_ VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__inv_2
XFILLER_0_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13804__1167 clknet_1_0__leaf__08465_ VGND VGND VPWR VPWR net1223 sky130_fd_sc_hd__inv_2
XFILLER_0_9_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09015_ _05359_ _05361_ _05366_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold130 mapped_spi_ram.rcv_data\[30\] VGND VGND VPWR VPWR net1427 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold141 mapped_spi_flash.rcv_data\[27\] VGND VGND VPWR VPWR net1438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 per_uart.uart0.txd_reg\[7\] VGND VGND VPWR VPWR net1449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 mapped_spi_ram.cmd_addr\[11\] VGND VGND VPWR VPWR net1460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 mapped_spi_ram.cmd_addr\[12\] VGND VGND VPWR VPWR net1471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 mapped_spi_ram.rcv_data\[12\] VGND VGND VPWR VPWR net1482 sky130_fd_sc_hd__dlygate4sd3_1
X_13933__93 clknet_1_1__leaf__08478_ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__inv_2
Xhold196 mapped_spi_flash.cmd_addr\[15\] VGND VGND VPWR VPWR net1493 sky130_fd_sc_hd__dlygate4sd3_1
X_09917_ _05526_ _05550_ _05553_ CPU.cycles\[12\] VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__a22o_1
X_17313__727 clknet_1_1__leaf__04981_ VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__inv_2
X_15671__468 clknet_1_1__leaf__03645_ VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__inv_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09848_ _05468_ _06183_ _05333_ VGND VGND VPWR VPWR _06184_ sky130_fd_sc_hd__o21ai_2
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _05514_ _05357_ _05520_ _06115_ _06117_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__a311o_1
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ net2030 _07322_ _07526_ VGND VGND VPWR VPWR _07532_ sky130_fd_sc_hd__mux2_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _08091_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__clkbuf_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _07495_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__clkbuf_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19195__53 VGND VGND VPWR VPWR _19195__53/HI net53 sky130_fd_sc_hd__conb_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11672_ _07458_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__clkbuf_1
X_14460_ CPU.registerFile\[5\]\[3\] CPU.registerFile\[4\]\[3\] _08576_ VGND VGND VPWR
+ VPWR _08703_ sky130_fd_sc_hd__mux2_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10623_ _06780_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__clkbuf_1
X_13411_ _08384_ VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14391_ _08425_ _08616_ _08635_ _08597_ VGND VGND VPWR VPWR _08636_ sky130_fd_sc_hd__a211o_1
XFILLER_0_119_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_21_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_16
X_16130_ _06855_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__clkbuf_4
X_10554_ net2035 _05805_ _06739_ VGND VGND VPWR VPWR _06743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13999__152 clknet_1_1__leaf__08485_ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__inv_2
XFILLER_0_161_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16061_ CPU.registerFile\[6\]\[1\] CPU.registerFile\[7\]\[1\] _03717_ VGND VGND VPWR
+ VPWR _03787_ sky130_fd_sc_hd__mux2_1
X_13273_ per_uart.uart0.enable16_counter\[9\] _08353_ VGND VGND VPWR VPWR _08354_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_161_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10485_ net2137 _05805_ _06702_ VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__mux2_1
X_12224_ mapped_spi_ram.rcv_bitcount\[2\] mapped_spi_ram.rcv_bitcount\[1\] mapped_spi_ram.rcv_bitcount\[0\]
+ VGND VGND VPWR VPWR _07780_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15012_ _02751_ _03074_ _03076_ _02759_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__a211o_1
XFILLER_0_121_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12155_ _07715_ _07731_ VGND VGND VPWR VPWR _07732_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13726__1097 clknet_1_0__leaf__08457_ VGND VGND VPWR VPWR net1153 sky130_fd_sc_hd__inv_2
X_11106_ mapped_spi_flash.state\[3\] VGND VGND VPWR VPWR _07130_ sky130_fd_sc_hd__inv_2
X_16963_ _04503_ _04664_ _04666_ _04509_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__a211o_1
X_12086_ net10 VGND VGND VPWR VPWR _07683_ sky130_fd_sc_hd__inv_2
X_18702_ net491 _02226_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[2\] sky130_fd_sc_hd__dfxtp_1
X_11037_ _07025_ _05601_ VGND VGND VPWR VPWR _07076_ sky130_fd_sc_hd__and2_1
X_16894_ _04389_ _04390_ CPU.registerFile\[1\]\[21\] VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__a21o_1
X_17288__704 clknet_1_1__leaf__04979_ VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__inv_2
X_18633_ clknet_leaf_17_clk _02157_ VGND VGND VPWR VPWR CPU.mem_wdata\[5\] sky130_fd_sc_hd__dfxtp_2
X_18564_ net385 net21 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_12988_ _08197_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__clkbuf_1
X_15648__448 clknet_1_1__leaf__03642_ VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__inv_2
X_17515_ _05088_ _05089_ _05058_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__a21oi_1
X_14727_ CPU.registerFile\[19\]\[10\] CPU.registerFile\[18\]\[10\] _02753_ VGND VGND
+ VPWR VPWR _02799_ sky130_fd_sc_hd__mux2_1
X_18495_ net316 _02019_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_11939_ _07600_ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14225__356 clknet_1_1__leaf__08507_ VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__inv_2
XFILLER_0_157_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17446_ _05016_ CPU.PC\[4\] _05032_ _05033_ _07002_ VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__o221a_1
XFILLER_0_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14658_ CPU.registerFile\[10\]\[8\] CPU.registerFile\[11\]\[8\] _08564_ VGND VGND
+ VPWR VPWR _02732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13609_ clknet_1_0__leaf__08440_ VGND VGND VPWR VPWR _08446_ sky130_fd_sc_hd__buf_1
XFILLER_0_83_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17377_ _04996_ _05003_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14589_ _08785_ _08826_ _08828_ _08590_ VGND VGND VPWR VPWR _08829_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_12_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19116_ net99 _02636_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_16328_ _03770_ _03771_ CPU.registerFile\[17\]\[7\] VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19047_ net789 _02567_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_16259_ _03703_ _03975_ _03978_ _03979_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_1__f__08473_ clknet_0__08473_ VGND VGND VPWR VPWR clknet_1_1__leaf__08473_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14119__261 clknet_1_1__leaf__08496_ VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__inv_2
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09702_ _06017_ _06043_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09633_ _05943_ _05975_ _05976_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__a21o_1
X_13743__1112 clknet_1_0__leaf__08459_ VGND VGND VPWR VPWR net1168 sky130_fd_sc_hd__inv_2
X_09564_ _05881_ _05895_ _05540_ _05907_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_78_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09495_ mapped_spi_ram.rcv_data\[1\] _05761_ _05762_ net1640 VGND VGND VPWR VPWR
+ _05841_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15707__501 clknet_1_1__leaf__03648_ VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__inv_2
XFILLER_0_77_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10270_ net1689 _06169_ _06569_ VGND VGND VPWR VPWR _06575_ sky130_fd_sc_hd__mux2_1
X_12911_ _06054_ net2447 _08156_ VGND VGND VPWR VPWR _08157_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__08493_ clknet_0__08493_ VGND VGND VPWR VPWR clknet_1_0__leaf__08493_
+ sky130_fd_sc_hd__clkbuf_16
X_15630_ clknet_1_0__leaf__08506_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__buf_1
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _08108_ VGND VGND VPWR VPWR _08120_ sky130_fd_sc_hd__buf_4
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ CPU.registerFile\[28\]\[31\] CPU.registerFile\[29\]\[31\] _08410_ VGND VGND
+ VPWR VPWR _03612_ sky130_fd_sc_hd__mux2_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _08082_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__clkbuf_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ CPU.registerFile\[17\]\[5\] _06456_ VGND VGND VPWR VPWR _08753_ sky130_fd_sc_hd__or2_1
X_11724_ _07485_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__clkbuf_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18280_ net1291 _01808_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_15492_ _08580_ _03542_ _03544_ _03218_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__a211o_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _04926_ _04927_ _06535_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__mux2_1
X_11655_ _07448_ VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14443_ _08410_ VGND VGND VPWR VPWR _08686_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17162_ CPU.registerFile\[24\]\[28\] _03724_ _04569_ _04860_ VGND VGND VPWR VPWR
+ _04861_ sky130_fd_sc_hd__o211a_1
X_10606_ net1880 _06486_ _06761_ VGND VGND VPWR VPWR _06770_ sky130_fd_sc_hd__mux2_1
X_14374_ _08617_ _08618_ _08562_ VGND VGND VPWR VPWR _08619_ sky130_fd_sc_hd__mux2_1
X_11586_ _07411_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16113_ CPU.registerFile\[27\]\[2\] CPU.registerFile\[26\]\[2\] _03837_ VGND VGND
+ VPWR VPWR _03838_ sky130_fd_sc_hd__mux2_1
X_10537_ net2013 _06486_ _06724_ VGND VGND VPWR VPWR _06733_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17093_ CPU.registerFile\[22\]\[26\] CPU.registerFile\[23\]\[26\] _03761_ VGND VGND
+ VPWR VPWR _04794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16044_ _03750_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__clkbuf_4
X_10468_ _06655_ net2409 _06687_ VGND VGND VPWR VPWR _06696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12207_ _07670_ _07671_ _07767_ _07749_ VGND VGND VPWR VPWR _07768_ sky130_fd_sc_hd__a22o_1
X_13187_ net1616 _08303_ VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__xor2_1
X_10399_ _06657_ net1733 _06639_ VGND VGND VPWR VPWR _06658_ sky130_fd_sc_hd__mux2_1
X_12138_ mapped_spi_ram.cmd_addr\[18\] _07045_ _07704_ VGND VGND VPWR VPWR _07720_
+ sky130_fd_sc_hd__mux2_1
X_15654__452 clknet_1_1__leaf__03644_ VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__inv_2
X_13803__1166 clknet_1_1__leaf__08465_ VGND VGND VPWR VPWR net1222 sky130_fd_sc_hd__inv_2
X_17995_ net1006 _01523_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_13912__74 clknet_1_1__leaf__08476_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__inv_2
X_12069_ net2055 _07376_ _07634_ VGND VGND VPWR VPWR _07669_ sky130_fd_sc_hd__mux2_1
X_16946_ _04479_ _04645_ _04650_ _04446_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_1_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_126_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16877_ _06109_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__clkbuf_4
X_18616_ net437 _02140_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13376__870 clknet_1_1__leaf__08369_ VGND VGND VPWR VPWR net926 sky130_fd_sc_hd__inv_2
XFILLER_0_48_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18547_ net368 _02071_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09280_ _05630_ _05631_ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__nor2_1
X_18478_ net299 _02002_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17429_ CPU.PC\[2\] _08311_ _08331_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__or3_1
XFILLER_0_142_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08456_ clknet_0__08456_ VGND VGND VPWR VPWR clknet_1_1__leaf__08456_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__08487_ _08487_ VGND VGND VPWR VPWR clknet_0__08487_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14052__201 clknet_1_0__leaf__08489_ VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__inv_2
X_08995_ _05340_ _05346_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09616_ CPU.PC\[3\] _05958_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09547_ CPU.PC\[17\] _05890_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__and2_1
X_17412__34 clknet_1_1__leaf__05014_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__inv_2
XFILLER_0_148_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09478_ net2341 _05825_ _05742_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__mux2_1
X_13725__1096 clknet_1_0__leaf__08457_ VGND VGND VPWR VPWR net1152 sky130_fd_sc_hd__inv_2
XFILLER_0_148_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11440_ _05838_ VGND VGND VPWR VPWR _07322_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11371_ _07282_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10322_ _06605_ net1848 _06597_ VGND VGND VPWR VPWR _06606_ sky130_fd_sc_hd__mux2_1
X_13110_ _08254_ _08260_ _08261_ _08253_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_132_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13041_ net1380 VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__clkbuf_1
X_10253_ net1678 _05873_ _06558_ VGND VGND VPWR VPWR _06566_ sky130_fd_sc_hd__mux2_1
X_14254__382 clknet_1_0__leaf__08510_ VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__inv_2
X_10184_ CPU.cycles\[2\] _05759_ _06491_ net1422 VGND VGND VPWR VPWR _06507_ sky130_fd_sc_hd__a211o_2
X_16800_ CPU.registerFile\[8\]\[19\] _04505_ _04506_ _04507_ VGND VGND VPWR VPWR _04508_
+ sky130_fd_sc_hd__o211a_1
X_17780_ net860 _01342_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_14992_ _03056_ _03057_ _02937_ VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__mux2_1
X_16731_ _08396_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16662_ _04141_ _04353_ _04373_ _04096_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__a211o_1
XFILLER_0_159_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18401_ net222 _01929_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[1\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__08476_ clknet_0__08476_ VGND VGND VPWR VPWR clknet_1_0__leaf__08476_
+ sky130_fd_sc_hd__clkbuf_16
X_13514__906 clknet_1_1__leaf__08436_ VGND VGND VPWR VPWR net962 sky130_fd_sc_hd__inv_2
X_12825_ _08111_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__clkbuf_1
X_16593_ CPU.registerFile\[6\]\[14\] CPU.registerFile\[7\]\[14\] _04022_ VGND VGND
+ VPWR VPWR _04306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18332_ net153 _01860_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15544_ _08567_ _08569_ CPU.registerFile\[1\]\[30\] VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__a21o_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _08073_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11707_ net2342 _07356_ _07475_ VGND VGND VPWR VPWR _07477_ sky130_fd_sc_hd__mux2_1
X_18263_ net1274 _01791_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15475_ _03520_ _03528_ _03241_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__o21a_1
X_12687_ _06611_ net2469 _08029_ VGND VGND VPWR VPWR _08037_ sky130_fd_sc_hd__mux2_1
X_17214_ CPU.registerFile\[8\]\[30\] _03707_ _03708_ _04910_ VGND VGND VPWR VPWR _04911_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14426_ _08581_ _08667_ _08669_ _08590_ VGND VGND VPWR VPWR _08670_ sky130_fd_sc_hd__a211o_1
X_11638_ net1994 _07356_ _07438_ VGND VGND VPWR VPWR _07440_ sky130_fd_sc_hd__mux2_1
X_18194_ net1205 _01722_ VGND VGND VPWR VPWR mapped_spi_ram.snd_bitcount\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17145_ CPU.registerFile\[13\]\[28\] _03767_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14357_ _08415_ _08599_ _08601_ _08420_ VGND VGND VPWR VPWR _08602_ sky130_fd_sc_hd__a211o_1
X_11569_ net1901 _07356_ _07401_ VGND VGND VPWR VPWR _07403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold707 CPU.registerFile\[29\]\[13\] VGND VGND VPWR VPWR net2004 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold718 CPU.registerFile\[17\]\[27\] VGND VGND VPWR VPWR net2015 sky130_fd_sc_hd__dlygate4sd3_1
X_17076_ CPU.registerFile\[6\]\[26\] CPU.registerFile\[7\]\[26\] _04426_ VGND VGND
+ VPWR VPWR _04777_ sky130_fd_sc_hd__mux2_1
Xhold729 per_uart.uart0.tx_bitcount\[2\] VGND VGND VPWR VPWR net2026 sky130_fd_sc_hd__dlygate4sd3_1
X_14288_ _08521_ _08524_ _08531_ _08533_ VGND VGND VPWR VPWR _08534_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__08341_ _08341_ VGND VGND VPWR VPWR clknet_0__08341_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_733 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16027_ _03702_ _03746_ _03753_ _08400_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17978_ net989 _01506_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16929_ CPU.registerFile\[5\]\[22\] CPU.registerFile\[4\]\[22\] _04428_ VGND VGND
+ VPWR VPWR _04634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09401_ _05414_ _05510_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09332_ _05659_ _05678_ _05679_ _05683_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__a211o_1
XFILLER_0_158_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09263_ _05613_ _05614_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09194_ _05422_ _05538_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1__f__08508_ clknet_0__08508_ VGND VGND VPWR VPWR clknet_1_1__leaf__08508_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08439_ clknet_0__08439_ VGND VGND VPWR VPWR clknet_1_1__leaf__08439_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold12 _01726_ VGND VGND VPWR VPWR net1309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 mapped_spi_ram.div_counter\[0\] VGND VGND VPWR VPWR net1320 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ CPU.rs2\[14\] _05245_ _05249_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__o21a_1
Xhold34 CPU.aluReg\[9\] VGND VGND VPWR VPWR net1331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 _01734_ VGND VGND VPWR VPWR net1342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 _06315_ VGND VGND VPWR VPWR net1353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 per_uart.uart0.uart_rxd1 VGND VGND VPWR VPWR net1364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 mapped_spi_flash.rcv_data\[30\] VGND VGND VPWR VPWR net1375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 _08243_ VGND VGND VPWR VPWR net1386 sky130_fd_sc_hd__dlygate4sd3_1
X_15865__611 clknet_1_1__leaf__03681_ VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__inv_2
XFILLER_0_97_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10940_ mapped_spi_flash.cmd_addr\[26\] _06983_ _06985_ mapped_spi_flash.cmd_addr\[25\]
+ VGND VGND VPWR VPWR _06997_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10871_ CPU.aluReg\[10\] CPU.aluReg\[8\] _06939_ VGND VGND VPWR VPWR _06943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12610_ _07996_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__clkbuf_1
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13963__121 clknet_1_1__leaf__08480_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__inv_2
X_12541_ net2368 _07316_ _07957_ VGND VGND VPWR VPWR _07960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13802__1165 clknet_1_1__leaf__08465_ VGND VGND VPWR VPWR net1221 sky130_fd_sc_hd__inv_2
X_15260_ net1644 _03201_ _03319_ _02993_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12472_ net1811 _07316_ _07920_ VGND VGND VPWR VPWR _07923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11423_ _05739_ _05737_ _05738_ VGND VGND VPWR VPWR _07310_ sky130_fd_sc_hd__or3b_4
XFILLER_0_105_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15191_ _03078_ _03249_ _03251_ _03043_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__a211o_1
X_14059__207 clknet_1_0__leaf__08490_ VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__inv_2
XANTENNA_9 _03354_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14142_ clknet_1_0__leaf__08495_ VGND VGND VPWR VPWR _08499_ sky130_fd_sc_hd__buf_1
XFILLER_0_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11354_ _06813_ _07199_ VGND VGND VPWR VPWR _07273_ sky130_fd_sc_hd__nor2b_4
X_10305_ _05733_ VGND VGND VPWR VPWR _06593_ sky130_fd_sc_hd__clkbuf_4
X_11285_ _05736_ CPU.writeBack _05735_ VGND VGND VPWR VPWR _07236_ sky130_fd_sc_hd__nand3b_4
X_18950_ net724 _02470_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13024_ _06813_ _07310_ VGND VGND VPWR VPWR _08216_ sky130_fd_sc_hd__nor2_4
X_17901_ clknet_leaf_22_clk _01429_ VGND VGND VPWR VPWR CPU.Bimm\[1\] sky130_fd_sc_hd__dfxtp_2
X_10236_ _06556_ VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__clkbuf_1
X_18881_ net655 _02401_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_17832_ net912 _01394_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_10167_ _06488_ _06489_ VGND VGND VPWR VPWR _06490_ sky130_fd_sc_hd__xor2_1
X_17763_ net843 _01325_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_10098_ _06423_ _05963_ VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__xor2_1
X_14975_ CPU.registerFile\[21\]\[16\] _02960_ VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__or2_1
X_16714_ CPU.registerFile\[12\]\[17\] _04421_ _04422_ _04423_ VGND VGND VPWR VPWR
+ _04424_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17694_ _05220_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16645_ CPU.registerFile\[27\]\[15\] CPU.registerFile\[26\]\[15\] _04242_ VGND VGND
+ VPWR VPWR _04357_ sky130_fd_sc_hd__mux2_1
X_15766__553 clknet_1_0__leaf__03655_ VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__08459_ clknet_0__08459_ VGND VGND VPWR VPWR clknet_1_0__leaf__08459_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12808_ _05287_ _06864_ VGND VGND VPWR VPWR _08101_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16576_ CPU.registerFile\[19\]\[13\] CPU.registerFile\[18\]\[13\] _03923_ VGND VGND
+ VPWR VPWR _04290_ sky130_fd_sc_hd__mux2_1
X_18315_ net136 _01843_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15527_ _08566_ _08568_ CPU.registerFile\[25\]\[30\] VGND VGND VPWR VPWR _03579_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12739_ _06663_ _07633_ VGND VGND VPWR VPWR _08064_ sky130_fd_sc_hd__nand2_4
XFILLER_0_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18246_ net1257 _01774_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15458_ _03202_ _03499_ _03503_ _03511_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__a31o_1
Xclkbuf_0__04984_ _04984_ VGND VGND VPWR VPWR clknet_0__04984_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_154_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14409_ _08535_ _08648_ _08652_ _08554_ VGND VGND VPWR VPWR _08653_ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18177_ net1188 net1537 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[16\] sky130_fd_sc_hd__dfxtp_1
X_15389_ _03443_ _03444_ _08541_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__mux2_1
X_17128_ _04479_ _04823_ _04827_ _08403_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__o211a_1
Xhold504 CPU.registerFile\[21\]\[12\] VGND VGND VPWR VPWR net1801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 mapped_spi_flash.rcv_data\[11\] VGND VGND VPWR VPWR net1812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold526 CPU.registerFile\[10\]\[24\] VGND VGND VPWR VPWR net1823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 CPU.registerFile\[10\]\[9\] VGND VGND VPWR VPWR net1834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold548 CPU.registerFile\[20\]\[24\] VGND VGND VPWR VPWR net1845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 CPU.registerFile\[5\]\[4\] VGND VGND VPWR VPWR net1856 sky130_fd_sc_hd__dlygate4sd3_1
X_17059_ _04759_ _04760_ _03742_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__mux2_1
X_09950_ _06281_ _05975_ VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08901_ CPU.aluIn1\[30\] _05252_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__and2_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _05333_ _05523_ _06215_ VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__o21ai_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13724__1095 clknet_1_0__leaf__08457_ VGND VGND VPWR VPWR net1151 sky130_fd_sc_hd__inv_2
XFILLER_0_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13341__839 clknet_1_1__leaf__08365_ VGND VGND VPWR VPWR net895 sky130_fd_sc_hd__inv_2
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1204 CPU.registerFile\[2\]\[15\] VGND VGND VPWR VPWR net2501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1215 CPU.registerFile\[12\]\[27\] VGND VGND VPWR VPWR net2512 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 CPU.registerFile\[14\]\[20\] VGND VGND VPWR VPWR net2523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 CPU.registerFile\[7\]\[5\] VGND VGND VPWR VPWR net2534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 CPU.registerFile\[2\]\[14\] VGND VGND VPWR VPWR net2545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1259 CPU.registerFile\[23\]\[25\] VGND VGND VPWR VPWR net2556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09315_ CPU.PC\[16\] _05636_ _05666_ _05235_ VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09246_ CPU.aluIn1\[10\] CPU.Bimm\[10\] VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09177_ CPU.aluIn1\[31\] _05525_ _05528_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13543__932 clknet_1_0__leaf__08439_ VGND VGND VPWR VPWR net988 sky130_fd_sc_hd__inv_2
XFILLER_0_102_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11070_ net1492 _07054_ _07103_ _07069_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__o211a_1
X_10021_ _05266_ _05749_ VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__nor2_1
X_14760_ _08568_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__clkbuf_4
X_11972_ _07617_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__clkbuf_1
X_14030__181 clknet_1_1__leaf__08487_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__inv_2
X_10923_ _06984_ VGND VGND VPWR VPWR _06985_ sky130_fd_sc_hd__clkbuf_4
X_14691_ _08837_ _02761_ _02763_ _08802_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__a211o_1
X_16430_ CPU.registerFile\[15\]\[10\] CPU.registerFile\[14\]\[10\] _04146_ VGND VGND
+ VPWR VPWR _04147_ sky130_fd_sc_hd__mux2_1
X_13642_ clknet_1_0__leaf__08440_ VGND VGND VPWR VPWR _08449_ sky130_fd_sc_hd__buf_1
X_10854_ CPU.aluReg\[14\] CPU.aluReg\[12\] _06906_ VGND VGND VPWR VPWR _06930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16361_ _05689_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__clkbuf_4
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10785_ CPU.aluIn1\[29\] _06876_ _06861_ VGND VGND VPWR VPWR _06877_ sky130_fd_sc_hd__mux2_1
X_18100_ net1111 _01628_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[10\] sky130_fd_sc_hd__dfxtp_1
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15312_ _06013_ _03365_ _03369_ _03092_ VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__o211a_1
X_12524_ net2063 _07368_ _07942_ VGND VGND VPWR VPWR _07950_ sky130_fd_sc_hd__mux2_1
X_19080_ clknet_leaf_27_clk _02600_ VGND VGND VPWR VPWR per_uart.uart0.rxd_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16292_ CPU.registerFile\[9\]\[7\] _03698_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__or2_1
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18031_ net1042 _01559_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_15243_ _03301_ _03302_ _02937_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12455_ _07913_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11406_ net1726 _06386_ _07296_ VGND VGND VPWR VPWR _07301_ sky130_fd_sc_hd__mux2_1
X_15174_ _08568_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__clkbuf_4
X_12386_ _06651_ net1859 _07870_ VGND VGND VPWR VPWR _07877_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__03651_ _03651_ VGND VGND VPWR VPWR clknet_0__03651_ sky130_fd_sc_hd__clkbuf_16
X_11337_ _07264_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__clkbuf_1
X_18933_ net707 _02453_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11268_ _07227_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13007_ _08207_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__clkbuf_1
X_10219_ _06532_ _06533_ _06536_ _06539_ VGND VGND VPWR VPWR _06540_ sky130_fd_sc_hd__o211a_1
X_18864_ net638 _02384_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_11199_ _07182_ net1487 _07188_ VGND VGND VPWR VPWR _07189_ sky130_fd_sc_hd__mux2_1
X_17815_ net895 _01377_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_18795_ net584 _02319_ VGND VGND VPWR VPWR CPU.aluReg\[25\] sky130_fd_sc_hd__dfxtp_1
X_17746_ net831 _01312_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_14958_ _08540_ VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__buf_4
X_13909_ clknet_1_1__leaf__08473_ VGND VGND VPWR VPWR _08476_ sky130_fd_sc_hd__buf_1
XFILLER_0_134_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17677_ _06854_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__buf_2
X_14889_ CPU.registerFile\[16\]\[14\] _02755_ _02956_ _02757_ VGND VGND VPWR VPWR
+ _02957_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16628_ CPU.registerFile\[15\]\[15\] CPU.registerFile\[14\]\[15\] _04146_ VGND VGND
+ VPWR VPWR _04340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16559_ CPU.registerFile\[0\]\[13\] _04233_ _04068_ _04272_ VGND VGND VPWR VPWR _04273_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09100_ _05314_ _05313_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09031_ CPU.rs2\[25\] _05247_ _05251_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__o21a_1
X_18229_ net1240 _01757_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold301 per_uart.uart0.enable16_counter\[13\] VGND VGND VPWR VPWR net1598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 CPU.cycles\[1\] VGND VGND VPWR VPWR net1609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 CPU.cycles\[16\] VGND VGND VPWR VPWR net1620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 per_uart.uart0.rx_bitcount\[2\] VGND VGND VPWR VPWR net1631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 _08224_ VGND VGND VPWR VPWR net1642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 _06852_ VGND VGND VPWR VPWR net1653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold367 CPU.registerFile\[24\]\[1\] VGND VGND VPWR VPWR net1664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 CPU.registerFile\[10\]\[28\] VGND VGND VPWR VPWR net1675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 CPU.registerFile\[5\]\[23\] VGND VGND VPWR VPWR net1686 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ _06249_ _06250_ _06261_ _06265_ VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__or4b_4
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _06199_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__buf_4
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801__1164 clknet_1_1__leaf__08465_ VGND VGND VPWR VPWR net1220 sky130_fd_sc_hd__inv_2
Xhold1001 CPU.registerFile\[16\]\[6\] VGND VGND VPWR VPWR net2298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 CPU.registerFile\[14\]\[5\] VGND VGND VPWR VPWR net2309 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 CPU.registerFile\[24\]\[28\] VGND VGND VPWR VPWR net2320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1034 CPU.registerFile\[14\]\[1\] VGND VGND VPWR VPWR net2331 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ _05818_ _06129_ _06131_ _06132_ _05358_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__a32o_1
Xhold1045 CPU.registerFile\[8\]\[10\] VGND VGND VPWR VPWR net2342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1056 CPU.registerFile\[8\]\[8\] VGND VGND VPWR VPWR net2353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 CPU.registerFile\[1\]\[19\] VGND VGND VPWR VPWR net2364 sky130_fd_sc_hd__dlygate4sd3_1
X_14088__233 clknet_1_1__leaf__08493_ VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__inv_2
Xhold1078 CPU.registerFile\[12\]\[20\] VGND VGND VPWR VPWR net2375 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03640_ clknet_0__03640_ VGND VGND VPWR VPWR clknet_1_0__leaf__03640_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1089 CPU.registerFile\[2\]\[10\] VGND VGND VPWR VPWR net2386 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10570_ _06751_ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09229_ _05577_ _05579_ _05580_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_91_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12240_ mapped_spi_ram.rcv_data\[27\] _07787_ VGND VGND VPWR VPWR _07792_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12171_ net1490 _07738_ _07743_ _07737_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11122_ net1591 _07133_ _07141_ _07138_ VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__o211a_1
Xhold890 CPU.registerFile\[23\]\[4\] VGND VGND VPWR VPWR net2187 sky130_fd_sc_hd__dlygate4sd3_1
X_13324__823 clknet_1_0__leaf__08364_ VGND VGND VPWR VPWR net879 sky130_fd_sc_hd__inv_2
X_11053_ _07082_ _07089_ _07031_ VGND VGND VPWR VPWR _07090_ sky130_fd_sc_hd__o21ai_1
X_10004_ _05855_ _06203_ _05841_ _06204_ _06333_ VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__o32a_1
X_17600_ _05156_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__clkbuf_4
X_14812_ _02751_ _02879_ _02881_ _02759_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__a211o_1
X_18580_ net401 net37 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_15792_ per_uart.uart0.enable16_counter\[3\] _08347_ VGND VGND VPWR VPWR _03664_
+ sky130_fd_sc_hd__and2_1
X_17531_ _08335_ _06070_ _05073_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__o21ai_1
X_14743_ _08764_ _02811_ _02813_ _02814_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11955_ _07608_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17462_ _08311_ _06357_ _08331_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__or3_1
X_10906_ _06969_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__clkbuf_1
X_14674_ _02738_ _02747_ _08594_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__o21a_2
XFILLER_0_58_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11886_ _06615_ net1820 _07562_ VGND VGND VPWR VPWR _07572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16413_ CPU.registerFile\[20\]\[9\] CPU.registerFile\[21\]\[9\] _03883_ VGND VGND
+ VPWR VPWR _04131_ sky130_fd_sc_hd__mux2_1
X_10837_ CPU.aluReg\[18\] CPU.aluReg\[16\] _06906_ VGND VGND VPWR VPWR _06917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15843__591 clknet_1_1__leaf__03679_ VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__inv_2
X_19132_ clknet_leaf_16_clk _02652_ VGND VGND VPWR VPWR CPU.PC\[14\] sky130_fd_sc_hd__dfxtp_2
X_16344_ _04015_ _04060_ _04062_ _03979_ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__a211o_1
X_13723__1094 clknet_1_1__leaf__08457_ VGND VGND VPWR VPWR net1150 sky130_fd_sc_hd__inv_2
XFILLER_0_82_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10768_ _05799_ _05534_ VGND VGND VPWR VPWR _06862_ sky130_fd_sc_hd__nand2_1
X_18570__27 VGND VGND VPWR VPWR _18570__27/HI net27 sky130_fd_sc_hd__conb_1
XFILLER_0_137_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12507_ net2228 _07351_ _07931_ VGND VGND VPWR VPWR _07941_ sky130_fd_sc_hd__mux2_1
X_19063_ net805 _02583_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_16275_ _03749_ _03751_ CPU.registerFile\[25\]\[6\] VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__a21o_1
X_13487_ clknet_1_1__leaf__08366_ VGND VGND VPWR VPWR _08434_ sky130_fd_sc_hd__buf_1
X_10699_ net1810 _05839_ _06816_ VGND VGND VPWR VPWR _06822_ sky130_fd_sc_hd__mux2_1
X_18014_ net1025 _01542_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_15226_ _03156_ _03283_ _03285_ _03163_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__a211o_1
XFILLER_0_152_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12438_ _07904_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15157_ _03006_ _03215_ _03217_ _03218_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12369_ _06634_ net1790 _07859_ VGND VGND VPWR VPWR _07868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14108_ clknet_1_1__leaf__08339_ VGND VGND VPWR VPWR _08495_ sky130_fd_sc_hd__buf_1
X_15088_ _02826_ _03146_ _03150_ _03151_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__o211a_1
X_18916_ net690 _02436_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_14037__187 clknet_1_1__leaf__08488_ VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__inv_2
XFILLER_0_38_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18847_ clknet_leaf_7_clk net1542 VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_09580_ CPU.Jimm\[19\] _05921_ _05923_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__a21o_1
X_18778_ net567 _02302_ VGND VGND VPWR VPWR CPU.aluReg\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17729_ net814 _01295_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15625__427 clknet_1_0__leaf__03640_ VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__inv_2
XFILLER_0_162_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09014_ _05365_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__clkbuf_2
X_13918__80 clknet_1_1__leaf__08476_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__inv_2
XFILLER_0_115_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold120 _06223_ VGND VGND VPWR VPWR net1417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold131 _01720_ VGND VGND VPWR VPWR net1428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_950 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold142 _06484_ VGND VGND VPWR VPWR net1439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 _02680_ VGND VGND VPWR VPWR net1450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 mapped_spi_ram.rcv_data\[10\] VGND VGND VPWR VPWR net1461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 mapped_spi_ram.cmd_addr\[15\] VGND VGND VPWR VPWR net1472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 _01702_ VGND VGND VPWR VPWR net1483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 mapped_spi_flash.cmd_addr\[12\] VGND VGND VPWR VPWR net1494 sky130_fd_sc_hd__dlygate4sd3_1
X_09916_ _06202_ _06248_ _06177_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__o21a_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09847_ _06181_ _06182_ _05457_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__a21boi_2
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _05354_ _05531_ _05534_ CPU.aluReg\[18\] _06116_ VGND VGND VPWR VPWR _06117_
+ sky130_fd_sc_hd__a221o_1
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _06605_ net1984 _07490_ VGND VGND VPWR VPWR _07495_ sky130_fd_sc_hd__mux2_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ net2070 _07320_ _07453_ VGND VGND VPWR VPWR _07458_ sky130_fd_sc_hd__mux2_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ _05736_ _06364_ _00000_ VGND VGND VPWR VPWR _08384_ sky130_fd_sc_hd__mux2_1
X_10622_ net2516 _05786_ _06777_ VGND VGND VPWR VPWR _06780_ sky130_fd_sc_hd__mux2_1
X_14390_ _08625_ _08634_ _08594_ VGND VGND VPWR VPWR _08635_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10553_ _06742_ VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16060_ _03703_ _03783_ _03785_ _03714_ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__a211o_1
X_13272_ net1610 _08352_ VGND VGND VPWR VPWR _08353_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10484_ _06705_ VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15011_ CPU.registerFile\[16\]\[17\] _02755_ _03075_ _02757_ VGND VGND VPWR VPWR
+ _03076_ sky130_fd_sc_hd__o211a_1
X_12223_ net1298 VGND VGND VPWR VPWR _07779_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12154_ mapped_spi_ram.cmd_addr\[13\] _07079_ _07724_ VGND VGND VPWR VPWR _07731_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11105_ mapped_spi_flash.rcv_bitcount\[5\] _07128_ VGND VGND VPWR VPWR _07129_ sky130_fd_sc_hd__or2_2
X_16962_ CPU.registerFile\[8\]\[23\] _04505_ _04506_ _04665_ VGND VGND VPWR VPWR _04666_
+ sky130_fd_sc_hd__o211a_1
X_12085_ _07682_ VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18701_ net490 _02225_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[1\] sky130_fd_sc_hd__dfxtp_1
X_11036_ net1512 _07054_ _07075_ _07069_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__o211a_1
X_16893_ CPU.registerFile\[2\]\[21\] CPU.registerFile\[3\]\[21\] _04431_ VGND VGND
+ VPWR VPWR _04599_ sky130_fd_sc_hd__mux2_1
X_17418__40 clknet_1_0__leaf__05014_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__inv_2
X_15844_ clknet_1_0__leaf__03654_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__buf_1
X_18632_ clknet_leaf_17_clk _02156_ VGND VGND VPWR VPWR CPU.mem_wdata\[4\] sky130_fd_sc_hd__dfxtp_2
X_18563_ net384 _02087_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_15775_ clknet_1_0__leaf__03654_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__buf_1
X_12987_ net1912 _07341_ _08192_ VGND VGND VPWR VPWR _08197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17514_ _05075_ _05025_ _06135_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__o21bai_1
X_14726_ _05876_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__clkbuf_4
X_18494_ net315 _02018_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_11938_ _06599_ net2127 _07598_ VGND VGND VPWR VPWR _07600_ sky130_fd_sc_hd__mux2_1
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13294__796 clknet_1_0__leaf__08361_ VGND VGND VPWR VPWR net852 sky130_fd_sc_hd__inv_2
X_17445_ _05022_ _06444_ _08256_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__o21ai_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14657_ _02729_ _02730_ _08695_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__mux2_1
X_11869_ _07563_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17376_ per_uart.uart0.rxd_reg\[6\] _04992_ _04993_ per_uart.uart0.rxd_reg\[5\] VGND
+ VGND VPWR VPWR _05003_ sky130_fd_sc_hd__a22o_1
X_14588_ CPU.registerFile\[0\]\[6\] _08706_ _08827_ _08588_ VGND VGND VPWR VPWR _08828_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19115_ net98 _02635_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_13800__1163 clknet_1_1__leaf__08465_ VGND VGND VPWR VPWR net1219 sky130_fd_sc_hd__inv_2
X_16327_ CPU.registerFile\[19\]\[7\] CPU.registerFile\[18\]\[7\] _03923_ VGND VGND
+ VPWR VPWR _04047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19046_ net788 _02566_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_16258_ _03713_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1__f__08472_ clknet_0__08472_ VGND VGND VPWR VPWR clknet_1_1__leaf__08472_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_152_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15209_ _03098_ _03266_ _03269_ _02903_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__a211o_1
X_16189_ CPU.registerFile\[28\]\[4\] CPU.registerFile\[29\]\[4\] _03739_ VGND VGND
+ VPWR VPWR _03912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13604__987 clknet_1_1__leaf__08445_ VGND VGND VPWR VPWR net1043 sky130_fd_sc_hd__inv_2
XFILLER_0_10_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09701_ _05488_ _05898_ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09632_ CPU.PC\[11\] _05942_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09563_ _05373_ _05896_ _05897_ _05906_ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09494_ _05840_ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_867 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13579__964 clknet_1_0__leaf__08443_ VGND VGND VPWR VPWR net1020 sky130_fd_sc_hd__inv_2
X_13722__1093 clknet_1_0__leaf__08457_ VGND VGND VPWR VPWR net1149 sky130_fd_sc_hd__inv_2
X_12910_ _08144_ VGND VGND VPWR VPWR _08156_ sky130_fd_sc_hd__buf_4
XFILLER_0_88_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__08492_ clknet_0__08492_ VGND VGND VPWR VPWR clknet_1_0__leaf__08492_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12841_ _08119_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__clkbuf_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ CPU.registerFile\[30\]\[31\] CPU.registerFile\[31\]\[31\] _03291_ VGND VGND
+ VPWR VPWR _03611_ sky130_fd_sc_hd__mux2_1
X_12772_ _06628_ net2167 _08076_ VGND VGND VPWR VPWR _08082_ sky130_fd_sc_hd__mux2_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ CPU.registerFile\[19\]\[5\] CPU.registerFile\[18\]\[5\] _06064_ VGND VGND
+ VPWR VPWR _08752_ sky130_fd_sc_hd__mux2_1
X_11723_ net2417 _07372_ _07475_ VGND VGND VPWR VPWR _07485_ sky130_fd_sc_hd__mux2_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ CPU.registerFile\[24\]\[29\] _08582_ _03543_ _08540_ VGND VGND VPWR VPWR
+ _03544_ sky130_fd_sc_hd__o211a_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ CPU.registerFile\[28\]\[30\] CPU.registerFile\[29\]\[30\] _03717_ VGND VGND
+ VPWR VPWR _04927_ sky130_fd_sc_hd__mux2_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ CPU.registerFile\[27\]\[3\] CPU.registerFile\[26\]\[3\] _06063_ VGND VGND
+ VPWR VPWR _08685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11654_ net2345 _07372_ _07438_ VGND VGND VPWR VPWR _07448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17161_ _03726_ _03727_ CPU.registerFile\[25\]\[28\] VGND VGND VPWR VPWR _04860_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10605_ _06769_ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__clkbuf_1
X_14373_ CPU.registerFile\[13\]\[1\] CPU.registerFile\[12\]\[1\] _08560_ VGND VGND
+ VPWR VPWR _08618_ sky130_fd_sc_hd__mux2_1
X_11585_ net1681 _07372_ _07401_ VGND VGND VPWR VPWR _07411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16112_ _03744_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__clkbuf_4
X_17092_ _04479_ _04788_ _04792_ _04446_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__o211a_1
X_10536_ _06732_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16043_ _03748_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__clkbuf_4
X_10467_ _06695_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12206_ _07759_ _07766_ VGND VGND VPWR VPWR _07767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13186_ _08303_ _08304_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__nor2_1
X_10398_ _06507_ VGND VGND VPWR VPWR _06657_ sky130_fd_sc_hd__clkbuf_4
X_12137_ net1408 _07714_ _07719_ _07713_ VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__o211a_1
X_17994_ net1005 _01522_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12068_ _07668_ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__clkbuf_1
X_16945_ _04441_ _04647_ _04649_ _04612_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__a211o_1
X_11019_ CPU.PC\[11\] _07031_ _07058_ _07060_ _05703_ VGND VGND VPWR VPWR _07061_
+ sky130_fd_sc_hd__o221a_1
X_16876_ _04367_ _04578_ _04582_ _04410_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18615_ net436 _02139_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18546_ net367 _02070_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_14149__288 clknet_1_1__leaf__08499_ VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__inv_2
XFILLER_0_47_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14709_ CPU.registerFile\[8\]\[9\] _08776_ _02781_ _08622_ VGND VGND VPWR VPWR _02782_
+ sky130_fd_sc_hd__o211a_1
X_18477_ net298 _02001_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17428_ _08379_ _05017_ _06490_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_56_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17359_ per_uart.uart0.rx_bitcount\[2\] per_uart.uart0.rx_bitcount\[0\] per_uart.uart0.rx_bitcount\[1\]
+ per_uart.uart0.rx_bitcount\[3\] VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_42_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19029_ net771 _02549_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[14\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__08455_ clknet_0__08455_ VGND VGND VPWR VPWR clknet_1_1__leaf__08455_
+ sky130_fd_sc_hd__clkbuf_16
X_15737__528 clknet_1_1__leaf__03651_ VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__inv_2
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08486_ _08486_ VGND VGND VPWR VPWR clknet_0__08486_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08994_ CPU.aluIn1\[17\] _05345_ VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09615_ CPU.PC\[3\] _05958_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__xor2_1
X_09546_ CPU.PC\[16\] CPU.PC\[15\] _05889_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_918 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09477_ _05824_ VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11370_ net1860 _05873_ _07274_ VGND VGND VPWR VPWR _07282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10321_ net1339 VGND VGND VPWR VPWR _06605_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_132_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13040_ CPU.registerFile\[4\]\[24\] _05872_ _08217_ VGND VGND VPWR VPWR _08225_ sky130_fd_sc_hd__mux2_1
X_10252_ _06565_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__clkbuf_1
X_10183_ _06176_ _06497_ _06505_ _05541_ VGND VGND VPWR VPWR _06506_ sky130_fd_sc_hd__a22o_1
X_14991_ CPU.registerFile\[13\]\[16\] CPU.registerFile\[12\]\[16\] _02935_ VGND VGND
+ VPWR VPWR _03057_ sky130_fd_sc_hd__mux2_1
X_13942_ clknet_1_0__leaf__08473_ VGND VGND VPWR VPWR _08479_ sky130_fd_sc_hd__buf_1
X_16730_ _04438_ _04439_ _04279_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__mux2_1
X_16661_ _04361_ _04372_ _04138_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__o21a_1
Xclkbuf_1_0__f__08475_ clknet_0__08475_ VGND VGND VPWR VPWR clknet_1_0__leaf__08475_
+ sky130_fd_sc_hd__clkbuf_16
X_18400_ net221 _01928_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12824_ _05767_ net2282 _08109_ VGND VGND VPWR VPWR _08111_ sky130_fd_sc_hd__mux2_1
X_16592_ _03713_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__clkbuf_4
X_15543_ CPU.registerFile\[2\]\[30\] CPU.registerFile\[3\]\[30\] _03275_ VGND VGND
+ VPWR VPWR _03595_ sky130_fd_sc_hd__mux2_1
X_18331_ net152 _01859_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ _06611_ net2223 _08065_ VGND VGND VPWR VPWR _08073_ sky130_fd_sc_hd__mux2_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _07476_ VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__clkbuf_1
X_18262_ net1273 _01790_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15474_ _03230_ _03523_ _03527_ _05876_ VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12686_ _08036_ VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__clkbuf_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17213_ CPU.registerFile\[9\]\[30\] _03709_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__or2_1
X_14425_ CPU.registerFile\[0\]\[2\] _08584_ _08668_ _08588_ VGND VGND VPWR VPWR _08669_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11637_ _07439_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__clkbuf_1
X_18193_ net1204 _01721_ VGND VGND VPWR VPWR mapped_spi_ram.snd_bitcount\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13940__100 clknet_1_0__leaf__08478_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__inv_2
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17144_ CPU.registerFile\[15\]\[28\] CPU.registerFile\[14\]\[28\] _04550_ VGND VGND
+ VPWR VPWR _04843_ sky130_fd_sc_hd__mux2_1
X_14356_ CPU.registerFile\[16\]\[1\] _08412_ _08600_ _06037_ VGND VGND VPWR VPWR _08601_
+ sky130_fd_sc_hd__o211a_1
X_11568_ _07402_ VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold708 CPU.registerFile\[13\]\[24\] VGND VGND VPWR VPWR net2005 sky130_fd_sc_hd__dlygate4sd3_1
X_17075_ _04419_ _04773_ _04775_ _03716_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__a211o_1
Xhold719 CPU.registerFile\[22\]\[14\] VGND VGND VPWR VPWR net2016 sky130_fd_sc_hd__dlygate4sd3_1
X_10519_ _06723_ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14287_ _08532_ VGND VGND VPWR VPWR _08533_ sky130_fd_sc_hd__clkbuf_4
X_11499_ _06385_ VGND VGND VPWR VPWR _07362_ sky130_fd_sc_hd__buf_4
Xclkbuf_0__08340_ _08340_ VGND VGND VPWR VPWR clknet_0__08340_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16026_ CPU.registerFile\[24\]\[0\] _08393_ _03747_ _03752_ VGND VGND VPWR VPWR _03753_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13169_ _08293_ net1561 VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17977_ net988 _01505_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_16928_ CPU.registerFile\[6\]\[22\] CPU.registerFile\[7\]\[22\] _04426_ VGND VGND
+ VPWR VPWR _04633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16859_ CPU.registerFile\[28\]\[20\] CPU.registerFile\[29\]\[20\] _04526_ VGND VGND
+ VPWR VPWR _04566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09400_ _05253_ _05533_ _05536_ CPU.aluReg\[30\] VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09331_ _05682_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__buf_8
X_14082__228 clknet_1_0__leaf__08492_ VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__inv_2
X_18529_ net350 _02053_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09262_ CPU.aluIn1\[14\] _05543_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_910 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09193_ _05544_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__buf_4
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13721__1092 clknet_1_0__leaf__08457_ VGND VGND VPWR VPWR net1148 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__08507_ clknet_0__08507_ VGND VGND VPWR VPWR clknet_1_1__leaf__08507_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_114_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08438_ clknet_0__08438_ VGND VGND VPWR VPWR clknet_1_1__leaf__08438_
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0__08469_ _08469_ VGND VGND VPWR VPWR clknet_0__08469_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__08369_ clknet_0__08369_ VGND VGND VPWR VPWR clknet_1_1__leaf__08369_
+ sky130_fd_sc_hd__clkbuf_16
X_13888__52 clknet_1_0__leaf__08474_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__inv_2
Xhold13 mapped_spi_ram.rcv_bitcount\[3\] VGND VGND VPWR VPWR net1310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 _07827_ VGND VGND VPWR VPWR net1321 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ _05328_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__inv_2
Xhold35 _06336_ VGND VGND VPWR VPWR net1332 sky130_fd_sc_hd__clkbuf_2
Xhold46 mapped_spi_ram.cmd_addr\[3\] VGND VGND VPWR VPWR net1343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 _08241_ VGND VGND VPWR VPWR net1354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 mapped_spi_ram.cmd_addr\[30\] VGND VGND VPWR VPWR net1365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 _06398_ VGND VGND VPWR VPWR net1376 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10870_ _06942_ VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09529_ net2031 _05873_ _05742_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__mux2_1
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12540_ _07959_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12471_ _07922_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11422_ _05733_ VGND VGND VPWR VPWR _07309_ sky130_fd_sc_hd__buf_4
X_15190_ CPU.registerFile\[20\]\[21\] _03080_ _03250_ _03082_ VGND VGND VPWR VPWR
+ _03251_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11353_ _07272_ VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10304_ _06592_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11284_ _07235_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13023_ _08215_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__clkbuf_1
X_17900_ clknet_leaf_22_clk _01428_ VGND VGND VPWR VPWR CPU.Bimm\[11\] sky130_fd_sc_hd__dfxtp_2
X_10235_ net2258 _06555_ net15 VGND VGND VPWR VPWR _06556_ sky130_fd_sc_hd__mux2_1
X_18880_ net654 _02400_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_17831_ net911 _01393_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_10166_ _05956_ _05955_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__and2b_1
X_17762_ net842 _01324_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_10097_ _05964_ _05949_ VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__or2b_1
X_14974_ CPU.registerFile\[22\]\[16\] CPU.registerFile\[23\]\[16\] _02998_ VGND VGND
+ VPWR VPWR _03040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16713_ CPU.registerFile\[13\]\[17\] _04380_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17693_ _05207_ _05219_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__and2_1
XFILLER_0_159_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16644_ _04354_ _04355_ _04279_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__08458_ clknet_0__08458_ VGND VGND VPWR VPWR clknet_1_0__leaf__08458_
+ sky130_fd_sc_hd__clkbuf_16
X_12807_ CPU.aluShamt\[4\] _06859_ VGND VGND VPWR VPWR _08100_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13787_ clknet_1_0__leaf__08462_ VGND VGND VPWR VPWR _08464_ sky130_fd_sc_hd__buf_1
X_16575_ _04286_ _04288_ _03961_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__mux2_1
X_10999_ _05606_ _07042_ _05609_ VGND VGND VPWR VPWR _07043_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18314_ net135 _01842_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15526_ CPU.registerFile\[27\]\[30\] CPU.registerFile\[26\]\[30\] _08576_ VGND VGND
+ VPWR VPWR _03578_ sky130_fd_sc_hd__mux2_1
X_12738_ _08063_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18245_ net1256 _01773_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_15457_ _06013_ _03506_ _03510_ _08422_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__o211a_1
Xclkbuf_0__04983_ _04983_ VGND VGND VPWR VPWR clknet_0__04983_ sky130_fd_sc_hd__clkbuf_16
X_12669_ _06661_ net2115 _07992_ VGND VGND VPWR VPWR _08027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14408_ _08543_ _08649_ _08651_ _08552_ VGND VGND VPWR VPWR _08652_ sky130_fd_sc_hd__a211o_1
X_15388_ CPU.registerFile\[13\]\[26\] CPU.registerFile\[12\]\[26\] _08794_ VGND VGND
+ VPWR VPWR _03444_ sky130_fd_sc_hd__mux2_1
X_18176_ net1187 _01704_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14339_ _08566_ VGND VGND VPWR VPWR _08585_ sky130_fd_sc_hd__clkbuf_4
X_17127_ _03722_ _04824_ _04826_ _04612_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__a211o_1
XFILLER_0_123_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold505 CPU.registerFile\[11\]\[10\] VGND VGND VPWR VPWR net1802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 CPU.registerFile\[18\]\[20\] VGND VGND VPWR VPWR net1813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 CPU.registerFile\[10\]\[26\] VGND VGND VPWR VPWR net1824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 CPU.registerFile\[5\]\[27\] VGND VGND VPWR VPWR net1835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17058_ CPU.registerFile\[20\]\[25\] CPU.registerFile\[21\]\[25\] _03737_ VGND VGND
+ VPWR VPWR _04760_ sky130_fd_sc_hd__mux2_1
Xhold549 CPU.registerFile\[6\]\[12\] VGND VGND VPWR VPWR net1846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16009_ _06171_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__clkbuf_4
X_08900_ CPU.rs2\[30\] _05247_ _05251_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__o21a_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _05427_ _06212_ _06214_ _05800_ VGND VGND VPWR VPWR _06215_ sky130_fd_sc_hd__a211o_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1205 CPU.registerFile\[25\]\[29\] VGND VGND VPWR VPWR net2502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 CPU.registerFile\[31\]\[16\] VGND VGND VPWR VPWR net2513 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 CPU.registerFile\[25\]\[27\] VGND VGND VPWR VPWR net2524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1238 CPU.registerFile\[8\]\[15\] VGND VGND VPWR VPWR net2535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 CPU.registerFile\[25\]\[11\] VGND VGND VPWR VPWR net2546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18576__33 VGND VGND VPWR VPWR _18576__33/HI net33 sky130_fd_sc_hd__conb_1
XFILLER_0_88_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13947__106 clknet_1_0__leaf__08479_ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__inv_2
X_09314_ _05664_ _05665_ _05636_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09245_ CPU.aluIn1\[10\] CPU.Bimm\[10\] VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15895__638 clknet_1_0__leaf__03684_ VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__inv_2
X_09176_ _05526_ _05527_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__nor2_2
XFILLER_0_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13993__148 clknet_1_1__leaf__08483_ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__inv_2
X_10020_ _06126_ _06345_ _06348_ _05818_ VGND VGND VPWR VPWR _06349_ sky130_fd_sc_hd__o211a_1
X_11971_ _06632_ net2116 _07609_ VGND VGND VPWR VPWR _07617_ sky130_fd_sc_hd__mux2_1
X_10922_ mapped_spi_flash.state\[1\] _06981_ VGND VGND VPWR VPWR _06984_ sky130_fd_sc_hd__and2_1
X_14690_ CPU.registerFile\[20\]\[9\] _08839_ _02762_ _08841_ VGND VGND VPWR VPWR _02763_
+ sky130_fd_sc_hd__o211a_1
X_13741__1111 clknet_1_0__leaf__08458_ VGND VGND VPWR VPWR net1167 sky130_fd_sc_hd__inv_2
XFILLER_0_39_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14065__212 clknet_1_0__leaf__08491_ VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__inv_2
X_10853_ _06929_ VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16360_ CPU.registerFile\[27\]\[8\] CPU.registerFile\[26\]\[8\] _03837_ VGND VGND
+ VPWR VPWR _04079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10784_ CPU.aluReg\[30\] CPU.aluReg\[28\] _06872_ VGND VGND VPWR VPWR _06876_ sky130_fd_sc_hd__mux2_1
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15311_ _03006_ _03366_ _03368_ _03218_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__a211o_1
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12523_ _07949_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__clkbuf_1
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16291_ CPU.registerFile\[10\]\[7\] CPU.registerFile\[11\]\[7\] _03931_ VGND VGND
+ VPWR VPWR _04011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_915 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18030_ net1041 _01558_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_15242_ CPU.registerFile\[13\]\[22\] CPU.registerFile\[12\]\[22\] _02935_ VGND VGND
+ VPWR VPWR _03302_ sky130_fd_sc_hd__mux2_1
X_12454_ net1756 _07366_ _07906_ VGND VGND VPWR VPWR _07913_ sky130_fd_sc_hd__mux2_1
X_11405_ _07300_ VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__clkbuf_1
X_15173_ _08566_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_62_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12385_ _07876_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__03650_ _03650_ VGND VGND VPWR VPWR clknet_0__03650_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_22_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11336_ net2663 _06361_ _07260_ VGND VGND VPWR VPWR _07264_ sky130_fd_sc_hd__mux2_1
X_18932_ net706 _02452_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_11267_ _06645_ net2022 _07223_ VGND VGND VPWR VPWR _07227_ sky130_fd_sc_hd__mux2_1
X_13006_ net2084 _07360_ _08203_ VGND VGND VPWR VPWR _08207_ sky130_fd_sc_hd__mux2_1
X_10218_ _05724_ _06537_ _06538_ _06391_ VGND VGND VPWR VPWR _06539_ sky130_fd_sc_hd__a211o_1
X_18863_ net637 _02383_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_11198_ _07183_ _07184_ _07186_ _00004_ VGND VGND VPWR VPWR _07188_ sky130_fd_sc_hd__a211o_2
X_17814_ net894 _01376_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_10149_ _05691_ _06287_ VGND VGND VPWR VPWR _06473_ sky130_fd_sc_hd__or2_1
X_18794_ net583 _02318_ VGND VGND VPWR VPWR CPU.aluReg\[24\] sky130_fd_sc_hd__dfxtp_1
X_13301__802 clknet_1_0__leaf__08362_ VGND VGND VPWR VPWR net858 sky130_fd_sc_hd__inv_2
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17745_ net830 _01311_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_14957_ CPU.registerFile\[5\]\[15\] CPU.registerFile\[4\]\[15\] _08864_ VGND VGND
+ VPWR VPWR _03024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17676_ _05206_ VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14888_ CPU.registerFile\[17\]\[14\] _08795_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__or2_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16627_ _04099_ _04336_ _04338_ _04105_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__a211o_1
X_13258__778 clknet_1_1__leaf__08344_ VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__inv_2
XFILLER_0_134_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13490__884 clknet_1_1__leaf__08434_ VGND VGND VPWR VPWR net940 sky130_fd_sc_hd__inv_2
X_16558_ _03985_ _03986_ CPU.registerFile\[1\]\[13\] VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15509_ _08414_ _03559_ _03561_ _08419_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__a211o_1
XFILLER_0_155_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16489_ CPU.registerFile\[27\]\[11\] CPU.registerFile\[26\]\[11\] _03837_ VGND VGND
+ VPWR VPWR _04205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09030_ _05373_ _05376_ _05372_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__a21oi_2
X_18228_ net1239 _01756_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[29\] sky130_fd_sc_hd__dfxtp_1
X_15820__570 clknet_1_0__leaf__03656_ VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__inv_2
XFILLER_0_13_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14194__329 clknet_1_0__leaf__08503_ VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__inv_2
X_18159_ net1170 _01687_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_bitcount\[5\] sky130_fd_sc_hd__dfxtp_1
Xhold302 mapped_spi_flash.rcv_data\[17\] VGND VGND VPWR VPWR net1599 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold313 per_uart.uart0.enable16_counter\[8\] VGND VGND VPWR VPWR net1610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold324 CPU.cycles\[13\] VGND VGND VPWR VPWR net1621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 _02697_ VGND VGND VPWR VPWR net1632 sky130_fd_sc_hd__dlygate4sd3_1
X_13663__1041 clknet_1_1__leaf__08450_ VGND VGND VPWR VPWR net1097 sky130_fd_sc_hd__inv_2
Xhold346 mapped_spi_flash.rcv_data\[6\] VGND VGND VPWR VPWR net1643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 _02326_ VGND VGND VPWR VPWR net1654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09932_ _05911_ _06263_ _06264_ _06197_ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold368 CPU.rs2\[12\] VGND VGND VPWR VPWR net1665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 CPU.registerFile\[6\]\[30\] VGND VGND VPWR VPWR net1676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03679_ clknet_0__03679_ VGND VGND VPWR VPWR clknet_1_1__leaf__03679_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ _06178_ _06179_ _06194_ _06198_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__or4b_4
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 CPU.registerFile\[11\]\[5\] VGND VGND VPWR VPWR net2299 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 CPU.registerFile\[26\]\[28\] VGND VGND VPWR VPWR net2310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 CPU.registerFile\[13\]\[1\] VGND VGND VPWR VPWR net2321 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _05346_ _05523_ _05749_ VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__o21ai_1
Xhold1035 CPU.registerFile\[29\]\[19\] VGND VGND VPWR VPWR net2332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1046 CPU.registerFile\[10\]\[13\] VGND VGND VPWR VPWR net2343 sky130_fd_sc_hd__dlygate4sd3_1
X_14014__166 clknet_1_0__leaf__08486_ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__inv_2
Xhold1057 CPU.registerFile\[31\]\[8\] VGND VGND VPWR VPWR net2354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1068 CPU.registerFile\[16\]\[15\] VGND VGND VPWR VPWR net2365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 CPU.registerFile\[30\]\[4\] VGND VGND VPWR VPWR net2376 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13573__959 clknet_1_1__leaf__08442_ VGND VGND VPWR VPWR net1015 sky130_fd_sc_hd__inv_2
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15903__645 clknet_1_0__leaf__03685_ VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__inv_2
XFILLER_0_76_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09228_ CPU.aluIn1\[1\] _05578_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15602__406 clknet_1_0__leaf__03638_ VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__inv_2
XFILLER_0_91_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09159_ _05252_ CPU.aluIn1\[30\] VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__and2b_1
XFILLER_0_161_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12170_ _07739_ _07742_ VGND VGND VPWR VPWR _07743_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11121_ net1438 _07135_ VGND VGND VPWR VPWR _07141_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold880 CPU.registerFile\[8\]\[17\] VGND VGND VPWR VPWR net2177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 CPU.registerFile\[22\]\[4\] VGND VGND VPWR VPWR net2188 sky130_fd_sc_hd__dlygate4sd3_1
X_11052_ _05570_ _05592_ VGND VGND VPWR VPWR _07089_ sky130_fd_sc_hd__and2_1
X_10003_ net1599 _05698_ _05717_ per_uart.tx_busy _06332_ VGND VGND VPWR VPWR _06333_
+ sky130_fd_sc_hd__a221o_1
X_14811_ CPU.registerFile\[16\]\[12\] _02755_ _02880_ _02757_ VGND VGND VPWR VPWR
+ _02881_ sky130_fd_sc_hd__o211a_1
X_15791_ _03663_ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17530_ _05100_ _05101_ _05058_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__a21oi_1
X_14742_ _06396_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__clkbuf_4
X_11954_ _06615_ net2274 _07598_ VGND VGND VPWR VPWR _07608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10905_ CPU.aluReg\[1\] _06968_ _06868_ VGND VGND VPWR VPWR _06969_ sky130_fd_sc_hd__mux2_1
X_14673_ _08574_ _02741_ _02745_ _02746_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__o211a_1
X_17461_ _08379_ _05017_ _06355_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_39_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11885_ _07571_ VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16412_ CPU.registerFile\[22\]\[9\] CPU.registerFile\[23\]\[9\] _03958_ VGND VGND
+ VPWR VPWR _04130_ sky130_fd_sc_hd__mux2_1
X_10836_ _06916_ VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19131_ clknet_leaf_10_clk _02651_ VGND VGND VPWR VPWR CPU.PC\[13\] sky130_fd_sc_hd__dfxtp_2
X_16343_ CPU.registerFile\[12\]\[8\] _04017_ _04018_ _04061_ VGND VGND VPWR VPWR _04062_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10767_ _06860_ VGND VGND VPWR VPWR _06861_ sky130_fd_sc_hd__buf_4
X_15878__622 clknet_1_1__leaf__03683_ VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__inv_2
X_12506_ _07940_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16274_ CPU.registerFile\[27\]\[6\] CPU.registerFile\[26\]\[6\] _03837_ VGND VGND
+ VPWR VPWR _03995_ sky130_fd_sc_hd__mux2_1
X_19062_ net804 _02582_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10698_ _06821_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18013_ net1024 _01541_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_15225_ CPU.registerFile\[16\]\[22\] _03159_ _03284_ _03161_ VGND VGND VPWR VPWR
+ _03285_ sky130_fd_sc_hd__o211a_1
X_12437_ net2343 _07349_ _07895_ VGND VGND VPWR VPWR _07904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15156_ _06396_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__clkbuf_4
X_12368_ _07867_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13976__132 clknet_1_1__leaf__08482_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__inv_2
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11319_ net2412 _06169_ _07249_ VGND VGND VPWR VPWR _07255_ sky130_fd_sc_hd__mux2_1
X_15087_ _05875_ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__clkbuf_4
X_12299_ mapped_spi_ram.rcv_data\[1\] _07786_ VGND VGND VPWR VPWR _07825_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18915_ net689 _02435_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_13299__801 clknet_1_1__leaf__08361_ VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__inv_2
X_18846_ clknet_leaf_7_clk _02370_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_18777_ net566 _02301_ VGND VGND VPWR VPWR CPU.aluReg\[7\] sky130_fd_sc_hd__dfxtp_1
X_15989_ _03713_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17728_ net813 _01294_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17659_ per_uart.uart0.rx_busy _04988_ _05185_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_148_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14202__336 clknet_1_0__leaf__08504_ VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__inv_2
XFILLER_0_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09013_ _05363_ _05364_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold110 _08238_ VGND VGND VPWR VPWR net1407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold121 _08236_ VGND VGND VPWR VPWR net1418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 mapped_spi_ram.rcv_data\[26\] VGND VGND VPWR VPWR net1429 sky130_fd_sc_hd__dlygate4sd3_1
X_13619__1001 clknet_1_1__leaf__08446_ VGND VGND VPWR VPWR net1057 sky130_fd_sc_hd__inv_2
XFILLER_0_79_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold143 _08248_ VGND VGND VPWR VPWR net1440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13740__1110 clknet_1_0__leaf__08458_ VGND VGND VPWR VPWR net1166 sky130_fd_sc_hd__inv_2
Xhold154 per_uart.uart0.txd_reg\[0\] VGND VGND VPWR VPWR net1451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 mapped_spi_ram.cmd_addr\[9\] VGND VGND VPWR VPWR net1462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold176 mapped_spi_ram.rcv_data\[4\] VGND VGND VPWR VPWR net1473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 mapped_spi_ram.rcv_data\[2\] VGND VGND VPWR VPWR net1484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 mapped_spi_ram.cmd_addr\[16\] VGND VGND VPWR VPWR net1495 sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ CPU.Jimm\[13\] _06203_ _05788_ _06204_ _06247_ VGND VGND VPWR VPWR _06248_
+ sky130_fd_sc_hd__o32a_1
X_09846_ CPU.aluIn1\[12\] _05317_ VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__nand2_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _05355_ _05747_ VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__nor2_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827__576 clknet_1_1__leaf__03678_ VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__inv_2
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13883__1239 clknet_1_1__leaf__08472_ VGND VGND VPWR VPWR net1295 sky130_fd_sc_hd__inv_2
X_11670_ _07457_ VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ _06779_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10552_ net1855 _05786_ _06739_ VGND VGND VPWR VPWR _06742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14177__313 clknet_1_0__leaf__08502_ VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__inv_2
X_13271_ net1596 _08351_ VGND VGND VPWR VPWR _08352_ sky130_fd_sc_hd__or2_1
X_10483_ net2255 _05786_ _06702_ VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__mux2_1
X_15010_ CPU.registerFile\[17\]\[17\] _03036_ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__or2_1
X_12222_ net1324 _07764_ _07776_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12153_ net1472 _07714_ _07730_ _07713_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11104_ mapped_spi_flash.rcv_bitcount\[4\] _07127_ VGND VGND VPWR VPWR _07128_ sky130_fd_sc_hd__or2_1
X_16961_ CPU.registerFile\[9\]\[23\] _04460_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__or2_1
X_12084_ _06992_ _07681_ VGND VGND VPWR VPWR _07682_ sky130_fd_sc_hd__and2_1
X_18700_ net489 _02224_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[0\] sky130_fd_sc_hd__dfxtp_1
X_11035_ _07048_ _07074_ VGND VGND VPWR VPWR _07075_ sky130_fd_sc_hd__or2_1
X_16892_ _04596_ _04597_ _04557_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__mux2_1
X_18631_ clknet_leaf_24_clk _02155_ VGND VGND VPWR VPWR CPU.mem_wdata\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_99_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13556__943 clknet_1_1__leaf__08441_ VGND VGND VPWR VPWR net999 sky130_fd_sc_hd__inv_2
X_18562_ net383 _02086_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_12986_ _08196_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17513_ _08311_ _06137_ _08331_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__or3_1
XFILLER_0_115_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14725_ _08513_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__buf_2
X_18493_ net314 _02017_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_13662__1040 clknet_1_1__leaf__08450_ VGND VGND VPWR VPWR net1096 sky130_fd_sc_hd__inv_2
X_11937_ _07599_ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _05030_ _05031_ _05020_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__a21oi_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14656_ CPU.registerFile\[13\]\[8\] CPU.registerFile\[12\]\[8\] _08693_ VGND VGND
+ VPWR VPWR _02730_ sky130_fd_sc_hd__mux2_1
X_11868_ _06593_ net2008 _07562_ VGND VGND VPWR VPWR _07563_ sky130_fd_sc_hd__mux2_1
X_10819_ CPU.aluReg\[22\] CPU.aluReg\[20\] _06872_ VGND VGND VPWR VPWR _06903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17375_ _05002_ VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__clkbuf_1
X_11799_ _07525_ VGND VGND VPWR VPWR _07526_ sky130_fd_sc_hd__buf_4
X_14587_ _08585_ _08586_ CPU.registerFile\[1\]\[6\] VGND VGND VPWR VPWR _08827_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19114_ net97 _02634_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_16326_ _04044_ _04045_ _03961_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14043__192 clknet_1_1__leaf__08489_ VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__inv_2
X_19045_ net787 _02565_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16257_ CPU.registerFile\[12\]\[6\] _03707_ _03708_ _03977_ VGND VGND VPWR VPWR _03978_
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_1__f__08471_ clknet_0__08471_ VGND VGND VPWR VPWR clknet_1_1__leaf__08471_
+ sky130_fd_sc_hd__clkbuf_16
X_13469_ CPU.Iimm\[4\] _08425_ _08416_ VGND VGND VPWR VPWR _08426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15208_ CPU.registerFile\[8\]\[21\] _03018_ _03267_ _03268_ VGND VGND VPWR VPWR _03269_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_871 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16188_ CPU.registerFile\[30\]\[4\] CPU.registerFile\[31\]\[4\] _03796_ VGND VGND
+ VPWR VPWR _03911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15139_ _08513_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__buf_2
XFILLER_0_49_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15932__671 clknet_1_0__leaf__03688_ VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__inv_2
X_09700_ _05488_ _06041_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09631_ _05944_ _05973_ _05974_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15631__432 clknet_1_0__leaf__03641_ VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__inv_2
X_18829_ net618 _02353_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_13496__890 clknet_1_0__leaf__08434_ VGND VGND VPWR VPWR net946 sky130_fd_sc_hd__inv_2
X_09562_ _05424_ _05901_ _05905_ _05516_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09493_ net2347 _05839_ _05742_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14126__267 clknet_1_0__leaf__08497_ VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__inv_2
XFILLER_0_148_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15714__507 clknet_1_1__leaf__03649_ VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__inv_2
X_09829_ _05881_ _06156_ _06165_ _05744_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_1_0__f__08491_ clknet_0__08491_ VGND VGND VPWR VPWR clknet_1_0__leaf__08491_
+ sky130_fd_sc_hd__clkbuf_16
X_12840_ _06032_ net2481 _08109_ VGND VGND VPWR VPWR _08119_ sky130_fd_sc_hd__mux2_1
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15909__651 clknet_1_1__leaf__03685_ VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__inv_2
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _08081_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__clkbuf_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11722_ _07484_ VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__clkbuf_1
X_14510_ CPU.mem_wdata\[4\] _08514_ _08750_ _08751_ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__o211a_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15490_ _08566_ _08568_ CPU.registerFile\[25\]\[29\] VGND VGND VPWR VPWR _03543_
+ sky130_fd_sc_hd__a21o_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _07447_ VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__clkbuf_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ _08682_ _08683_ _08609_ VGND VGND VPWR VPWR _08684_ sky130_fd_sc_hd__mux2_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760__549 clknet_1_1__leaf__03653_ VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__inv_2
XFILLER_0_154_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10604_ net1963 _06465_ _06761_ VGND VGND VPWR VPWR _06769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14372_ CPU.registerFile\[15\]\[1\] CPU.registerFile\[14\]\[1\] _08558_ VGND VGND
+ VPWR VPWR _08617_ sky130_fd_sc_hd__mux2_1
X_17160_ CPU.registerFile\[27\]\[28\] CPU.registerFile\[26\]\[28\] _04646_ VGND VGND
+ VPWR VPWR _04859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11584_ _07410_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16111_ _03834_ _03835_ _03742_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10535_ net1970 _06465_ _06724_ VGND VGND VPWR VPWR _06732_ sky130_fd_sc_hd__mux2_1
X_17091_ _04441_ _04789_ _04791_ _04612_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__a211o_1
XFILLER_0_101_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16042_ _06534_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__buf_4
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10466_ _06653_ net2271 _06687_ VGND VGND VPWR VPWR _06695_ sky130_fd_sc_hd__mux2_1
X_17294__710 clknet_1_0__leaf__04979_ VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__inv_2
XFILLER_0_32_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12205_ mapped_spi_ram.snd_bitcount\[4\] _07758_ VGND VGND VPWR VPWR _07766_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13185_ net1562 _08301_ VGND VGND VPWR VPWR _08304_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10397_ _06656_ VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12136_ _07715_ _07718_ VGND VGND VPWR VPWR _07719_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17993_ net1004 _01521_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_12067_ net1664 _07374_ _07634_ VGND VGND VPWR VPWR _07668_ sky130_fd_sc_hd__mux2_1
X_16944_ CPU.registerFile\[24\]\[22\] _04319_ _04569_ _04648_ VGND VGND VPWR VPWR
+ _04649_ sky130_fd_sc_hd__o211a_1
X_11018_ _07031_ _07059_ VGND VGND VPWR VPWR _07060_ sky130_fd_sc_hd__nand2_1
X_16875_ CPU.registerFile\[16\]\[20\] _04252_ _04494_ _04581_ VGND VGND VPWR VPWR
+ _04582_ sky130_fd_sc_hd__o211a_1
X_18614_ net435 _02138_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18545_ net366 _02069_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_12969_ _08187_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__clkbuf_1
X_13618__1000 clknet_1_1__leaf__08446_ VGND VGND VPWR VPWR net1056 sky130_fd_sc_hd__inv_2
XFILLER_0_157_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14708_ _02733_ _02734_ CPU.registerFile\[9\]\[9\] VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__a21o_1
X_18476_ net297 _02000_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17427_ _08330_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__buf_2
XFILLER_0_118_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14639_ CPU.registerFile\[16\]\[8\] _08412_ _08876_ _06037_ VGND VGND VPWR VPWR _08877_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17358_ _04986_ _04988_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13610__992 clknet_1_0__leaf__08446_ VGND VGND VPWR VPWR net1048 sky130_fd_sc_hd__inv_2
XFILLER_0_42_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16309_ _03985_ _03986_ CPU.registerFile\[1\]\[7\] VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19028_ net770 _02548_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[13\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__08454_ clknet_0__08454_ VGND VGND VPWR VPWR clknet_1_1__leaf__08454_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08485_ _08485_ VGND VGND VPWR VPWR clknet_0__08485_ sky130_fd_sc_hd__clkbuf_16
X_13383__876 clknet_1_1__leaf__08370_ VGND VGND VPWR VPWR net932 sky130_fd_sc_hd__inv_2
X_13882__1238 clknet_1_1__leaf__08472_ VGND VGND VPWR VPWR net1294 sky130_fd_sc_hd__inv_2
X_08993_ CPU.rs2\[17\] _05246_ _05250_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09614_ CPU.Iimm\[3\] CPU.instr\[3\] _05922_ _05737_ VGND VGND VPWR VPWR _05958_
+ sky130_fd_sc_hd__a22o_1
X_09545_ CPU.PC\[14\] _05888_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09476_ _05745_ _05820_ _05821_ _05823_ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__a211o_2
XFILLER_0_19_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_871 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15939__677 clknet_1_1__leaf__03689_ VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__inv_2
X_10320_ _06604_ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10251_ net1685 _05853_ _06558_ VGND VGND VPWR VPWR _06565_ sky130_fd_sc_hd__mux2_1
X_10182_ _05282_ _05769_ _05536_ net1421 _06504_ VGND VGND VPWR VPWR _06505_ sky130_fd_sc_hd__a221o_2
X_14990_ CPU.registerFile\[15\]\[16\] CPU.registerFile\[14\]\[16\] _03013_ VGND VGND
+ VPWR VPWR _03056_ sky130_fd_sc_hd__mux2_1
X_16660_ _04170_ _04366_ _04371_ _04180_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__08474_ clknet_0__08474_ VGND VGND VPWR VPWR clknet_1_0__leaf__08474_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12823_ _08110_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__clkbuf_1
X_16591_ _04015_ _04301_ _04303_ _03979_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18330_ net151 _01858_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_15542_ _03592_ _03593_ _08562_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__mux2_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _08072_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__clkbuf_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17326__739 clknet_1_1__leaf__04982_ VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__inv_2
XFILLER_0_56_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ net2287 _07353_ _07475_ VGND VGND VPWR VPWR _07476_ sky130_fd_sc_hd__mux2_1
X_18261_ net1272 _01789_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _06609_ net2616 _08029_ VGND VGND VPWR VPWR _08036_ sky130_fd_sc_hd__mux2_1
X_15473_ _08414_ _03524_ _03526_ _08419_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__a211o_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ CPU.registerFile\[10\]\[30\] CPU.registerFile\[11\]\[30\] _06173_ VGND VGND
+ VPWR VPWR _04909_ sky130_fd_sc_hd__mux2_1
X_11636_ net2370 _07353_ _07438_ VGND VGND VPWR VPWR _07439_ sky130_fd_sc_hd__mux2_1
X_14424_ _08585_ _08586_ CPU.registerFile\[1\]\[2\] VGND VGND VPWR VPWR _08668_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18192_ net1203 net1428 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17143_ _04503_ _04839_ _04841_ _04509_ VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__a211o_1
X_11567_ net1716 _07353_ _07401_ VGND VGND VPWR VPWR _07402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14355_ CPU.registerFile\[17\]\[1\] _06456_ VGND VGND VPWR VPWR _08600_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10518_ net2017 _06267_ _06713_ VGND VGND VPWR VPWR _06723_ sky130_fd_sc_hd__mux2_1
X_17074_ CPU.registerFile\[12\]\[26\] _04421_ _04422_ _04774_ VGND VGND VPWR VPWR
+ _04775_ sky130_fd_sc_hd__o211a_1
Xhold709 CPU.registerFile\[10\]\[14\] VGND VGND VPWR VPWR net2006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14286_ _06012_ VGND VGND VPWR VPWR _08532_ sky130_fd_sc_hd__buf_4
X_11498_ _07361_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__clkbuf_1
X_16025_ _03749_ _03751_ CPU.registerFile\[25\]\[0\] VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__a21o_1
X_10449_ _06636_ net2126 _06676_ VGND VGND VPWR VPWR _06686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13168_ CPU.cycles\[19\] _08291_ net1560 VGND VGND VPWR VPWR _08294_ sky130_fd_sc_hd__a21oi_1
X_14155__293 clknet_1_0__leaf__08500_ VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__inv_2
X_12119_ net1312 _07671_ VGND VGND VPWR VPWR _07706_ sky130_fd_sc_hd__nor2_4
X_13099_ net1301 _07675_ _06856_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__o21a_1
X_17976_ net987 _01504_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_16927_ _04419_ _04629_ _04631_ _04383_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16858_ CPU.registerFile\[30\]\[20\] CPU.registerFile\[31\]\[20\] _04201_ VGND VGND
+ VPWR VPWR _04565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15809_ net1587 _08354_ net1624 VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__o21ai_1
X_16789_ _04170_ _04492_ _04497_ _04180_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__o211a_1
X_09330_ _05642_ _05651_ _05681_ _05657_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__and4bb_1
X_18528_ net349 _02052_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09261_ CPU.aluIn1\[14\] _05543_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__nand2_1
X_15743__533 clknet_1_0__leaf__03652_ VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__inv_2
X_18459_ net280 _01987_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09192_ _05543_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__buf_2
XFILLER_0_16_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08506_ clknet_0__08506_ VGND VGND VPWR VPWR clknet_1_1__leaf__08506_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08437_ clknet_0__08437_ VGND VGND VPWR VPWR clknet_1_1__leaf__08437_
+ sky130_fd_sc_hd__clkbuf_16
X_14238__368 clknet_1_1__leaf__08508_ VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__inv_2
X_17720__51 clknet_1_0__leaf__05015_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__inv_2
XFILLER_0_30_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__08468_ _08468_ VGND VGND VPWR VPWR clknet_0__08468_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__08368_ clknet_0__08368_ VGND VGND VPWR VPWR clknet_1_1__leaf__08368_
+ sky130_fd_sc_hd__clkbuf_16
Xhold14 mapped_spi_ram.rcv_bitcount\[5\] VGND VGND VPWR VPWR net1311 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ _05326_ _05327_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__or2_2
Xhold25 _07828_ VGND VGND VPWR VPWR net1322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 _08242_ VGND VGND VPWR VPWR net1333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 _01730_ VGND VGND VPWR VPWR net1344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 mapped_spi_ram.cmd_addr\[4\] VGND VGND VPWR VPWR net1355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 mapped_spi_flash.rcv_data\[29\] VGND VGND VPWR VPWR net1366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09528_ _05872_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__clkbuf_4
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09459_ _05393_ _05522_ _05748_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12470_ net2097 _07314_ _07920_ VGND VGND VPWR VPWR _07922_ sky130_fd_sc_hd__mux2_1
X_13679__1054 clknet_1_0__leaf__08453_ VGND VGND VPWR VPWR net1110 sky130_fd_sc_hd__inv_2
XFILLER_0_152_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11421_ _07308_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11352_ net2355 _06555_ _07237_ VGND VGND VPWR VPWR _07272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15872__617 clknet_1_1__leaf__03682_ VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__inv_2
XFILLER_0_132_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10303_ net2077 _06555_ _06557_ VGND VGND VPWR VPWR _06592_ sky130_fd_sc_hd__mux2_1
X_11283_ _06661_ net2039 _07200_ VGND VGND VPWR VPWR _07235_ sky130_fd_sc_hd__mux2_1
X_13022_ net1866 _07376_ _08180_ VGND VGND VPWR VPWR _08215_ sky130_fd_sc_hd__mux2_1
X_10234_ _06554_ VGND VGND VPWR VPWR _06555_ sky130_fd_sc_hd__clkbuf_4
X_17830_ net910 _01392_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_10165_ CPU.PC\[1\] _05952_ VGND VGND VPWR VPWR _06488_ sky130_fd_sc_hd__nand2_1
X_13970__127 clknet_1_1__leaf__08481_ VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__inv_2
X_17761_ net841 _01323_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_10096_ _05883_ _06421_ VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__nor2_1
X_14973_ _02751_ _03035_ _03038_ _02759_ VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__a211o_1
X_16712_ _06149_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__clkbuf_4
X_17692_ CPU.mem_wdata\[0\] per_uart.d_in_uart\[0\] _05218_ VGND VGND VPWR VPWR _05219_
+ sky130_fd_sc_hd__mux2_1
X_16643_ CPU.registerFile\[28\]\[15\] CPU.registerFile\[29\]\[15\] _04122_ VGND VGND
+ VPWR VPWR _04355_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__08457_ clknet_0__08457_ VGND VGND VPWR VPWR clknet_1_0__leaf__08457_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12806_ _08099_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16574_ CPU.registerFile\[20\]\[13\] CPU.registerFile\[21\]\[13\] _04287_ VGND VGND
+ VPWR VPWR _04288_ sky130_fd_sc_hd__mux2_1
X_10998_ _07024_ _07026_ VGND VGND VPWR VPWR _07042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18313_ net134 _01841_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15525_ _03575_ _03576_ _03255_ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _06661_ net2621 _08028_ VGND VGND VPWR VPWR _08063_ sky130_fd_sc_hd__mux2_1
X_13881__1237 clknet_1_0__leaf__08472_ VGND VGND VPWR VPWR net1293 sky130_fd_sc_hd__inv_2
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ net1255 _01772_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15456_ _08580_ _03507_ _03509_ _03218_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__a211o_1
Xclkbuf_0__04982_ _04982_ VGND VGND VPWR VPWR clknet_0__04982_ sky130_fd_sc_hd__clkbuf_16
X_12668_ _08026_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__clkbuf_1
X_14407_ CPU.registerFile\[24\]\[2\] _08545_ _08650_ _08550_ VGND VGND VPWR VPWR _08651_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11619_ net2047 _07337_ _07427_ VGND VGND VPWR VPWR _07430_ sky130_fd_sc_hd__mux2_1
X_18175_ net1186 _01703_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[14\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_142_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15387_ CPU.registerFile\[15\]\[26\] CPU.registerFile\[14\]\[26\] _08560_ VGND VGND
+ VPWR VPWR _03443_ sky130_fd_sc_hd__mux2_1
X_12599_ net2405 _07374_ _07956_ VGND VGND VPWR VPWR _07990_ sky130_fd_sc_hd__mux2_1
X_17126_ CPU.registerFile\[24\]\[27\] _03724_ _04569_ _04825_ VGND VGND VPWR VPWR
+ _04826_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14338_ _08410_ VGND VGND VPWR VPWR _08584_ sky130_fd_sc_hd__clkbuf_8
Xhold506 CPU.registerFile\[9\]\[31\] VGND VGND VPWR VPWR net1803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold517 CPU.registerFile\[28\]\[15\] VGND VGND VPWR VPWR net1814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 CPU.registerFile\[13\]\[12\] VGND VGND VPWR VPWR net1825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 CPU.registerFile\[6\]\[1\] VGND VGND VPWR VPWR net1836 sky130_fd_sc_hd__dlygate4sd3_1
X_17057_ CPU.registerFile\[22\]\[25\] CPU.registerFile\[23\]\[25\] _03761_ VGND VGND
+ VPWR VPWR _04759_ sky130_fd_sc_hd__mux2_1
X_14269_ _05876_ VGND VGND VPWR VPWR _08515_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16008_ _03713_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 CPU.registerFile\[8\]\[4\] VGND VGND VPWR VPWR net2503 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1217 CPU.registerFile\[25\]\[4\] VGND VGND VPWR VPWR net2514 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ net970 _01487_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xhold1228 CPU.registerFile\[17\]\[11\] VGND VGND VPWR VPWR net2525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1239 CPU.registerFile\[25\]\[22\] VGND VGND VPWR VPWR net2536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17309__723 clknet_1_0__leaf__04981_ VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__inv_2
XFILLER_0_48_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15667__464 clknet_1_0__leaf__03645_ VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__inv_2
X_09313_ _05625_ _05617_ _05623_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__and3_1
XFILLER_0_158_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_721 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18591__48 VGND VGND VPWR VPWR _18591__48/HI net48 sky130_fd_sc_hd__conb_1
X_09244_ CPU.aluIn1\[11\] CPU.Bimm\[12\] VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__nor2_1
X_13235__757 clknet_1_0__leaf__08342_ VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__inv_2
XFILLER_0_91_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09175_ CPU.Jimm\[14\] CPU.Jimm\[13\] VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14171__308 clknet_1_1__leaf__08501_ VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__inv_2
XFILLER_0_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08959_ _05263_ _05265_ _05307_ _05308_ _05310_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__o311a_1
X_11970_ _07616_ VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__clkbuf_1
X_10921_ _06982_ VGND VGND VPWR VPWR _06983_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10852_ CPU.aluReg\[14\] _06928_ _06922_ VGND VGND VPWR VPWR _06929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10783_ _06875_ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__clkbuf_1
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15310_ CPU.registerFile\[24\]\[24\] _08582_ _03367_ _03175_ VGND VGND VPWR VPWR
+ _03368_ sky130_fd_sc_hd__o211a_1
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12522_ net2299 _07366_ _07942_ VGND VGND VPWR VPWR _07949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16290_ net2654 _03566_ _04010_ _03855_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_927 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15241_ CPU.registerFile\[15\]\[22\] CPU.registerFile\[14\]\[22\] _03013_ VGND VGND
+ VPWR VPWR _03301_ sky130_fd_sc_hd__mux2_1
X_12453_ _07912_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11404_ net1735 _06361_ _07296_ VGND VGND VPWR VPWR _07300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12384_ _06649_ net1888 _07870_ VGND VGND VPWR VPWR _07876_ sky130_fd_sc_hd__mux2_1
X_15172_ CPU.registerFile\[2\]\[20\] CPU.registerFile\[3\]\[20\] _02871_ VGND VGND
+ VPWR VPWR _03234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11335_ _07263_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18931_ net705 _02451_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_11266_ _07226_ VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__clkbuf_1
X_13005_ _08206_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__clkbuf_1
X_10217_ _05724_ _06534_ VGND VGND VPWR VPWR _06538_ sky130_fd_sc_hd__nor2_1
X_18862_ net636 _02382_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11197_ net1395 VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__inv_2
X_17813_ net893 _01375_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_10148_ net1438 _05859_ _05719_ per_uart.rx_data\[3\] _06471_ VGND VGND VPWR VPWR
+ _06472_ sky130_fd_sc_hd__a221o_1
X_18793_ net582 _02317_ VGND VGND VPWR VPWR CPU.aluReg\[23\] sky130_fd_sc_hd__dfxtp_1
X_17744_ net829 _01310_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_14956_ CPU.registerFile\[6\]\[15\] CPU.registerFile\[7\]\[15\] _02982_ VGND VGND
+ VPWR VPWR _03023_ sky130_fd_sc_hd__mux2_1
X_10079_ _05300_ _06373_ VGND VGND VPWR VPWR _06406_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17675_ _05180_ _05205_ _06855_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__and3b_1
Xclkbuf_1_0__f__08509_ clknet_0__08509_ VGND VGND VPWR VPWR clknet_1_0__leaf__08509_
+ sky130_fd_sc_hd__clkbuf_16
X_14887_ CPU.registerFile\[19\]\[14\] CPU.registerFile\[18\]\[14\] _02753_ VGND VGND
+ VPWR VPWR _02955_ sky130_fd_sc_hd__mux2_1
X_16626_ CPU.registerFile\[8\]\[15\] _04101_ _04102_ _04337_ VGND VGND VPWR VPWR _04338_
+ sky130_fd_sc_hd__o211a_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16557_ CPU.registerFile\[2\]\[13\] CPU.registerFile\[3\]\[13\] _04027_ VGND VGND
+ VPWR VPWR _04271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15508_ CPU.registerFile\[0\]\[29\] _08411_ _03560_ _06036_ VGND VGND VPWR VPWR _03561_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16488_ _04202_ _04203_ _03875_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18227_ net1238 _01755_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[28\] sky130_fd_sc_hd__dfxtp_1
X_15439_ _03485_ _03493_ _03241_ VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18158_ net1169 _01686_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_bitcount\[4\] sky130_fd_sc_hd__dfxtp_1
X_13527__918 clknet_1_0__leaf__08437_ VGND VGND VPWR VPWR net974 sky130_fd_sc_hd__inv_2
XFILLER_0_5_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold303 mapped_spi_flash.rcv_data\[14\] VGND VGND VPWR VPWR net1600 sky130_fd_sc_hd__clkdlybuf4s25_1
X_17109_ CPU.registerFile\[13\]\[27\] _03767_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__or2_1
Xhold314 mapped_spi_flash.rcv_data\[15\] VGND VGND VPWR VPWR net1611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold325 CPU.cycles\[7\] VGND VGND VPWR VPWR net1622 sky130_fd_sc_hd__dlygate4sd3_1
X_18089_ net1100 _01617_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold336 CPU.rs2\[13\] VGND VGND VPWR VPWR net1633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold347 CPU.rs2\[22\] VGND VGND VPWR VPWR net1644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 CPU.registerFile\[31\]\[1\] VGND VGND VPWR VPWR net1655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 CPU.rs2\[30\] VGND VGND VPWR VPWR net1666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09931_ CPU.PC\[12\] _05887_ VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03678_ clknet_0__03678_ VGND VGND VPWR VPWR clknet_1_1__leaf__03678_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _05911_ _06195_ _06196_ _06197_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__o22a_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1003 CPU.registerFile\[21\]\[13\] VGND VGND VPWR VPWR net2300 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13678__1053 clknet_1_0__leaf__08453_ VGND VGND VPWR VPWR net1109 sky130_fd_sc_hd__inv_2
Xhold1014 CPU.registerFile\[22\]\[27\] VGND VGND VPWR VPWR net2311 sky130_fd_sc_hd__dlygate4sd3_1
X_09793_ _05425_ _06130_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1025 CPU.registerFile\[16\]\[4\] VGND VGND VPWR VPWR net2322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 CPU.registerFile\[16\]\[10\] VGND VGND VPWR VPWR net2333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 CPU.registerFile\[28\]\[0\] VGND VGND VPWR VPWR net2344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 CPU.registerFile\[2\]\[0\] VGND VGND VPWR VPWR net2355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1069 CPU.registerFile\[3\]\[11\] VGND VGND VPWR VPWR net2366 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09227_ CPU.aluIn1\[1\] _05578_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_118_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09158_ _05410_ _05408_ _05506_ _05509_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09089_ _05435_ _05439_ _05440_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11120_ net1438 _07133_ _07140_ _07138_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__o211a_1
Xhold870 CPU.registerFile\[26\]\[16\] VGND VGND VPWR VPWR net2167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 CPU.registerFile\[16\]\[29\] VGND VGND VPWR VPWR net2178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 CPU.registerFile\[21\]\[1\] VGND VGND VPWR VPWR net2189 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ net1505 _07054_ _07088_ _07069_ VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__o211a_1
X_13759__1127 clknet_1_0__leaf__08460_ VGND VGND VPWR VPWR net1183 sky130_fd_sc_hd__inv_2
X_10002_ mapped_spi_ram.rcv_data\[17\] _05685_ VGND VGND VPWR VPWR _06332_ sky130_fd_sc_hd__and2_1
X_13880__1236 clknet_1_0__leaf__08472_ VGND VGND VPWR VPWR net1292 sky130_fd_sc_hd__inv_2
X_14810_ CPU.registerFile\[17\]\[12\] _08795_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__or2_1
X_15790_ _03660_ _03662_ _08347_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__or3b_1
X_14741_ CPU.registerFile\[24\]\[10\] _08686_ _02812_ _02771_ VGND VGND VPWR VPWR
+ _02813_ sky130_fd_sc_hd__o211a_1
X_11953_ _07607_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17460_ _05016_ CPU.PC\[7\] _05043_ _05044_ _07002_ VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__o221a_1
X_10904_ CPU.aluIn1\[1\] _06967_ _06880_ VGND VGND VPWR VPWR _06968_ sky130_fd_sc_hd__mux2_1
X_14672_ _05876_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11884_ _06613_ net2351 _07562_ VGND VGND VPWR VPWR _07571_ sky130_fd_sc_hd__mux2_1
X_16411_ _04075_ _04124_ _04128_ _04042_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__o211a_1
X_10835_ net2662 _06915_ _06889_ VGND VGND VPWR VPWR _06916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_16
X_19130_ clknet_leaf_10_clk _02650_ VGND VGND VPWR VPWR CPU.PC\[12\] sky130_fd_sc_hd__dfxtp_2
X_16342_ CPU.registerFile\[13\]\[8\] _03976_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__or2_1
X_13554_ clknet_1_1__leaf__08440_ VGND VGND VPWR VPWR _08441_ sky130_fd_sc_hd__buf_1
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10766_ CPU.aluShamt\[4\] _06859_ VGND VGND VPWR VPWR _06860_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12505_ net2399 _07349_ _07931_ VGND VGND VPWR VPWR _07940_ sky130_fd_sc_hd__mux2_1
X_19061_ net803 _02581_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16273_ _03992_ _03993_ _03875_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__mux2_1
X_10697_ net2438 _05825_ _06816_ VGND VGND VPWR VPWR _06821_ sky130_fd_sc_hd__mux2_1
X_18012_ net1023 _01540_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15224_ CPU.registerFile\[17\]\[22\] _03036_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12436_ _07903_ VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15155_ CPU.registerFile\[24\]\[20\] _02928_ _03216_ _03175_ VGND VGND VPWR VPWR
+ _03217_ sky130_fd_sc_hd__o211a_1
X_12367_ _06632_ net2045 _07859_ VGND VGND VPWR VPWR _07867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11318_ _07254_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__clkbuf_1
X_15086_ _03027_ _03147_ _03149_ _03111_ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__a211o_1
X_12298_ net1469 _07812_ _07824_ _07822_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__o211a_1
X_18914_ net688 _02434_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_11249_ _07217_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13264__783 clknet_1_1__leaf__08345_ VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__inv_2
X_18845_ clknet_leaf_7_clk _02369_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_15850__597 clknet_1_1__leaf__03680_ VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__inv_2
X_18776_ net565 _02300_ VGND VGND VPWR VPWR CPU.aluReg\[6\] sky130_fd_sc_hd__dfxtp_1
X_15988_ _03703_ _03706_ _03711_ _03714_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17727_ net812 _01293_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_14939_ _06418_ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17658_ net1453 _05189_ _05193_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16609_ _04037_ _04318_ _04321_ _04208_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__a211o_1
XFILLER_0_147_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17589_ per_uart.uart0.tx_bitcount\[0\] _05116_ _05120_ _05148_ _06854_ VGND VGND
+ VPWR VPWR _05149_ sky130_fd_sc_hd__o311a_1
XFILLER_0_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09012_ CPU.aluIn1\[20\] _05362_ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15779__565 clknet_1_1__leaf__03656_ VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__inv_2
XFILLER_0_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold100 _08240_ VGND VGND VPWR VPWR net1397 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold111 mapped_spi_ram.cmd_addr\[20\] VGND VGND VPWR VPWR net1408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 mapped_spi_flash.rcv_data\[10\] VGND VGND VPWR VPWR net1419 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold133 _01716_ VGND VGND VPWR VPWR net1430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 CPU.aluReg\[26\] VGND VGND VPWR VPWR net1441 sky130_fd_sc_hd__dlygate4sd3_1
X_13308__809 clknet_1_1__leaf__08362_ VGND VGND VPWR VPWR net865 sky130_fd_sc_hd__inv_2
Xhold155 _02673_ VGND VGND VPWR VPWR net1452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 per_uart.uart0.txd_reg\[1\] VGND VGND VPWR VPWR net1463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 per_uart.uart0.txd_reg\[3\] VGND VGND VPWR VPWR net1474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 mapped_spi_ram.cmd_addr\[17\] VGND VGND VPWR VPWR net1485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold199 mapped_spi_ram.rcv_data\[14\] VGND VGND VPWR VPWR net1496 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ mapped_spi_ram.rcv_data\[20\] _05761_ _05762_ mapped_spi_flash.rcv_data\[20\]
+ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09845_ _06180_ _05455_ _05319_ VGND VGND VPWR VPWR _06181_ sky130_fd_sc_hd__o21ai_2
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ _05424_ _06112_ _06114_ _05516_ VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__o211a_1
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_917 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10620_ net2521 _05767_ _06777_ VGND VGND VPWR VPWR _06779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10551_ _06741_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13270_ per_uart.uart0.enable16_counter\[6\] _08350_ VGND VGND VPWR VPWR _08351_
+ sky130_fd_sc_hd__or2_1
X_10482_ _06704_ VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__clkbuf_1
X_12221_ _07778_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__clkbuf_1
X_12152_ _07715_ _07729_ VGND VGND VPWR VPWR _07730_ sky130_fd_sc_hd__or2_1
X_13924__85 clknet_1_0__leaf__08477_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__inv_2
X_11103_ mapped_spi_flash.rcv_bitcount\[3\] _07126_ VGND VGND VPWR VPWR _07127_ sky130_fd_sc_hd__or2_1
X_16960_ CPU.registerFile\[10\]\[23\] CPU.registerFile\[11\]\[23\] _04335_ VGND VGND
+ VPWR VPWR _04664_ sky130_fd_sc_hd__mux2_1
X_12083_ _07670_ _07680_ _07674_ _07677_ CPU.mem_wbusy VGND VGND VPWR VPWR _07681_
+ sky130_fd_sc_hd__a32o_1
X_11034_ mapped_spi_flash.cmd_addr\[8\] _07073_ _07039_ VGND VGND VPWR VPWR _07074_
+ sky130_fd_sc_hd__mux2_1
X_15911_ clknet_1_1__leaf__03686_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__buf_1
X_16891_ CPU.registerFile\[5\]\[21\] CPU.registerFile\[4\]\[21\] _04428_ VGND VGND
+ VPWR VPWR _04597_ sky130_fd_sc_hd__mux2_1
X_18630_ clknet_leaf_24_clk _02154_ VGND VGND VPWR VPWR CPU.mem_wdata\[2\] sky130_fd_sc_hd__dfxtp_4
X_18561_ net382 _02085_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_12985_ net1907 _07339_ _08192_ VGND VGND VPWR VPWR _08196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17512_ _05069_ net2605 _05086_ _05087_ _05053_ VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__o221a_1
X_14724_ net2051 _08514_ _02796_ _08751_ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__o211a_1
X_18492_ net313 _02016_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_11936_ _06593_ net2312 _07598_ VGND VGND VPWR VPWR _07599_ sky130_fd_sc_hd__mux2_1
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17443_ _08311_ _06453_ _08331_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__or3_1
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14655_ CPU.registerFile\[15\]\[8\] CPU.registerFile\[14\]\[8\] _08771_ VGND VGND
+ VPWR VPWR _02729_ sky130_fd_sc_hd__mux2_1
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _07561_ VGND VGND VPWR VPWR _07562_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10818_ _06902_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__clkbuf_1
X_17374_ _04996_ _05001_ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__and2_1
X_14586_ CPU.registerFile\[2\]\[6\] CPU.registerFile\[3\]\[6\] _08629_ VGND VGND VPWR
+ VPWR _08826_ sky130_fd_sc_hd__mux2_1
X_11798_ _06774_ _07451_ VGND VGND VPWR VPWR _07525_ sky130_fd_sc_hd__nor2_4
XFILLER_0_28_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19113_ net96 _02633_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_16325_ CPU.registerFile\[20\]\[7\] CPU.registerFile\[21\]\[7\] _03883_ VGND VGND
+ VPWR VPWR _04045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10749_ net2567 _06508_ _06838_ VGND VGND VPWR VPWR _06848_ sky130_fd_sc_hd__mux2_1
X_13677__1052 clknet_1_0__leaf__08453_ VGND VGND VPWR VPWR net1108 sky130_fd_sc_hd__inv_2
XFILLER_0_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19044_ net786 _02564_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16256_ CPU.registerFile\[13\]\[6\] _03976_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_1__f__08470_ clknet_0__08470_ VGND VGND VPWR VPWR clknet_1_1__leaf__08470_
+ sky130_fd_sc_hd__clkbuf_16
X_13468_ _06339_ VGND VGND VPWR VPWR _08425_ sky130_fd_sc_hd__buf_2
XFILLER_0_113_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15207_ _08549_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__clkbuf_4
X_12419_ _07894_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16187_ _08404_ _03896_ _03900_ _03909_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__a31o_2
XFILLER_0_112_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13399_ CPU.instr\[2\] _06493_ _00000_ VGND VGND VPWR VPWR _08378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15138_ net1627 _02797_ _03200_ _02993_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15069_ _08532_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_4_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_16
X_09630_ CPU.PC\[10\] CPU.Bimm\[10\] _05914_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__and3_1
X_18828_ net617 _02352_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_09561_ _05424_ _05904_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__nand2_1
X_17424__45 clknet_1_1__leaf__05015_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__inv_2
X_18759_ net548 _02283_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[21\] sky130_fd_sc_hd__dfxtp_1
X_09492_ _05838_ VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13758__1126 clknet_1_0__leaf__08460_ VGND VGND VPWR VPWR net1182 sky130_fd_sc_hd__inv_2
XFILLER_0_129_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13505__898 clknet_1_1__leaf__08435_ VGND VGND VPWR VPWR net954 sky130_fd_sc_hd__inv_2
X_13360__855 clknet_1_0__leaf__08368_ VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__inv_2
X_09828_ _06161_ _06163_ _06164_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__or3_1
Xclkbuf_1_0__f__08490_ clknet_0__08490_ VGND VGND VPWR VPWR clknet_1_0__leaf__08490_
+ sky130_fd_sc_hd__clkbuf_16
X_09759_ _05350_ _06089_ _06098_ VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__o21ai_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _06626_ net2252 _08076_ VGND VGND VPWR VPWR _08081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ net2482 _07370_ _07475_ VGND VGND VPWR VPWR _07484_ sky130_fd_sc_hd__mux2_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_920 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ CPU.registerFile\[28\]\[3\] CPU.registerFile\[29\]\[3\] _08538_ VGND VGND
+ VPWR VPWR _08683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11652_ net2395 _07370_ _07438_ VGND VGND VPWR VPWR _07447_ sky130_fd_sc_hd__mux2_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10603_ _06768_ VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14371_ _08515_ _08602_ _08606_ _08615_ VGND VGND VPWR VPWR _08616_ sky130_fd_sc_hd__a31o_1
XFILLER_0_153_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11583_ net1693 _07370_ _07401_ VGND VGND VPWR VPWR _07410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16110_ CPU.registerFile\[28\]\[2\] CPU.registerFile\[29\]\[2\] _03739_ VGND VGND
+ VPWR VPWR _03835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13322_ clknet_1_1__leaf__08341_ VGND VGND VPWR VPWR _08364_ sky130_fd_sc_hd__buf_1
X_17090_ CPU.registerFile\[24\]\[26\] _03724_ _04569_ _04790_ VGND VGND VPWR VPWR
+ _04791_ sky130_fd_sc_hd__o211a_1
X_10534_ _06731_ VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16041_ CPU.registerFile\[19\]\[0\] CPU.registerFile\[18\]\[0\] _03767_ VGND VGND
+ VPWR VPWR _03768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10465_ _06694_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12204_ net1308 _07764_ mapped_spi_ram.snd_bitcount\[5\] _07765_ VGND VGND VPWR VPWR
+ _01726_ sky130_fd_sc_hd__a2bb2o_1
X_10396_ _06655_ net1861 _06639_ VGND VGND VPWR VPWR _06656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13184_ CPU.cycles\[27\] _08301_ VGND VGND VPWR VPWR _08303_ sky130_fd_sc_hd__and2_1
X_15916__656 clknet_1_1__leaf__03687_ VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__inv_2
X_12135_ mapped_spi_ram.cmd_addr\[19\] _07038_ _07704_ VGND VGND VPWR VPWR _07718_
+ sky130_fd_sc_hd__mux2_1
X_17992_ net1003 _01520_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16943_ _04484_ _04485_ CPU.registerFile\[25\]\[22\] VGND VGND VPWR VPWR _04648_
+ sky130_fd_sc_hd__a21o_1
X_12066_ _07667_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__clkbuf_1
X_11017_ _05595_ _05596_ _05597_ _07057_ VGND VGND VPWR VPWR _07059_ sky130_fd_sc_hd__or4_1
X_16874_ _04579_ _04580_ CPU.registerFile\[17\]\[20\] VGND VGND VPWR VPWR _04581_
+ sky130_fd_sc_hd__a21o_1
X_18613_ net434 _02137_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18544_ net365 _02068_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_12968_ net2113 _07322_ _08181_ VGND VGND VPWR VPWR _08187_ sky130_fd_sc_hd__mux2_1
X_13337__835 clknet_1_0__leaf__08365_ VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__inv_2
X_14707_ CPU.registerFile\[10\]\[9\] CPU.registerFile\[11\]\[9\] _02779_ VGND VGND
+ VPWR VPWR _02780_ sky130_fd_sc_hd__mux2_1
X_18475_ net296 _01999_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11919_ _07589_ VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__clkbuf_1
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15962__698 clknet_1_0__leaf__03691_ VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__inv_2
X_12899_ _08150_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ _08255_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_942 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14638_ CPU.registerFile\[17\]\[8\] _08795_ VGND VGND VPWR VPWR _08876_ sky130_fd_sc_hd__or2_1
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17357_ per_uart.uart0.rx_count16\[3\] per_uart.uart0.rx_count16\[2\] _04987_ VGND
+ VGND VPWR VPWR _04988_ sky130_fd_sc_hd__or3_1
X_17303__718 clknet_1_1__leaf__04980_ VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__inv_2
X_14569_ _06059_ VGND VGND VPWR VPWR _08809_ sky130_fd_sc_hd__clkbuf_4
X_15661__459 clknet_1_0__leaf__03644_ VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__inv_2
XFILLER_0_43_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16308_ CPU.registerFile\[2\]\[7\] CPU.registerFile\[3\]\[7\] _04027_ VGND VGND VPWR
+ VPWR _04028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19027_ net769 _02547_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_16239_ _03741_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__buf_4
XFILLER_0_113_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__08453_ clknet_0__08453_ VGND VGND VPWR VPWR clknet_1_1__leaf__08453_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08484_ _08484_ VGND VGND VPWR VPWR clknet_0__08484_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08992_ _05336_ _05338_ _05343_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__a21oi_4
X_13903__66 clknet_1_1__leaf__08475_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__inv_2
X_14132__272 clknet_1_0__leaf__08498_ VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__inv_2
X_09613_ CPU.PC\[1\] _05952_ _05955_ _05956_ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__a31o_1
X_09544_ CPU.PC\[13\] CPU.PC\[12\] _05887_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09475_ _05556_ _05822_ _05731_ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_690 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15720__512 clknet_1_0__leaf__03650_ VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__inv_2
XFILLER_0_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13585__970 clknet_1_1__leaf__08443_ VGND VGND VPWR VPWR net1026 sky130_fd_sc_hd__inv_2
XFILLER_0_21_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10250_ _06564_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__clkbuf_1
X_15638__439 clknet_1_1__leaf__03641_ VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__inv_2
X_10181_ _05517_ _06499_ _06502_ _06503_ _05271_ VGND VGND VPWR VPWR _06504_ sky130_fd_sc_hd__a32o_1
XFILLER_0_30_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__08473_ clknet_0__08473_ VGND VGND VPWR VPWR clknet_1_0__leaf__08473_
+ sky130_fd_sc_hd__clkbuf_16
X_12822_ _05734_ net2426 _08109_ VGND VGND VPWR VPWR _08110_ sky130_fd_sc_hd__mux2_1
X_16590_ CPU.registerFile\[12\]\[14\] _04017_ _04018_ _04302_ VGND VGND VPWR VPWR
+ _04303_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17403__26 clknet_1_0__leaf__05013_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__inv_2
X_15541_ CPU.registerFile\[5\]\[30\] CPU.registerFile\[4\]\[30\] _08558_ VGND VGND
+ VPWR VPWR _03593_ sky130_fd_sc_hd__mux2_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12753_ _06609_ net2196 _08065_ VGND VGND VPWR VPWR _08072_ sky130_fd_sc_hd__mux2_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _07452_ VGND VGND VPWR VPWR _07475_ sky130_fd_sc_hd__clkbuf_4
X_18260_ net1271 _01788_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15472_ CPU.registerFile\[0\]\[28\] _08411_ _03525_ _03195_ VGND VGND VPWR VPWR _03526_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12684_ _08035_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14261__389 clknet_1_0__leaf__08510_ VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__inv_2
XFILLER_0_126_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17211_ net2540 _08513_ _04908_ _04663_ VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14423_ CPU.registerFile\[2\]\[2\] CPU.registerFile\[3\]\[2\] _08629_ VGND VGND VPWR
+ VPWR _08667_ sky130_fd_sc_hd__mux2_1
X_11635_ _07415_ VGND VGND VPWR VPWR _07438_ sky130_fd_sc_hd__clkbuf_4
X_18191_ net1202 _01719_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17142_ CPU.registerFile\[8\]\[28\] _04505_ _04506_ _04840_ VGND VGND VPWR VPWR _04841_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14354_ CPU.registerFile\[19\]\[1\] CPU.registerFile\[18\]\[1\] _06064_ VGND VGND
+ VPWR VPWR _08599_ sky130_fd_sc_hd__mux2_1
X_11566_ _07378_ VGND VGND VPWR VPWR _07401_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17073_ CPU.registerFile\[13\]\[26\] _03767_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10517_ _06722_ VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__clkbuf_1
X_14285_ CPU.registerFile\[20\]\[0\] _08527_ _08529_ _08530_ VGND VGND VPWR VPWR _08531_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11497_ net2380 _07360_ _07354_ VGND VGND VPWR VPWR _07361_ sky130_fd_sc_hd__mux2_1
X_16024_ _03750_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__clkbuf_4
X_10448_ _06685_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13167_ CPU.cycles\[19\] CPU.cycles\[20\] _08291_ VGND VGND VPWR VPWR _08293_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10379_ _06644_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12118_ net1316 _07693_ _07705_ _07175_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__o211a_1
X_17975_ net986 _01503_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_13098_ net1652 _06975_ _06856_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__o21a_1
X_13757__1125 clknet_1_0__leaf__08460_ VGND VGND VPWR VPWR net1181 sky130_fd_sc_hd__inv_2
X_16926_ CPU.registerFile\[12\]\[22\] _04421_ _04422_ _04630_ VGND VGND VPWR VPWR
+ _04631_ sky130_fd_sc_hd__o211a_1
X_12049_ CPU.registerFile\[24\]\[10\] _07356_ _07657_ VGND VGND VPWR VPWR _07659_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16857_ _04502_ _04549_ _04554_ _04563_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__a31o_2
X_15808_ _08355_ _03672_ _03661_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__a21oi_1
X_16788_ _04367_ _04493_ _04496_ _04410_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__a211o_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18527_ net348 _02051_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09260_ _05611_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__inv_2
X_18458_ net279 _01986_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09191_ CPU.Bimm\[12\] VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__buf_2
X_17409_ clknet_1_1__leaf__08340_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__buf_1
XFILLER_0_145_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18389_ net210 _01917_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__08505_ clknet_0__08505_ VGND VGND VPWR VPWR clknet_1_1__leaf__08505_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__08436_ clknet_0__08436_ VGND VGND VPWR VPWR clknet_1_1__leaf__08436_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08467_ _08467_ VGND VGND VPWR VPWR clknet_0__08467_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08367_ clknet_0__08367_ VGND VGND VPWR VPWR clknet_1_1__leaf__08367_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08975_ CPU.aluIn1\[15\] _05325_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__nor2_1
Xhold15 net2674 VGND VGND VPWR VPWR net1312 sky130_fd_sc_hd__buf_4
Xhold26 _07830_ VGND VGND VPWR VPWR net1323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 mapped_spi_ram.cmd_addr\[24\] VGND VGND VPWR VPWR net1334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 mapped_spi_ram.cmd_addr\[2\] VGND VGND VPWR VPWR net1345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 mapped_spi_flash.rcv_data\[24\] VGND VGND VPWR VPWR net1356 sky130_fd_sc_hd__dlygate4sd3_1
X_09527_ _05764_ _05862_ _05871_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__a21o_4
X_15945__682 clknet_1_0__leaf__03690_ VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__inv_2
X_13617__999 clknet_1_1__leaf__08446_ VGND VGND VPWR VPWR net1055 sky130_fd_sc_hd__inv_2
XFILLER_0_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09458_ _05806_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09389_ _05735_ _05736_ _05740_ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_47_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17343__4 clknet_1_1__leaf__04984_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__inv_2
XFILLER_0_152_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11420_ net2344 _06555_ _07273_ VGND VGND VPWR VPWR _07308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11351_ _07271_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10302_ _06591_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__clkbuf_1
X_13817__1179 clknet_1_0__leaf__08466_ VGND VGND VPWR VPWR net1235 sky130_fd_sc_hd__inv_2
XFILLER_0_21_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11282_ _07234_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13366__861 clknet_1_1__leaf__08368_ VGND VGND VPWR VPWR net917 sky130_fd_sc_hd__inv_2
X_13021_ _08214_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__clkbuf_1
X_10233_ CPU.cycles\[0\] _05759_ _06176_ net1357 _06553_ VGND VGND VPWR VPWR _06554_
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_30_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10164_ _06487_ VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__clkbuf_1
X_17332__744 clknet_1_0__leaf__04983_ VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__inv_2
X_15690__485 clknet_1_0__leaf__03647_ VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__inv_2
X_17760_ net840 _01322_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_10095_ CPU.PC\[5\] _05882_ VGND VGND VPWR VPWR _06421_ sky130_fd_sc_hd__nor2_1
X_14972_ CPU.registerFile\[16\]\[16\] _02755_ _03037_ _02757_ VGND VGND VPWR VPWR
+ _03038_ sky130_fd_sc_hd__o211a_1
X_16711_ _08393_ VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__clkbuf_4
X_17691_ _05719_ _07673_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__nand2_4
XFILLER_0_159_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16642_ CPU.registerFile\[30\]\[15\] CPU.registerFile\[31\]\[15\] _04201_ VGND VGND
+ VPWR VPWR _04354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__08456_ clknet_0__08456_ VGND VGND VPWR VPWR clknet_1_0__leaf__08456_
+ sky130_fd_sc_hd__clkbuf_16
X_12805_ _06661_ net2483 _08064_ VGND VGND VPWR VPWR _08099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16573_ _03736_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__buf_4
X_10997_ net1504 _07007_ _07041_ _07014_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15524_ CPU.registerFile\[28\]\[30\] CPU.registerFile\[29\]\[30\] _08410_ VGND VGND
+ VPWR VPWR _03576_ sky130_fd_sc_hd__mux2_1
X_18312_ net133 _01840_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _08062_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ net1254 _01771_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__04981_ _04981_ VGND VGND VPWR VPWR clknet_0__04981_ sky130_fd_sc_hd__clkbuf_16
X_15455_ CPU.registerFile\[24\]\[28\] _08582_ _03508_ _03175_ VGND VGND VPWR VPWR
+ _03509_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12667_ _06659_ net2234 _07992_ VGND VGND VPWR VPWR _08026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14406_ _08546_ _08547_ CPU.registerFile\[25\]\[2\] VGND VGND VPWR VPWR _08650_ sky130_fd_sc_hd__a21o_1
X_11618_ _07429_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__clkbuf_1
X_18174_ net1185 net1483 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[13\] sky130_fd_sc_hd__dfxtp_1
X_15386_ _03202_ _03429_ _03433_ _03441_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__a31o_1
XFILLER_0_108_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12598_ _07989_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17125_ _04484_ _04485_ CPU.registerFile\[25\]\[27\] VGND VGND VPWR VPWR _04825_
+ sky130_fd_sc_hd__a21o_1
X_14337_ CPU.registerFile\[2\]\[0\] CPU.registerFile\[3\]\[0\] _08582_ VGND VGND VPWR
+ VPWR _08583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11549_ _07392_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold507 CPU.registerFile\[13\]\[9\] VGND VGND VPWR VPWR net1804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 CPU.registerFile\[6\]\[26\] VGND VGND VPWR VPWR net1815 sky130_fd_sc_hd__dlygate4sd3_1
X_17056_ _04479_ _04753_ _04757_ _04446_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__o211a_1
Xhold529 CPU.registerFile\[28\]\[21\] VGND VGND VPWR VPWR net1826 sky130_fd_sc_hd__dlygate4sd3_1
X_14268_ _08513_ VGND VGND VPWR VPWR _08514_ sky130_fd_sc_hd__buf_2
X_16007_ _08404_ _03701_ _03715_ _03733_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__a31o_1
XFILLER_0_150_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13219_ _05241_ _08310_ CPU.instr\[2\] VGND VGND VPWR VPWR _08333_ sky130_fd_sc_hd__or3b_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1207 CPU.registerFile\[26\]\[5\] VGND VGND VPWR VPWR net2504 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ net969 _01486_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[28\] sky130_fd_sc_hd__dfxtp_1
Xhold1218 CPU.registerFile\[26\]\[4\] VGND VGND VPWR VPWR net2515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1229 CPU.registerFile\[8\]\[20\] VGND VGND VPWR VPWR net2526 sky130_fd_sc_hd__dlygate4sd3_1
X_16909_ CPU.registerFile\[22\]\[21\] CPU.registerFile\[23\]\[21\] _04362_ VGND VGND
+ VPWR VPWR _04615_ sky130_fd_sc_hd__mux2_1
X_17889_ _00012_ _00014_ VGND VGND VPWR VPWR CPU.mem_rstrb sky130_fd_sc_hd__dlxtn_1
XFILLER_0_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09312_ _05617_ _05623_ _05625_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14244__373 clknet_1_0__leaf__08509_ VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__inv_2
XFILLER_0_146_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09243_ CPU.aluIn1\[11\] CPU.Bimm\[12\] VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09174_ CPU.Jimm\[12\] VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__buf_4
XFILLER_0_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08958_ _05261_ _05309_ VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__nor2_2
X_08889_ CPU.instr\[4\] CPU.instr\[6\] CPU.instr\[5\] VGND VGND VPWR VPWR _05241_
+ sky130_fd_sc_hd__nand3b_4
X_10920_ mapped_spi_flash.state\[2\] mapped_spi_flash.state\[1\] _06981_ VGND VGND
+ VPWR VPWR _06982_ sky130_fd_sc_hd__o21ai_1
X_18567__24 VGND VGND VPWR VPWR _18567__24/HI net24 sky130_fd_sc_hd__conb_1
X_10851_ CPU.aluIn1\[14\] _06927_ _06914_ VGND VGND VPWR VPWR _06928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13550__939 clknet_1_1__leaf__08439_ VGND VGND VPWR VPWR net995 sky130_fd_sc_hd__inv_2
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10782_ net2643 _06874_ _06869_ VGND VGND VPWR VPWR _06875_ sky130_fd_sc_hd__mux2_1
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12521_ _07948_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15240_ _03202_ _03286_ _03290_ _03299_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__a31o_1
XFILLER_0_136_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12452_ net1910 _07364_ _07906_ VGND VGND VPWR VPWR _07912_ sky130_fd_sc_hd__mux2_1
X_13756__1124 clknet_1_0__leaf__08460_ VGND VGND VPWR VPWR net1180 sky130_fd_sc_hd__inv_2
XFILLER_0_125_939 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11403_ _07299_ VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15171_ _03231_ _03232_ _03025_ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__mux2_1
X_12383_ _07875_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11334_ net2618 _06337_ _07260_ VGND VGND VPWR VPWR _07263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14053_ clknet_1_0__leaf__08484_ VGND VGND VPWR VPWR _08490_ sky130_fd_sc_hd__buf_1
X_18930_ net704 _02450_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_11265_ _06643_ net2033 _07223_ VGND VGND VPWR VPWR _07226_ sky130_fd_sc_hd__mux2_1
X_13004_ net1734 _07358_ _08203_ VGND VGND VPWR VPWR _08206_ sky130_fd_sc_hd__mux2_1
X_10216_ _06339_ _06341_ _06203_ VGND VGND VPWR VPWR _06537_ sky130_fd_sc_hd__mux2_1
X_18861_ net635 _02381_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_11196_ _07129_ net1394 _05703_ VGND VGND VPWR VPWR _07187_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17812_ net892 _01374_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_10147_ mapped_spi_ram.rcv_data\[27\] _05761_ VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18792_ net581 _02316_ VGND VGND VPWR VPWR CPU.aluReg\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17743_ net828 _01309_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_14955_ _02728_ _03016_ _03021_ _02784_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__o211a_1
X_10078_ _05447_ _06404_ VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__and2_1
Xclkbuf_1_0__f__08508_ clknet_0__08508_ VGND VGND VPWR VPWR clknet_1_0__leaf__08508_
+ sky130_fd_sc_hd__clkbuf_16
X_17674_ _05179_ per_uart.rx_error _05168_ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__a21o_1
X_14886_ net1633 _02797_ _02954_ _08751_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16625_ CPU.registerFile\[9\]\[15\] _04056_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_0__f__08439_ clknet_0__08439_ VGND VGND VPWR VPWR clknet_1_0__leaf__08439_
+ sky130_fd_sc_hd__clkbuf_16
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16556_ _04268_ _04269_ _04153_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15507_ _03235_ _03236_ CPU.registerFile\[1\]\[29\] VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__a21o_1
X_12719_ _06643_ net2568 _08051_ VGND VGND VPWR VPWR _08054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16487_ CPU.registerFile\[28\]\[11\] CPU.registerFile\[29\]\[11\] _04122_ VGND VGND
+ VPWR VPWR _04203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18226_ net1237 _01754_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[27\] sky130_fd_sc_hd__dfxtp_1
X_15438_ _03230_ _03488_ _03492_ _03151_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18157_ net1168 _01685_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_bitcount\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15369_ net1594 _03201_ _03425_ _03390_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17108_ CPU.registerFile\[15\]\[27\] CPU.registerFile\[14\]\[27\] _04550_ VGND VGND
+ VPWR VPWR _04808_ sky130_fd_sc_hd__mux2_1
Xhold304 _08227_ VGND VGND VPWR VPWR net1601 sky130_fd_sc_hd__dlygate4sd3_1
X_18088_ net1099 _01616_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[30\] sky130_fd_sc_hd__dfxtp_1
Xhold315 CPU.registerFile\[31\]\[9\] VGND VGND VPWR VPWR net1612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 CPU.state\[3\] VGND VGND VPWR VPWR net1623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 CPU.aluShamt\[0\] VGND VGND VPWR VPWR net1634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 CPU.cycles\[25\] VGND VGND VPWR VPWR net1645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17039_ _04419_ _04738_ _04740_ _04383_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__a211o_1
X_09930_ _05977_ _06262_ VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__xor2_1
XFILLER_0_110_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold359 CPU.rs2\[17\] VGND VGND VPWR VPWR net1656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ _05881_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__buf_2
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _05477_ _06093_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__xor2_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1004 CPU.registerFile\[16\]\[3\] VGND VGND VPWR VPWR net2301 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1015 CPU.registerFile\[23\]\[31\] VGND VGND VPWR VPWR net2312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1026 CPU.registerFile\[3\]\[22\] VGND VGND VPWR VPWR net2323 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1037 CPU.registerFile\[31\]\[4\] VGND VGND VPWR VPWR net2334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 CPU.registerFile\[7\]\[2\] VGND VGND VPWR VPWR net2345 sky130_fd_sc_hd__dlygate4sd3_1
X_13241__762 clknet_1_0__leaf__08343_ VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__inv_2
Xhold1059 CPU.registerFile\[16\]\[18\] VGND VGND VPWR VPWR net2356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13816__1178 clknet_1_0__leaf__08466_ VGND VGND VPWR VPWR net1234 sky130_fd_sc_hd__inv_2
XFILLER_0_9_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09226_ CPU.Iimm\[1\] CPU.Bimm\[1\] CPU.instr\[5\] VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__mux2_4
XFILLER_0_119_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09157_ _05408_ _05507_ _05508_ VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09088_ CPU.aluIn1\[2\] _05270_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__xor2_2
XFILLER_0_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold860 CPU.registerFile\[19\]\[22\] VGND VGND VPWR VPWR net2157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 CPU.registerFile\[13\]\[23\] VGND VGND VPWR VPWR net2168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold882 CPU.registerFile\[4\]\[23\] VGND VGND VPWR VPWR net2179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 CPU.registerFile\[3\]\[14\] VGND VGND VPWR VPWR net2190 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ _07048_ _07087_ VGND VGND VPWR VPWR _07088_ sky130_fd_sc_hd__or2_1
X_10001_ _05912_ _06328_ _06330_ VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14740_ _08808_ _08809_ CPU.registerFile\[25\]\[10\] VGND VGND VPWR VPWR _02812_
+ sky130_fd_sc_hd__a21o_1
X_11952_ _06613_ net2551 _07598_ VGND VGND VPWR VPWR _07607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10903_ CPU.aluReg\[2\] CPU.aluReg\[0\] _06939_ VGND VGND VPWR VPWR _06967_ sky130_fd_sc_hd__mux2_1
X_14671_ _08785_ _02742_ _02744_ _08870_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11883_ _07570_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__clkbuf_1
X_16410_ _04037_ _04125_ _04127_ _03803_ VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10834_ CPU.aluIn1\[18\] _06913_ _06914_ VGND VGND VPWR VPWR _06915_ sky130_fd_sc_hd__mux2_1
X_17390_ _05012_ VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16341_ CPU.registerFile\[15\]\[8\] CPU.registerFile\[14\]\[8\] _03705_ VGND VGND
+ VPWR VPWR _04060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13553_ clknet_1_0__leaf__08340_ VGND VGND VPWR VPWR _08440_ sky130_fd_sc_hd__buf_1
XFILLER_0_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10765_ CPU.aluShamt\[3\] CPU.aluShamt\[2\] CPU.aluShamt\[1\] CPU.aluShamt\[0\] VGND
+ VGND VPWR VPWR _06859_ sky130_fd_sc_hd__or4_2
X_19060_ net802 _02580_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_12504_ _07939_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16272_ CPU.registerFile\[28\]\[6\] CPU.registerFile\[29\]\[6\] _03739_ VGND VGND
+ VPWR VPWR _03993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13484_ _08433_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__buf_1
X_10696_ _06820_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18011_ net1022 _01539_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_15223_ CPU.registerFile\[19\]\[22\] CPU.registerFile\[18\]\[22\] _03157_ VGND VGND
+ VPWR VPWR _03283_ sky130_fd_sc_hd__mux2_1
X_12435_ net2006 _07347_ _07895_ VGND VGND VPWR VPWR _07903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15154_ _03049_ _03050_ CPU.registerFile\[25\]\[20\] VGND VGND VPWR VPWR _03216_
+ sky130_fd_sc_hd__a21o_1
X_12366_ _07866_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11317_ net2500 _06145_ _07249_ VGND VGND VPWR VPWR _07254_ sky130_fd_sc_hd__mux2_1
X_15085_ CPU.registerFile\[0\]\[18\] _02948_ _03148_ _02791_ VGND VGND VPWR VPWR _03149_
+ sky130_fd_sc_hd__o211a_1
X_15696__491 clknet_1_1__leaf__03647_ VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__inv_2
X_17338__750 clknet_1_1__leaf__04983_ VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__inv_2
XFILLER_0_10_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12297_ mapped_spi_ram.rcv_data\[2\] _07813_ VGND VGND VPWR VPWR _07824_ sky130_fd_sc_hd__or2_1
X_18913_ net687 _02433_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11248_ _06626_ net1892 _07212_ VGND VGND VPWR VPWR _07217_ sky130_fd_sc_hd__mux2_1
X_18844_ clknet_leaf_7_clk net1527 VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11179_ net2194 _07134_ VGND VGND VPWR VPWR _07173_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18775_ net564 _02299_ VGND VGND VPWR VPWR CPU.aluReg\[5\] sky130_fd_sc_hd__dfxtp_1
X_15987_ _03713_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__buf_4
XFILLER_0_54_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17726_ net811 _01292_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_14938_ _03003_ _03004_ _02851_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17657_ net1453 _05189_ _05192_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__o21ai_1
X_14869_ _02934_ _02936_ _02937_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__mux2_1
X_13533__923 clknet_1_0__leaf__08438_ VGND VGND VPWR VPWR net979 sky130_fd_sc_hd__inv_2
XFILLER_0_9_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16608_ CPU.registerFile\[24\]\[14\] _04319_ _04165_ _04320_ VGND VGND VPWR VPWR
+ _04321_ sky130_fd_sc_hd__o211a_1
X_17588_ _05120_ _05133_ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__nand2_1
X_16539_ CPU.registerFile\[16\]\[12\] _04252_ _04090_ _04253_ VGND VGND VPWR VPWR
+ _04254_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09011_ CPU.aluIn1\[20\] _05362_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__and2_1
X_18209_ net1220 _01737_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19189_ clknet_leaf_3_clk _02707_ VGND VGND VPWR VPWR per_uart.d_in_uart\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold101 mapped_spi_flash.rcv_data\[31\] VGND VGND VPWR VPWR net1398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 mapped_spi_flash.rcv_data\[7\] VGND VGND VPWR VPWR net1409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _08232_ VGND VGND VPWR VPWR net1420 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold134 mapped_spi_ram.rcv_data\[27\] VGND VGND VPWR VPWR net1431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _05837_ VGND VGND VPWR VPWR net1442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 per_uart.uart0.rx_count16\[3\] VGND VGND VPWR VPWR net1453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold167 _02674_ VGND VGND VPWR VPWR net1464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 _02676_ VGND VGND VPWR VPWR net1475 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _06246_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__clkbuf_1
Xhold189 mapped_spi_ram.rcv_data\[11\] VGND VGND VPWR VPWR net1486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09844_ _05466_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__inv_2
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ _06017_ _06113_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__nand2_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13755__1123 clknet_1_0__leaf__08460_ VGND VGND VPWR VPWR net1179 sky130_fd_sc_hd__inv_2
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10550_ net2079 _05767_ _06739_ VGND VGND VPWR VPWR _06741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14103__247 clknet_1_1__leaf__08494_ VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__inv_2
X_09209_ CPU.aluIn1\[19\] _05544_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__nand2_1
X_10481_ net1889 _05767_ _06702_ VGND VGND VPWR VPWR _06704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12220_ _07776_ _07777_ mapped_spi_ram.snd_bitcount\[1\] VGND VGND VPWR VPWR _07778_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12151_ mapped_spi_ram.cmd_addr\[14\] _07073_ _07724_ VGND VGND VPWR VPWR _07729_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11102_ net1433 mapped_spi_flash.rcv_bitcount\[1\] mapped_spi_flash.rcv_bitcount\[0\]
+ VGND VGND VPWR VPWR _07126_ sky130_fd_sc_hd__or3_1
X_12082_ CPU.mem_rstrb _05858_ VGND VGND VPWR VPWR _07680_ sky130_fd_sc_hd__nand2_1
Xhold690 CPU.registerFile\[30\]\[13\] VGND VGND VPWR VPWR net1987 sky130_fd_sc_hd__dlygate4sd3_1
X_15910_ clknet_1_0__leaf__08339_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__buf_1
X_11033_ CPU.PC\[9\] _07031_ _07071_ _07072_ _05703_ VGND VGND VPWR VPWR _07073_ sky130_fd_sc_hd__o221a_1
X_16890_ CPU.registerFile\[6\]\[21\] CPU.registerFile\[7\]\[21\] _04426_ VGND VGND
+ VPWR VPWR _04596_ sky130_fd_sc_hd__mux2_1
X_18560_ net381 _02084_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_12984_ _08195_ VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__clkbuf_1
X_17511_ _08335_ _06159_ _05073_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__o21ai_1
X_14723_ _02750_ _02775_ _02795_ _08597_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__a211o_1
X_11935_ _07597_ VGND VGND VPWR VPWR _07598_ sky130_fd_sc_hd__buf_4
X_18491_ net312 _02015_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14654_ _08532_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__clkbuf_4
X_17442_ _08379_ _05017_ _06451_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__o21bai_1
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _06663_ _06814_ VGND VGND VPWR VPWR _07561_ sky130_fd_sc_hd__nand2_2
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10817_ net2660 _06901_ _06889_ VGND VGND VPWR VPWR _06902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14585_ _08823_ _08824_ _08783_ VGND VGND VPWR VPWR _08825_ sky130_fd_sc_hd__mux2_1
X_17373_ per_uart.uart0.rxd_reg\[5\] _04992_ _04993_ per_uart.uart0.rxd_reg\[4\] VGND
+ VGND VPWR VPWR _05001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11797_ _07524_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__clkbuf_1
X_19112_ net95 _02632_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_16324_ CPU.registerFile\[22\]\[7\] CPU.registerFile\[23\]\[7\] _03958_ VGND VGND
+ VPWR VPWR _04044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10748_ _06847_ VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16255_ _03697_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__buf_2
X_19043_ net785 _02563_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13467_ _08424_ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__clkbuf_1
X_10679_ _06809_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15206_ _03138_ _03139_ CPU.registerFile\[9\]\[21\] VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__a21o_1
X_14078__224 clknet_1_1__leaf__08492_ VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__inv_2
X_12418_ net1758 _07330_ _07884_ VGND VGND VPWR VPWR _07894_ sky130_fd_sc_hd__mux2_1
X_16186_ _03901_ _03904_ _03908_ _03732_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__o211a_1
X_13398_ _08377_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15137_ _03155_ _03179_ _03199_ _02839_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__a211o_1
XFILLER_0_140_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12349_ _07857_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__clkbuf_1
X_13815__1177 clknet_1_0__leaf__08466_ VGND VGND VPWR VPWR net1233 sky130_fd_sc_hd__inv_2
X_15068_ _02798_ _03119_ _03123_ _03131_ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__a31o_1
X_18827_ net616 _02351_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09560_ _05374_ _05903_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__xnor2_2
X_18758_ net547 _02282_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[20\] sky130_fd_sc_hd__dfxtp_1
X_17709_ _05230_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__clkbuf_1
X_09491_ CPU.Bimm\[6\] _05758_ _05759_ CPU.cycles\[26\] net1442 VGND VGND VPWR VPWR
+ _05838_ sky130_fd_sc_hd__a221o_4
X_18689_ net478 _02213_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13314__814 clknet_1_0__leaf__08363_ VGND VGND VPWR VPWR net870 sky130_fd_sc_hd__inv_2
XFILLER_0_129_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09827_ _05343_ _05522_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__nor2_1
X_09758_ _06017_ _06092_ _06097_ _05800_ VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__a211o_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _06031_ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__clkbuf_4
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _07483_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__clkbuf_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11651_ _07446_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10602_ net1978 _06440_ _06761_ VGND VGND VPWR VPWR _06768_ sky130_fd_sc_hd__mux2_1
X_14027__178 clknet_1_1__leaf__08487_ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__inv_2
X_14370_ _08535_ _08610_ _08614_ _08554_ VGND VGND VPWR VPWR _08615_ sky130_fd_sc_hd__o211a_1
X_11582_ _07409_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_691 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10533_ net2527 _06440_ _06724_ VGND VGND VPWR VPWR _06731_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16040_ _03744_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__buf_4
XFILLER_0_135_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10464_ _06651_ net2309 _06687_ VGND VGND VPWR VPWR _06694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12203_ _07694_ _07759_ _07764_ VGND VGND VPWR VPWR _07765_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13183_ _08301_ net1607 VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10395_ _06485_ VGND VGND VPWR VPWR _06655_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12134_ net1404 _07714_ _07717_ _07713_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17991_ net1002 _01519_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12065_ CPU.registerFile\[24\]\[2\] _07372_ _07657_ VGND VGND VPWR VPWR _07667_ sky130_fd_sc_hd__mux2_1
X_16942_ CPU.registerFile\[27\]\[22\] CPU.registerFile\[26\]\[22\] _04646_ VGND VGND
+ VPWR VPWR _04647_ sky130_fd_sc_hd__mux2_1
X_15615__418 clknet_1_0__leaf__03639_ VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__inv_2
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11016_ _05595_ _05596_ _05597_ _07057_ VGND VGND VPWR VPWR _07058_ sky130_fd_sc_hd__o22a_1
X_16873_ _03750_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__clkbuf_4
X_18612_ net433 _02136_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18543_ net364 _02067_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_12967_ _08186_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14706_ _08525_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__buf_4
X_11918_ _06647_ net2421 _07584_ VGND VGND VPWR VPWR _07589_ sky130_fd_sc_hd__mux2_1
X_18474_ net295 _01998_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12898_ _05825_ net2120 _08145_ VGND VGND VPWR VPWR _08150_ sky130_fd_sc_hd__mux2_1
X_15686_ clknet_1_0__leaf__03643_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__buf_1
XFILLER_0_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11849_ _07552_ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14637_ CPU.registerFile\[19\]\[8\] CPU.registerFile\[18\]\[8\] _06064_ VGND VGND
+ VPWR VPWR _08875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14568_ _06058_ VGND VGND VPWR VPWR _08808_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17356_ per_uart.uart0.rx_count16\[1\] per_uart.uart0.rx_count16\[0\] VGND VGND VPWR
+ VPWR _04987_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16307_ _06172_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14499_ CPU.registerFile\[6\]\[4\] CPU.registerFile\[7\]\[4\] _08740_ VGND VGND VPWR
+ VPWR _08741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13754__1122 clknet_1_0__leaf__08460_ VGND VGND VPWR VPWR net1178 sky130_fd_sc_hd__inv_2
XFILLER_0_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19026_ net768 _02546_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[11\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__08452_ clknet_0__08452_ VGND VGND VPWR VPWR clknet_1_1__leaf__08452_
+ sky130_fd_sc_hd__clkbuf_16
X_16238_ CPU.registerFile\[20\]\[5\] CPU.registerFile\[21\]\[5\] _03883_ VGND VGND
+ VPWR VPWR _03960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__08483_ _08483_ VGND VGND VPWR VPWR clknet_0__08483_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16169_ CPU.aluIn1\[3\] _03566_ _03892_ _03855_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08991_ _05342_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__clkbuf_2
X_09612_ _05953_ _05954_ CPU.PC\[2\] VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__a21boi_1
X_13989__144 clknet_1_0__leaf__08483_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__inv_2
X_09543_ CPU.PC\[11\] _05886_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09474_ mapped_spi_ram.rcv_data\[3\] _05685_ _05698_ net1338 VGND VGND VPWR VPWR
+ _05822_ sky130_fd_sc_hd__a22o_2
XFILLER_0_149_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_634 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10180_ _05282_ _05522_ _05748_ VGND VGND VPWR VPWR _06503_ sky130_fd_sc_hd__o21ai_1
X_14215__348 clknet_1_1__leaf__08505_ VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__inv_2
X_13284__787 clknet_1_0__leaf__08345_ VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__inv_2
XFILLER_0_100_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__08472_ clknet_0__08472_ VGND VGND VPWR VPWR clknet_1_0__leaf__08472_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12821_ _08108_ VGND VGND VPWR VPWR _08109_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15540_ CPU.registerFile\[6\]\[30\] CPU.registerFile\[7\]\[30\] _08536_ VGND VGND
+ VPWR VPWR _03592_ sky130_fd_sc_hd__mux2_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ _08071_ VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__clkbuf_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _07474_ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__clkbuf_1
X_13814__1176 clknet_1_1__leaf__08466_ VGND VGND VPWR VPWR net1232 sky130_fd_sc_hd__inv_2
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15471_ _03235_ _03236_ CPU.registerFile\[1\]\[28\] VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _06607_ net2579 _08029_ VGND VGND VPWR VPWR _08035_ sky130_fd_sc_hd__mux2_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _08664_ _08665_ _08578_ VGND VGND VPWR VPWR _08666_ sky130_fd_sc_hd__mux2_1
X_17210_ _04545_ _04890_ _04907_ _08596_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__a211o_2
XFILLER_0_126_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11634_ _07437_ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18190_ net1201 net1436 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17141_ CPU.registerFile\[9\]\[28\] _03709_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__or2_1
X_14353_ CPU.mem_wdata\[0\] _08514_ _08598_ _07822_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__o211a_1
X_11565_ _07400_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17072_ CPU.registerFile\[15\]\[26\] CPU.registerFile\[14\]\[26\] _04550_ VGND VGND
+ VPWR VPWR _04773_ sky130_fd_sc_hd__mux2_1
X_10516_ net2486 _06245_ _06713_ VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__mux2_1
X_14284_ _06036_ VGND VGND VPWR VPWR _08530_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11496_ _06360_ VGND VGND VPWR VPWR _07360_ sky130_fd_sc_hd__buf_4
X_16023_ _05690_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__clkbuf_8
X_10447_ _06634_ net2192 _06676_ VGND VGND VPWR VPWR _06685_ sky130_fd_sc_hd__mux2_1
X_13166_ net1629 _08291_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__xor2_1
X_10378_ _06643_ net1958 _06639_ VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__mux2_1
X_12117_ mapped_spi_ram.cmd_addr\[24\] _07704_ _07695_ VGND VGND VPWR VPWR _07705_
+ sky130_fd_sc_hd__or3_1
X_17974_ net985 _01502_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_13097_ net1573 _08253_ _08254_ _08256_ _05237_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__a221o_1
X_16925_ CPU.registerFile\[13\]\[22\] _04380_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12048_ _07658_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16856_ _04305_ _04558_ _04562_ _04476_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__o211a_1
X_15807_ net1587 _08354_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__nand2_1
X_16787_ CPU.registerFile\[16\]\[18\] _04252_ _04494_ _04495_ VGND VGND VPWR VPWR
+ _04496_ sky130_fd_sc_hd__o211a_1
X_18526_ net347 _02050_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_887 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18457_ net278 _01985_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09190_ _05519_ _05524_ _05529_ _05537_ _05541_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__o41a_1
X_18388_ net209 _01916_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13569__955 clknet_1_0__leaf__08442_ VGND VGND VPWR VPWR net1011 sky130_fd_sc_hd__inv_2
XFILLER_0_83_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08504_ clknet_0__08504_ VGND VGND VPWR VPWR clknet_1_1__leaf__08504_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19009_ clknet_leaf_11_clk _02529_ VGND VGND VPWR VPWR CPU.aluIn1\[26\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__08435_ clknet_0__08435_ VGND VGND VPWR VPWR clknet_1_1__leaf__08435_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__08466_ _08466_ VGND VGND VPWR VPWR clknet_0__08466_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__08366_ clknet_0__08366_ VGND VGND VPWR VPWR clknet_1_1__leaf__08366_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08974_ CPU.aluIn1\[15\] _05325_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__and2_1
Xhold16 _01723_ VGND VGND VPWR VPWR net1313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 mapped_spi_ram.snd_bitcount\[0\] VGND VGND VPWR VPWR net1324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 CPU.aluReg\[17\] VGND VGND VPWR VPWR net1335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 mapped_spi_flash.rcv_data\[6\] VGND VGND VPWR VPWR net1346 sky130_fd_sc_hd__dlygate4sd3_1
X_09526_ CPU.Iimm\[4\] _05758_ _05759_ CPU.cycles\[24\] _05870_ VGND VGND VPWR VPWR
+ _05871_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09457_ net2478 _05805_ _05742_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15644__444 clknet_1_0__leaf__03642_ VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__inv_2
XFILLER_0_35_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09388_ _05737_ _05738_ CPU.writeBack _05739_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_19_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14221__352 clknet_1_1__leaf__08507_ VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__inv_2
XFILLER_0_22_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11350_ net1933 _06530_ _07237_ VGND VGND VPWR VPWR _07271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10301_ net1789 _06530_ _06557_ VGND VGND VPWR VPWR _06591_ sky130_fd_sc_hd__mux2_1
X_11281_ _06659_ net2434 _07200_ VGND VGND VPWR VPWR _07234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13020_ net1677 _07374_ _08180_ VGND VGND VPWR VPWR _08214_ sky130_fd_sc_hd__mux2_1
X_14139__279 clknet_1_1__leaf__08498_ VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__inv_2
X_10232_ _06547_ _06552_ _05541_ VGND VGND VPWR VPWR _06553_ sky130_fd_sc_hd__o21a_1
X_10163_ net2301 _06486_ _06293_ VGND VGND VPWR VPWR _06487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10094_ _06392_ _06416_ _06419_ _05556_ VGND VGND VPWR VPWR _06420_ sky130_fd_sc_hd__a22o_1
X_14971_ CPU.registerFile\[17\]\[16\] _03036_ VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__or2_1
X_13894__58 clknet_1_1__leaf__08474_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__inv_2
X_16710_ CPU.registerFile\[15\]\[17\] CPU.registerFile\[14\]\[17\] _04146_ VGND VGND
+ VPWR VPWR _04420_ sky130_fd_sc_hd__mux2_1
X_17690_ _05217_ VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16641_ _04098_ _04339_ _04343_ _04352_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__a31o_2
X_13853_ clknet_1_1__leaf__08462_ VGND VGND VPWR VPWR _08470_ sky130_fd_sc_hd__buf_1
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__08455_ clknet_0__08455_ VGND VGND VPWR VPWR clknet_1_0__leaf__08455_
+ sky130_fd_sc_hd__clkbuf_16
X_12804_ _08098_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__clkbuf_1
X_15727__519 clknet_1_1__leaf__03650_ VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__inv_2
X_16572_ CPU.registerFile\[22\]\[13\] CPU.registerFile\[23\]\[13\] _03958_ VGND VGND
+ VPWR VPWR _04286_ sky130_fd_sc_hd__mux2_1
X_10996_ _07008_ _07040_ VGND VGND VPWR VPWR _07041_ sky130_fd_sc_hd__or2_1
X_18311_ net132 _01839_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15523_ CPU.registerFile\[30\]\[30\] CPU.registerFile\[31\]\[30\] _03291_ VGND VGND
+ VPWR VPWR _03575_ sky130_fd_sc_hd__mux2_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _06659_ net2598 _08028_ VGND VGND VPWR VPWR _08062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ net1253 _01770_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__04980_ _04980_ VGND VGND VPWR VPWR clknet_0__04980_ sky130_fd_sc_hd__clkbuf_16
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15454_ _08566_ _08568_ CPU.registerFile\[25\]\[28\] VGND VGND VPWR VPWR _03508_
+ sky130_fd_sc_hd__a21o_1
X_12666_ _08025_ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11617_ net2237 _07335_ _07427_ VGND VGND VPWR VPWR _07429_ sky130_fd_sc_hd__mux2_1
X_14405_ CPU.registerFile\[27\]\[2\] CPU.registerFile\[26\]\[2\] _06063_ VGND VGND
+ VPWR VPWR _08649_ sky130_fd_sc_hd__mux2_1
X_18173_ net1184 _01701_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[12\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_142_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12597_ CPU.registerFile\[12\]\[2\] _07372_ _07979_ VGND VGND VPWR VPWR _07989_ sky130_fd_sc_hd__mux2_1
X_15385_ _06013_ _03436_ _03440_ _03092_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17124_ CPU.registerFile\[27\]\[27\] CPU.registerFile\[26\]\[27\] _04646_ VGND VGND
+ VPWR VPWR _04824_ sky130_fd_sc_hd__mux2_1
X_11548_ net1739 _07335_ _07390_ VGND VGND VPWR VPWR _07392_ sky130_fd_sc_hd__mux2_1
X_14336_ _08525_ VGND VGND VPWR VPWR _08582_ sky130_fd_sc_hd__buf_4
XFILLER_0_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold508 CPU.registerFile\[19\]\[15\] VGND VGND VPWR VPWR net1805 sky130_fd_sc_hd__dlygate4sd3_1
X_17055_ _04441_ _04754_ _04756_ _04612_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__a211o_1
X_14267_ _08512_ VGND VGND VPWR VPWR _08513_ sky130_fd_sc_hd__buf_4
Xhold519 CPU.registerFile\[20\]\[18\] VGND VGND VPWR VPWR net1816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11479_ _07348_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16006_ _03716_ _03721_ _03731_ _03732_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__o211a_1
X_13218_ _08311_ _05880_ _08331_ CPU.state\[1\] VGND VGND VPWR VPWR _08332_ sky130_fd_sc_hd__o31a_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13149_ CPU.cycles\[12\] _08281_ VGND VGND VPWR VPWR _08283_ sky130_fd_sc_hd__and2_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ net968 _01485_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xhold1208 CPU.registerFile\[2\]\[3\] VGND VGND VPWR VPWR net2505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 CPU.registerFile\[1\]\[29\] VGND VGND VPWR VPWR net2516 sky130_fd_sc_hd__dlygate4sd3_1
X_16908_ _04479_ _04608_ _04613_ _04446_ VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__o211a_1
X_17888_ clknet_leaf_23_clk net1503 VGND VGND VPWR VPWR CPU.cycles\[31\] sky130_fd_sc_hd__dfxtp_1
X_16839_ CPU.registerFile\[10\]\[20\] CPU.registerFile\[11\]\[20\] _04335_ VGND VGND
+ VPWR VPWR _04546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09311_ _05558_ _05661_ _05662_ _05235_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__o211a_2
X_18509_ net330 _02033_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17394__18 clknet_1_1__leaf__04985_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__inv_2
XFILLER_0_146_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09242_ _05570_ _05592_ _05593_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09173_ CPU.rs2\[31\] _05247_ _05251_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__o21a_1
XFILLER_0_145_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13675__1051 clknet_1_0__leaf__08452_ VGND VGND VPWR VPWR net1107 sky130_fd_sc_hd__inv_2
XFILLER_0_4_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__08449_ _08449_ VGND VGND VPWR VPWR clknet_0__08449_ sky130_fd_sc_hd__clkbuf_16
X_13813__1175 clknet_1_1__leaf__08466_ VGND VGND VPWR VPWR net1231 sky130_fd_sc_hd__inv_2
X_08957_ CPU.aluIn1\[10\] _05260_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__nor2_1
X_08888_ CPU.instr\[6\] CPU.instr\[4\] CPU.instr\[5\] VGND VGND VPWR VPWR _05240_
+ sky130_fd_sc_hd__nand3b_4
X_10850_ CPU.aluReg\[15\] CPU.aluReg\[13\] _06906_ VGND VGND VPWR VPWR _06927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09509_ _05854_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__clkbuf_1
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10781_ CPU.aluIn1\[30\] _06873_ _06861_ VGND VGND VPWR VPWR _06874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12520_ net1829 _07364_ _07942_ VGND VGND VPWR VPWR _07948_ sky130_fd_sc_hd__mux2_1
X_18582__39 VGND VGND VPWR VPWR _18582__39/HI net39 sky130_fd_sc_hd__conb_1
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ _07911_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11402_ net2155 _06337_ _07296_ VGND VGND VPWR VPWR _07299_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15170_ CPU.registerFile\[5\]\[20\] CPU.registerFile\[4\]\[20\] _03105_ VGND VGND
+ VPWR VPWR _03232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12382_ _06647_ net1769 _07870_ VGND VGND VPWR VPWR _07875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11333_ _07262_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11264_ _07225_ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__clkbuf_1
X_14072__219 clknet_1_1__leaf__08491_ VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__inv_2
X_13003_ _08205_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__clkbuf_1
X_10215_ _06535_ _06204_ VGND VGND VPWR VPWR _06536_ sky130_fd_sc_hd__nand2_1
X_18860_ net634 _02380_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_11195_ _07185_ VGND VGND VPWR VPWR _07186_ sky130_fd_sc_hd__inv_2
X_17811_ net891 _01373_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_10146_ CPU.cycles\[3\] _05553_ _06368_ _06467_ _06469_ VGND VGND VPWR VPWR _06470_
+ sky130_fd_sc_hd__a221o_1
X_18791_ net580 _02315_ VGND VGND VPWR VPWR CPU.aluReg\[21\] sky130_fd_sc_hd__dfxtp_1
X_17742_ net827 _01308_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_14954_ _08857_ _03017_ _03020_ _02903_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__a211o_1
X_10077_ _05300_ _05430_ _05446_ VGND VGND VPWR VPWR _06404_ sky130_fd_sc_hd__nand3_1
XFILLER_0_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17673_ net1639 _05203_ _05204_ _05192_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_0__f__08507_ clknet_0__08507_ VGND VGND VPWR VPWR clknet_1_0__leaf__08507_
+ sky130_fd_sc_hd__clkbuf_16
X_14885_ _02750_ _02933_ _02953_ _02839_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__a211o_1
XFILLER_0_159_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16624_ CPU.registerFile\[10\]\[15\] CPU.registerFile\[11\]\[15\] _04335_ VGND VGND
+ VPWR VPWR _04336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__08438_ clknet_0__08438_ VGND VGND VPWR VPWR clknet_1_0__leaf__08438_
+ sky130_fd_sc_hd__clkbuf_16
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16555_ CPU.registerFile\[5\]\[13\] CPU.registerFile\[4\]\[13\] _04024_ VGND VGND
+ VPWR VPWR _04269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10979_ _05567_ _05569_ _05594_ VGND VGND VPWR VPWR _07025_ sky130_fd_sc_hd__and3_1
Xclkbuf_1_0__f__08369_ clknet_0__08369_ VGND VGND VPWR VPWR clknet_1_0__leaf__08369_
+ sky130_fd_sc_hd__clkbuf_16
X_15506_ CPU.registerFile\[2\]\[29\] CPU.registerFile\[3\]\[29\] _03275_ VGND VGND
+ VPWR VPWR _03559_ sky130_fd_sc_hd__mux2_1
X_12718_ _08053_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__clkbuf_1
X_16486_ CPU.registerFile\[30\]\[11\] CPU.registerFile\[31\]\[11\] _04201_ VGND VGND
+ VPWR VPWR _04202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13698_ clknet_1_1__leaf__08451_ VGND VGND VPWR VPWR _08455_ sky130_fd_sc_hd__buf_1
XFILLER_0_150_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18225_ net1236 _01753_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[26\] sky130_fd_sc_hd__dfxtp_1
X_15437_ _08414_ _03489_ _03491_ _08419_ VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__a211o_1
XFILLER_0_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12649_ _06641_ net2046 _08015_ VGND VGND VPWR VPWR _08017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18156_ net1167 net1305 VGND VGND VPWR VPWR mapped_spi_ram.rcv_bitcount\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15368_ _03155_ _03407_ _03424_ _03243_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__a211o_2
XFILLER_0_108_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17107_ _04503_ _04804_ _04806_ _04509_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__a211o_1
X_14319_ CPU.registerFile\[10\]\[0\] CPU.registerFile\[11\]\[0\] _08564_ VGND VGND
+ VPWR VPWR _08565_ sky130_fd_sc_hd__mux2_1
Xhold305 mapped_spi_flash.rcv_data\[21\] VGND VGND VPWR VPWR net1602 sky130_fd_sc_hd__dlygate4sd3_1
X_18087_ net1098 _01615_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xhold316 CPU.cycles\[10\] VGND VGND VPWR VPWR net1613 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15299_ CPU.registerFile\[16\]\[24\] _03159_ _03356_ _03161_ VGND VGND VPWR VPWR
+ _03357_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold327 per_uart.uart0.enable16_counter\[11\] VGND VGND VPWR VPWR net1624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 CPU.registerFile\[13\]\[30\] VGND VGND VPWR VPWR net1635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17038_ CPU.registerFile\[12\]\[25\] _04421_ _04422_ _04739_ VGND VGND VPWR VPWR
+ _04740_ sky130_fd_sc_hd__o211a_1
Xhold349 CPU.rs2\[16\] VGND VGND VPWR VPWR net1646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09860_ CPU.PC\[15\] _05889_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__xnor2_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15673__470 clknet_1_0__leaf__03645_ VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__inv_2
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _06126_ _06128_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__nand2_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ clknet_leaf_18_clk _02509_ VGND VGND VPWR VPWR CPU.aluIn1\[6\] sky130_fd_sc_hd__dfxtp_4
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 CPU.registerFile\[9\]\[29\] VGND VGND VPWR VPWR net2302 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1016 CPU.registerFile\[9\]\[21\] VGND VGND VPWR VPWR net2313 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1027 CPU.registerFile\[29\]\[16\] VGND VGND VPWR VPWR net2324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 CPU.registerFile\[7\]\[12\] VGND VGND VPWR VPWR net2335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 CPU.registerFile\[11\]\[31\] VGND VGND VPWR VPWR net2346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13510__902 clknet_1_0__leaf__08436_ VGND VGND VPWR VPWR net958 sky130_fd_sc_hd__inv_2
XFILLER_0_91_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09225_ CPU.aluIn1\[0\] _05576_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__nand2_8
XFILLER_0_63_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09156_ _05254_ CPU.aluIn1\[29\] VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__and2b_1
XFILLER_0_115_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09087_ _05436_ _05274_ _05438_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__a21o_1
X_15756__545 clknet_1_0__leaf__03653_ VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__inv_2
Xhold850 CPU.registerFile\[10\]\[1\] VGND VGND VPWR VPWR net2147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 CPU.registerFile\[31\]\[20\] VGND VGND VPWR VPWR net2158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold872 CPU.registerFile\[22\]\[30\] VGND VGND VPWR VPWR net2169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 CPU.registerFile\[18\]\[12\] VGND VGND VPWR VPWR net2180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 CPU.registerFile\[12\]\[22\] VGND VGND VPWR VPWR net2191 sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ CPU.cycles\[9\] _05553_ _06197_ _06329_ VGND VGND VPWR VPWR _06330_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_101_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09989_ _06272_ _06318_ VGND VGND VPWR VPWR _06319_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11951_ _07606_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__clkbuf_1
X_10902_ _06966_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__clkbuf_1
X_14670_ CPU.registerFile\[0\]\[8\] _08706_ _02743_ _08588_ VGND VGND VPWR VPWR _02744_
+ sky130_fd_sc_hd__o211a_1
X_11882_ _06611_ net1853 _07562_ VGND VGND VPWR VPWR _07570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10833_ _06880_ VGND VGND VPWR VPWR _06914_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16340_ _08398_ _04055_ _04058_ _08401_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__a211o_1
XFILLER_0_149_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10764_ _06857_ _06851_ net1653 _06858_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__o211ai_1
X_12503_ net2247 _07347_ _07931_ VGND VGND VPWR VPWR _07939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13483_ _05545_ _05687_ _08265_ VGND VGND VPWR VPWR _08433_ sky130_fd_sc_hd__mux2_1
X_16271_ CPU.registerFile\[30\]\[6\] CPU.registerFile\[31\]\[6\] _03796_ VGND VGND
+ VPWR VPWR _03992_ sky130_fd_sc_hd__mux2_1
X_10695_ net1895 _05805_ _06816_ VGND VGND VPWR VPWR _06820_ sky130_fd_sc_hd__mux2_1
X_18010_ net1021 _01538_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_12434_ _07902_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__clkbuf_1
X_15222_ net1657 _03201_ _03282_ _02993_ VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12365_ _06630_ net2149 _07859_ VGND VGND VPWR VPWR _07866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15153_ CPU.registerFile\[27\]\[20\] CPU.registerFile\[26\]\[20\] _03172_ VGND VGND
+ VPWR VPWR _03215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11316_ _07253_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15084_ _02831_ _02832_ CPU.registerFile\[1\]\[18\] VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__a21o_1
X_12296_ net1484 _07812_ _07823_ _07822_ VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__o211a_1
X_18912_ net686 _02432_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11247_ _07216_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__clkbuf_1
X_18843_ clknet_leaf_8_clk _02367_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11178_ net1640 _07160_ _07172_ _07164_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__o211a_1
X_10129_ CPU.cycles\[4\] _05552_ _06197_ _06453_ VGND VGND VPWR VPWR _06454_ sky130_fd_sc_hd__o2bb2a_1
X_18774_ net563 _02298_ VGND VGND VPWR VPWR CPU.aluReg\[4\] sky130_fd_sc_hd__dfxtp_1
X_15986_ _03712_ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__clkbuf_8
X_15885__629 clknet_1_0__leaf__03683_ VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__inv_2
X_17725_ net810 _01291_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_14937_ CPU.registerFile\[28\]\[15\] CPU.registerFile\[29\]\[15\] _02808_ VGND VGND
+ VPWR VPWR _03004_ sky130_fd_sc_hd__mux2_1
X_13379__872 clknet_1_1__leaf__08370_ VGND VGND VPWR VPWR net928 sky130_fd_sc_hd__inv_2
X_13674__1050 clknet_1_0__leaf__08452_ VGND VGND VPWR VPWR net1106 sky130_fd_sc_hd__inv_2
XFILLER_0_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17656_ _04986_ _05185_ _05236_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__a21oi_2
X_14868_ _08540_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__buf_4
X_16607_ _04080_ _04081_ CPU.registerFile\[25\]\[14\] VGND VGND VPWR VPWR _04320_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17587_ _05236_ _05120_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__nor2_1
X_14799_ _02868_ _02869_ _08783_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__mux2_1
X_13983__139 clknet_1_0__leaf__08482_ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__inv_2
XFILLER_0_161_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16538_ _04175_ _04176_ CPU.registerFile\[17\]\[12\] VGND VGND VPWR VPWR _04253_
+ sky130_fd_sc_hd__a21o_1
X_13812__1174 clknet_1_1__leaf__08466_ VGND VGND VPWR VPWR net1230 sky130_fd_sc_hd__inv_2
XFILLER_0_85_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16469_ CPU.registerFile\[9\]\[11\] _04056_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09010_ CPU.rs2\[20\] _05246_ _05250_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__o21a_1
X_18208_ net1219 _01736_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19188_ clknet_leaf_3_clk _02706_ VGND VGND VPWR VPWR per_uart.d_in_uart\[3\] sky130_fd_sc_hd__dfxtp_1
X_15705__499 clknet_1_1__leaf__03648_ VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__inv_2
XFILLER_0_54_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18139_ net1150 _01667_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold102 _06385_ VGND VGND VPWR VPWR net1399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold113 _05733_ VGND VGND VPWR VPWR net1410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 CPU.aluReg\[2\] VGND VGND VPWR VPWR net1421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _01717_ VGND VGND VPWR VPWR net1432 sky130_fd_sc_hd__dlygate4sd3_1
X_14055__203 clknet_1_0__leaf__08490_ VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__inv_2
XFILLER_0_13_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold146 _08223_ VGND VGND VPWR VPWR net1443 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 mapped_spi_ram.rcv_data\[7\] VGND VGND VPWR VPWR net1454 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold168 mapped_spi_ram.rcv_data\[8\] VGND VGND VPWR VPWR net1465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 per_uart.uart0.txd_reg\[4\] VGND VGND VPWR VPWR net1476 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ net2511 _06245_ _06055_ VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__mux2_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ CPU.Jimm\[15\] _05550_ _05553_ CPU.cycles\[15\] VGND VGND VPWR VPWR _06179_
+ sky130_fd_sc_hd__a22o_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _05357_ _06090_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__xnor2_2
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09208_ CPU.aluIn1\[21\] _05544_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10480_ _06703_ VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09139_ _05368_ CPU.aluIn1\[21\] VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__and2b_1
XFILLER_0_60_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12150_ net1495 _07714_ _07728_ _07713_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11101_ _07125_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__clkbuf_1
X_13248__769 clknet_1_1__leaf__08343_ VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__inv_2
X_12081_ _07679_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__clkbuf_1
Xhold680 CPU.registerFile\[18\]\[8\] VGND VGND VPWR VPWR net1977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold691 CPU.registerFile\[20\]\[30\] VGND VGND VPWR VPWR net1988 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ _05604_ _07070_ _07023_ VGND VGND VPWR VPWR _07072_ sky130_fd_sc_hd__a21o_1
X_12983_ net1673 _07337_ _08192_ VGND VGND VPWR VPWR _08195_ sky130_fd_sc_hd__mux2_1
X_17510_ _05084_ _05085_ _05058_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__a21oi_1
X_14722_ _02785_ _02794_ _08594_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__o21a_2
X_18490_ net311 _02014_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_11934_ _06595_ _06814_ VGND VGND VPWR VPWR _07597_ sky130_fd_sc_hd__nand2_2
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17441_ _05027_ _05028_ _05029_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__a21oi_1
X_14653_ _08515_ _08878_ _02718_ _02726_ VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__a31o_1
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11865_ _07560_ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__clkbuf_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03679_ clknet_0__03679_ VGND VGND VPWR VPWR clknet_1_0__leaf__03679_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10816_ CPU.aluIn1\[22\] _06900_ _06881_ VGND VGND VPWR VPWR _06901_ sky130_fd_sc_hd__mux2_1
X_17372_ _05000_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__clkbuf_1
X_14584_ CPU.registerFile\[5\]\[6\] CPU.registerFile\[4\]\[6\] _08576_ VGND VGND VPWR
+ VPWR _08824_ sky130_fd_sc_hd__mux2_1
X_11796_ _06661_ net2217 _07489_ VGND VGND VPWR VPWR _07524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19111_ net94 _02631_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16323_ _03735_ _04036_ _04041_ _04042_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10747_ net2244 _06486_ _06838_ VGND VGND VPWR VPWR _06847_ sky130_fd_sc_hd__mux2_1
X_19042_ net784 _02562_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16254_ CPU.registerFile\[15\]\[6\] CPU.registerFile\[14\]\[6\] _03705_ VGND VGND
+ VPWR VPWR _03975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10678_ CPU.registerFile\[1\]\[2\] _06508_ _06799_ VGND VGND VPWR VPWR _06809_ sky130_fd_sc_hd__mux2_1
X_13466_ CPU.Iimm\[3\] _08423_ _08416_ VGND VGND VPWR VPWR _08424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14004__157 clknet_1_1__leaf__08485_ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__inv_2
X_15205_ CPU.registerFile\[10\]\[21\] CPU.registerFile\[11\]\[21\] _03183_ VGND VGND
+ VPWR VPWR _03266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12417_ _07893_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16185_ _03722_ _03905_ _03907_ _03730_ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__a211o_1
X_13397_ _05538_ _05539_ _08371_ VGND VGND VPWR VPWR _08377_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15136_ _03189_ _03198_ _02837_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__o21a_2
XFILLER_0_140_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12348_ _06613_ net2168 _07848_ VGND VGND VPWR VPWR _07857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12279_ net1461 _07812_ _07814_ _07809_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__o211a_1
X_15067_ _02964_ _03126_ _03130_ _03092_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__o211a_1
X_18826_ net615 _02350_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_18757_ net546 _02281_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[19\] sky130_fd_sc_hd__dfxtp_1
X_15969_ _05689_ _05690_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__and2_1
X_14050__199 clknet_1_0__leaf__08489_ VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__inv_2
X_17708_ _05207_ _05229_ VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09490_ _05731_ _05828_ _05836_ _05541_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__a22o_1
X_18688_ net477 _02212_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17639_ per_uart.uart0.uart_rxd2 _05168_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09826_ _05340_ _05531_ _05534_ CPU.aluReg\[16\] _06162_ VGND VGND VPWR VPWR _06163_
+ sky130_fd_sc_hd__a221o_1
X_15868__613 clknet_1_0__leaf__03682_ VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__inv_2
X_09757_ _06017_ _06096_ VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__nor2_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _05764_ _06014_ _06027_ _06030_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__a211o_4
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13966__123 clknet_1_1__leaf__08481_ VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__inv_2
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11650_ net2028 _07368_ _07438_ VGND VGND VPWR VPWR _07446_ sky130_fd_sc_hd__mux2_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10601_ _06767_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__clkbuf_1
X_11581_ net1791 _07368_ _07401_ VGND VGND VPWR VPWR _07409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10532_ _06730_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10463_ _06693_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__clkbuf_1
X_13251_ clknet_1_1__leaf__08341_ VGND VGND VPWR VPWR _08344_ sky130_fd_sc_hd__buf_1
X_12202_ _07688_ _07763_ VGND VGND VPWR VPWR _07764_ sky130_fd_sc_hd__nand2_4
X_13182_ CPU.cycles\[25\] _08299_ net1606 VGND VGND VPWR VPWR _08302_ sky130_fd_sc_hd__a21oi_1
X_10394_ _06654_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12133_ _07715_ _07716_ VGND VGND VPWR VPWR _07717_ sky130_fd_sc_hd__or2_1
X_17990_ net1001 _01518_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16941_ _03744_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__buf_4
X_12064_ _07666_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__clkbuf_1
X_13811__1173 clknet_1_1__leaf__08466_ VGND VGND VPWR VPWR net1229 sky130_fd_sc_hd__inv_2
X_11015_ _05599_ _07056_ VGND VGND VPWR VPWR _07057_ sky130_fd_sc_hd__and2b_1
X_16872_ _03748_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__clkbuf_4
X_18611_ net432 _02135_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18542_ net363 _02066_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12966_ net2208 _07320_ _08181_ VGND VGND VPWR VPWR _08186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14705_ _02776_ _02777_ _08695_ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__mux2_1
X_18473_ net294 _01997_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_11917_ _07588_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__clkbuf_1
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _08149_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__clkbuf_1
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14636_ CPU.mem_wdata\[7\] _08514_ _08874_ _08751_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__o211a_1
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ net2626 _07360_ _07548_ VGND VGND VPWR VPWR _07552_ sky130_fd_sc_hd__mux2_1
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ per_uart.uart0.rx_busy VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__inv_2
X_14567_ CPU.registerFile\[27\]\[6\] CPU.registerFile\[26\]\[6\] _06063_ VGND VGND
+ VPWR VPWR _08807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11779_ _07515_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16306_ _04023_ _04025_ _03720_ VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14498_ _08525_ VGND VGND VPWR VPWR _08740_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19025_ net767 _02545_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08451_ clknet_0__08451_ VGND VGND VPWR VPWR clknet_1_1__leaf__08451_
+ sky130_fd_sc_hd__clkbuf_16
X_16237_ CPU.registerFile\[22\]\[5\] CPU.registerFile\[23\]\[5\] _03958_ VGND VGND
+ VPWR VPWR _03959_ sky130_fd_sc_hd__mux2_1
X_13449_ _08409_ VGND VGND VPWR VPWR _08410_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__08482_ _08482_ VGND VGND VPWR VPWR clknet_0__08482_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16168_ _03692_ _03872_ _03891_ _03601_ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__a211o_1
XFILLER_0_100_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15119_ _03180_ _03181_ _02937_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__mux2_1
X_08990_ _05340_ _05341_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__or2_1
X_16099_ CPU.registerFile\[6\]\[2\] CPU.registerFile\[7\]\[2\] _03717_ VGND VGND VPWR
+ VPWR _03824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09611_ CPU.PC\[2\] _05953_ _05954_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__nand3b_1
X_18809_ net598 _02333_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_14167__304 clknet_1_0__leaf__08501_ VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__inv_2
XFILLER_0_78_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09542_ CPU.PC\[10\] CPU.PC\[9\] _05885_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__and3_1
X_09473_ CPU.Bimm\[7\] _05758_ _05759_ CPU.cycles\[27\] VGND VGND VPWR VPWR _05821_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09809_ _06146_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__clkbuf_1
X_14033__183 clknet_1_0__leaf__08488_ VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__08471_ clknet_0__08471_ VGND VGND VPWR VPWR clknet_1_0__leaf__08471_
+ sky130_fd_sc_hd__clkbuf_16
X_12820_ _07488_ _07199_ VGND VGND VPWR VPWR _08108_ sky130_fd_sc_hd__nand2_4
X_13592__976 clknet_1_1__leaf__08444_ VGND VGND VPWR VPWR net1032 sky130_fd_sc_hd__inv_2
XFILLER_0_158_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _06607_ net2118 _08065_ VGND VGND VPWR VPWR _08071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ net2453 _07351_ _07464_ VGND VGND VPWR VPWR _07474_ sky130_fd_sc_hd__mux2_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ CPU.registerFile\[2\]\[28\] CPU.registerFile\[3\]\[28\] _03275_ VGND VGND
+ VPWR VPWR _03524_ sky130_fd_sc_hd__mux2_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _08034_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ CPU.registerFile\[5\]\[2\] CPU.registerFile\[4\]\[2\] _08576_ VGND VGND VPWR
+ VPWR _08665_ sky130_fd_sc_hd__mux2_1
X_11633_ net2335 _07351_ _07427_ VGND VGND VPWR VPWR _07437_ sky130_fd_sc_hd__mux2_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17140_ CPU.registerFile\[10\]\[28\] CPU.registerFile\[11\]\[28\] _06173_ VGND VGND
+ VPWR VPWR _04839_ sky130_fd_sc_hd__mux2_1
X_14352_ _08425_ _08556_ _08595_ _08597_ VGND VGND VPWR VPWR _08598_ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11564_ net1846 _07351_ _07390_ VGND VGND VPWR VPWR _07400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15621__423 clknet_1_1__leaf__03640_ VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__inv_2
XFILLER_0_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17071_ _04503_ _04769_ _04771_ _04509_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__a211o_1
XFILLER_0_80_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10515_ _06721_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__clkbuf_1
X_11495_ _07359_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__clkbuf_1
X_14283_ CPU.registerFile\[21\]\[0\] _08528_ VGND VGND VPWR VPWR _08529_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16022_ _03748_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__clkbuf_4
X_13486__881 clknet_1_0__leaf__08370_ VGND VGND VPWR VPWR net937 sky130_fd_sc_hd__inv_2
X_10446_ _06684_ VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10377_ _06336_ VGND VGND VPWR VPWR _06643_ sky130_fd_sc_hd__buf_4
X_13165_ _08291_ _08292_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__nor2_1
X_12116_ _07703_ VGND VGND VPWR VPWR _07704_ sky130_fd_sc_hd__buf_4
X_17973_ net984 _01501_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_13096_ _08255_ VGND VGND VPWR VPWR _08256_ sky130_fd_sc_hd__clkbuf_4
X_13343__841 clknet_1_1__leaf__08365_ VGND VGND VPWR VPWR net897 sky130_fd_sc_hd__inv_2
X_14116__258 clknet_1_1__leaf__08496_ VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__inv_2
X_16924_ CPU.registerFile\[15\]\[22\] CPU.registerFile\[14\]\[22\] _04550_ VGND VGND
+ VPWR VPWR _04629_ sky130_fd_sc_hd__mux2_1
X_12047_ CPU.registerFile\[24\]\[11\] _07353_ _07657_ VGND VGND VPWR VPWR _07658_
+ sky130_fd_sc_hd__mux2_1
X_16855_ _04347_ _04559_ _04561_ _04521_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__a211o_1
X_15806_ _08354_ _03671_ _03661_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18588__45 VGND VGND VPWR VPWR _18588__45/HI net45 sky130_fd_sc_hd__conb_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16786_ _04175_ _04176_ CPU.registerFile\[17\]\[18\] VGND VGND VPWR VPWR _04495_
+ sky130_fd_sc_hd__a21o_1
X_13998_ clknet_1_1__leaf__08484_ VGND VGND VPWR VPWR _08485_ sky130_fd_sc_hd__buf_1
X_18525_ net346 _02049_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12949_ _08176_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18456_ net277 _01984_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14619_ CPU.registerFile\[10\]\[7\] CPU.registerFile\[11\]\[7\] _08564_ VGND VGND
+ VPWR VPWR _08858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18387_ net208 _01915_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__08503_ clknet_0__08503_ VGND VGND VPWR VPWR clknet_1_1__leaf__08503_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17269_ _03726_ _03727_ CPU.registerFile\[25\]\[31\] VGND VGND VPWR VPWR _04965_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19008_ clknet_leaf_11_clk _02528_ VGND VGND VPWR VPWR CPU.aluIn1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__08434_ clknet_0__08434_ VGND VGND VPWR VPWR clknet_1_1__leaf__08434_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__08465_ _08465_ VGND VGND VPWR VPWR clknet_0__08465_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__08365_ clknet_0__08365_ VGND VGND VPWR VPWR clknet_1_1__leaf__08365_
+ sky130_fd_sc_hd__clkbuf_16
X_08973_ CPU.rs2\[15\] _05245_ _05249_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold17 mapped_spi_ram.cmd_addr\[1\] VGND VGND VPWR VPWR net1314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 mapped_spi_ram.cmd_addr\[26\] VGND VGND VPWR VPWR net1325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 _08233_ VGND VGND VPWR VPWR net1336 sky130_fd_sc_hd__dlygate4sd3_1
X_17284__701 clknet_1_1__leaf__03691_ VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__inv_2
X_09525_ _05866_ _05868_ _05869_ _05744_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__o31a_1
XFILLER_0_148_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09456_ _05804_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09387_ CPU.Bimm\[4\] VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13810__1172 clknet_1_1__leaf__08466_ VGND VGND VPWR VPWR net1228 sky130_fd_sc_hd__inv_2
X_13290__792 clknet_1_0__leaf__08361_ VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__inv_2
XFILLER_0_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10300_ _06590_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__clkbuf_1
X_11280_ _07233_ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__clkbuf_1
X_10231_ _06548_ _05533_ _05536_ net1617 _06551_ VGND VGND VPWR VPWR _06552_ sky130_fd_sc_hd__a221o_1
X_10162_ _06485_ VGND VGND VPWR VPWR _06486_ sky130_fd_sc_hd__clkbuf_4
X_10093_ _06241_ _06393_ _06417_ _06395_ _06418_ VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__a32o_1
X_14970_ _06062_ VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__buf_2
X_13600__983 clknet_1_0__leaf__08445_ VGND VGND VPWR VPWR net1039 sky130_fd_sc_hd__inv_2
X_16640_ _04305_ _04346_ _04351_ _04072_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__08454_ clknet_0__08454_ VGND VGND VPWR VPWR clknet_1_0__leaf__08454_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12803_ _06659_ net2602 _08064_ VGND VGND VPWR VPWR _08098_ sky130_fd_sc_hd__mux2_1
X_16571_ _04075_ _04280_ _04284_ _04042_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10995_ mapped_spi_flash.cmd_addr\[13\] _07038_ _07039_ VGND VGND VPWR VPWR _07040_
+ sky130_fd_sc_hd__mux2_1
X_18310_ net131 _01838_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15522_ _08581_ _03571_ _03573_ _08535_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__a211o_1
X_12734_ _08061_ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846__593 clknet_1_0__leaf__03680_ VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__inv_2
X_13373__867 clknet_1_1__leaf__08369_ VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__inv_2
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ net1252 _01769_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ CPU.registerFile\[27\]\[28\] CPU.registerFile\[26\]\[28\] _03172_ VGND VGND
+ VPWR VPWR _03507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12665_ _06657_ net2129 _08015_ VGND VGND VPWR VPWR _08025_ sky130_fd_sc_hd__mux2_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14404_ _08646_ _08647_ _08609_ VGND VGND VPWR VPWR _08648_ sky130_fd_sc_hd__mux2_1
X_11616_ _07428_ VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__clkbuf_1
X_18172_ net1183 _01700_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[11\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_108_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15384_ _08580_ _03437_ _03439_ _03218_ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__a211o_1
X_12596_ _07988_ VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17123_ _04821_ _04822_ _06535_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14335_ _08580_ VGND VGND VPWR VPWR _08581_ sky130_fd_sc_hd__buf_4
X_11547_ _07391_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold509 CPU.registerFile\[13\]\[25\] VGND VGND VPWR VPWR net1806 sky130_fd_sc_hd__dlygate4sd3_1
X_17054_ CPU.registerFile\[24\]\[25\] _03724_ _04569_ _04755_ VGND VGND VPWR VPWR
+ _04756_ sky130_fd_sc_hd__o211a_1
X_14266_ CPU.state\[2\] _08252_ VGND VGND VPWR VPWR _08512_ sky130_fd_sc_hd__and2_1
X_11478_ net1709 _07347_ _07333_ VGND VGND VPWR VPWR _07348_ sky130_fd_sc_hd__mux2_1
X_16005_ _06109_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__buf_4
XFILLER_0_111_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13217_ _08330_ VGND VGND VPWR VPWR _08331_ sky130_fd_sc_hd__buf_2
X_10429_ _06675_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__clkbuf_1
X_14197_ clknet_1_0__leaf__08495_ VGND VGND VPWR VPWR _08504_ sky130_fd_sc_hd__buf_1
XFILLER_0_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _08281_ net1529 VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__nor2_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ net1378 VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__clkbuf_1
X_17956_ net967 _01484_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[26\] sky130_fd_sc_hd__dfxtp_1
Xhold1209 CPU.registerFile\[30\]\[5\] VGND VGND VPWR VPWR net2506 sky130_fd_sc_hd__dlygate4sd3_1
X_16907_ _04441_ _04609_ _04611_ _04612_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__a211o_1
X_15591__396 clknet_1_0__leaf__08511_ VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__inv_2
X_17887_ clknet_leaf_21_clk _00038_ VGND VGND VPWR VPWR CPU.cycles\[30\] sky130_fd_sc_hd__dfxtp_1
X_16838_ _06085_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__clkbuf_4
X_15929__668 clknet_1_1__leaf__03688_ VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__inv_2
X_16769_ _04098_ _04463_ _04467_ _04477_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__a31o_2
X_09310_ CPU.PC\[18\] _05636_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__or2_1
X_18508_ net329 _02032_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_09241_ _05567_ _05568_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18439_ net260 _01967_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09172_ _05420_ _05523_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__nor2_1
XFILLER_0_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__08448_ _08448_ VGND VGND VPWR VPWR clknet_0__08448_ sky130_fd_sc_hd__clkbuf_16
X_08956_ CPU.aluIn1\[9\] _05264_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08887_ _05239_ VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__inv_2
X_09508_ net2083 _05853_ _05742_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__mux2_1
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10780_ CPU.aluReg\[31\] CPU.aluReg\[29\] _06872_ VGND VGND VPWR VPWR _06873_ sky130_fd_sc_hd__mux2_1
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09439_ mapped_spi_ram.rcv_data\[4\] _05761_ _05762_ net1401 VGND VGND VPWR VPWR
+ _05788_ sky130_fd_sc_hd__a22o_2
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14145__284 clknet_1_0__leaf__08499_ VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__inv_2
XFILLER_0_81_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12450_ net1809 _07362_ _07906_ VGND VGND VPWR VPWR _07911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11401_ _07298_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12381_ _07874_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_80 clknet_1_0__leaf__08444_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14120_ clknet_1_0__leaf__08495_ VGND VGND VPWR VPWR _08497_ sky130_fd_sc_hd__buf_1
X_11332_ net2386 _06316_ _07260_ VGND VGND VPWR VPWR _07262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11263_ _06641_ net2456 _07223_ VGND VGND VPWR VPWR _07225_ sky130_fd_sc_hd__mux2_1
X_13002_ net2135 _07356_ _08203_ VGND VGND VPWR VPWR _08205_ sky130_fd_sc_hd__mux2_1
X_10214_ _06534_ VGND VGND VPWR VPWR _06535_ sky130_fd_sc_hd__clkbuf_8
X_11194_ mapped_spi_flash.state\[1\] _06979_ VGND VGND VPWR VPWR _07185_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15733__524 clknet_1_0__leaf__03651_ VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__inv_2
X_10145_ _05911_ _06468_ VGND VGND VPWR VPWR _06469_ sky130_fd_sc_hd__nor2_1
X_17810_ net890 _01372_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_18790_ net579 _02314_ VGND VGND VPWR VPWR CPU.aluReg\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17741_ net826 _01307_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_14953_ CPU.registerFile\[8\]\[15\] _03018_ _03019_ _02864_ VGND VGND VPWR VPWR _03020_
+ sky130_fd_sc_hd__o211a_1
X_10076_ _05911_ _06400_ _06402_ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__o21ai_1
X_17672_ net1639 _05203_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__nand2_1
X_14884_ _02943_ _02952_ _02837_ VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__o21a_2
Xclkbuf_1_0__f__08506_ clknet_0__08506_ VGND VGND VPWR VPWR clknet_1_0__leaf__08506_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16623_ _03693_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__08437_ clknet_0__08437_ VGND VGND VPWR VPWR clknet_1_0__leaf__08437_
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_27_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_16
X_14228__359 clknet_1_0__leaf__08507_ VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__inv_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16554_ CPU.registerFile\[6\]\[13\] CPU.registerFile\[7\]\[13\] _04022_ VGND VGND
+ VPWR VPWR _04268_ sky130_fd_sc_hd__mux2_1
X_10978_ _05606_ _05607_ VGND VGND VPWR VPWR _07024_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__08368_ clknet_0__08368_ VGND VGND VPWR VPWR clknet_1_0__leaf__08368_
+ sky130_fd_sc_hd__clkbuf_16
X_15505_ _03556_ _03557_ _08562_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12717_ _06641_ net2655 _08051_ VGND VGND VPWR VPWR _08053_ sky130_fd_sc_hd__mux2_1
X_16485_ _03736_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18224_ net1235 net1317 VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[25\] sky130_fd_sc_hd__dfxtp_1
X_15436_ CPU.registerFile\[0\]\[27\] _08411_ _03490_ _03195_ VGND VGND VPWR VPWR _03491_
+ sky130_fd_sc_hd__o211a_1
X_12648_ _08016_ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18155_ net1166 net1300 VGND VGND VPWR VPWR mapped_spi_ram.rcv_bitcount\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15367_ _03415_ _03423_ _03241_ VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__o21a_2
XFILLER_0_142_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12579_ net2215 _07353_ _07979_ VGND VGND VPWR VPWR _07980_ sky130_fd_sc_hd__mux2_1
X_17106_ CPU.registerFile\[8\]\[27\] _04505_ _04506_ _04805_ VGND VGND VPWR VPWR _04806_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14318_ _08525_ VGND VGND VPWR VPWR _08564_ sky130_fd_sc_hd__clkbuf_8
X_18086_ net1097 _01614_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_15298_ CPU.registerFile\[17\]\[24\] _03036_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__or2_1
Xhold306 per_uart.uart0.enable16_counter\[14\] VGND VGND VPWR VPWR net1603 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold317 CPU.cycles\[22\] VGND VGND VPWR VPWR net1614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 mapped_spi_flash.rbusy VGND VGND VPWR VPWR net1625 sky130_fd_sc_hd__dlygate4sd3_1
X_17037_ CPU.registerFile\[13\]\[25\] _04380_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold339 CPU.rs2\[14\] VGND VGND VPWR VPWR net1636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _05477_ _06127_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__xnor2_2
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ clknet_leaf_18_clk _02508_ VGND VGND VPWR VPWR CPU.aluIn1\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1006 CPU.registerFile\[31\]\[6\] VGND VGND VPWR VPWR net2303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 CPU.registerFile\[23\]\[2\] VGND VGND VPWR VPWR net2314 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ net950 _01467_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[9\] sky130_fd_sc_hd__dfxtp_1
Xhold1028 CPU.registerFile\[31\]\[14\] VGND VGND VPWR VPWR net2325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 CPU.registerFile\[14\]\[14\] VGND VGND VPWR VPWR net2336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15862__608 clknet_1_1__leaf__03681_ VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_18_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09224_ CPU.Iimm\[0\] CPU.Bimm\[11\] CPU.instr\[5\] VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__mux2_2
XFILLER_0_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13960__118 clknet_1_1__leaf__08480_ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__inv_2
XFILLER_0_63_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09155_ _05257_ CPU.aluIn1\[28\] VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13752__1121 clknet_1_1__leaf__08459_ VGND VGND VPWR VPWR net1177 sky130_fd_sc_hd__inv_2
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09086_ CPU.Iimm\[0\] _05248_ _05275_ _05437_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13936__96 clknet_1_1__leaf__08478_ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__inv_2
XFILLER_0_13_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold840 CPU.registerFile\[17\]\[28\] VGND VGND VPWR VPWR net2137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 CPU.registerFile\[26\]\[27\] VGND VGND VPWR VPWR net2148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 CPU.registerFile\[26\]\[20\] VGND VGND VPWR VPWR net2159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 CPU.registerFile\[11\]\[22\] VGND VGND VPWR VPWR net2170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold884 CPU.registerFile\[3\]\[29\] VGND VGND VPWR VPWR net2181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold895 CPU.registerFile\[14\]\[13\] VGND VGND VPWR VPWR net2192 sky130_fd_sc_hd__dlygate4sd3_1
X_09988_ _05451_ _05460_ _06271_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__nand3_1
X_08939_ CPU.aluIn1\[3\] _05268_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11950_ _06611_ net2221 _07598_ VGND VGND VPWR VPWR _07606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10901_ net2671 _06965_ _06868_ VGND VGND VPWR VPWR _06966_ sky130_fd_sc_hd__mux2_1
X_19198__56 VGND VGND VPWR VPWR _19198__56/HI net56 sky130_fd_sc_hd__conb_1
X_11881_ _07569_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__clkbuf_1
X_13620_ clknet_1_0__leaf__08440_ VGND VGND VPWR VPWR _08447_ sky130_fd_sc_hd__buf_1
X_10832_ CPU.aluReg\[19\] CPU.aluReg\[17\] _06906_ VGND VGND VPWR VPWR _06913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10763_ _06855_ VGND VGND VPWR VPWR _06858_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12502_ _07938_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__clkbuf_1
X_16270_ _08404_ _03974_ _03980_ _03990_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__a31o_2
X_13482_ _08432_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__clkbuf_1
X_10694_ _06819_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15221_ _03155_ _03262_ _03281_ _03243_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__a211o_1
X_12433_ net1999 _07345_ _07895_ VGND VGND VPWR VPWR _07902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15152_ _03211_ _03213_ _02851_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__mux2_1
X_15958__694 clknet_1_1__leaf__03691_ VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__inv_2
X_12364_ _07865_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11315_ net1917 _06124_ _07249_ VGND VGND VPWR VPWR _07253_ sky130_fd_sc_hd__mux2_1
X_15083_ CPU.registerFile\[2\]\[18\] CPU.registerFile\[3\]\[18\] _02871_ VGND VGND
+ VPWR VPWR _03147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12295_ net1468 _07813_ VGND VGND VPWR VPWR _07823_ sky130_fd_sc_hd__or2_1
X_15657__455 clknet_1_1__leaf__03644_ VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__inv_2
X_18911_ net685 _02431_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_11246_ _06624_ net2096 _07212_ VGND VGND VPWR VPWR _07216_ sky130_fd_sc_hd__mux2_1
X_18842_ clknet_leaf_8_clk _02366_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11177_ net1592 _07134_ VGND VGND VPWR VPWR _07172_ sky130_fd_sc_hd__or2_1
X_10128_ _05882_ _06452_ VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__or2_1
X_15985_ mapped_spi_ram.rcv_data\[9\] _05858_ _05860_ mapped_spi_flash.rcv_data\[9\]
+ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__a22oi_4
X_18773_ net562 _02297_ VGND VGND VPWR VPWR CPU.aluReg\[3\] sky130_fd_sc_hd__dfxtp_1
X_17724_ net809 _01290_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_14936_ CPU.registerFile\[30\]\[15\] CPU.registerFile\[31\]\[15\] _02887_ VGND VGND
+ VPWR VPWR _03003_ sky130_fd_sc_hd__mux2_1
X_10059_ net2308 _06386_ _06293_ VGND VGND VPWR VPWR _06387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14867_ CPU.registerFile\[13\]\[13\] CPU.registerFile\[12\]\[13\] _02935_ VGND VGND
+ VPWR VPWR _02936_ sky130_fd_sc_hd__mux2_1
X_17655_ _05237_ _05191_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16606_ _03847_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__clkbuf_4
X_17586_ _05146_ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14798_ CPU.registerFile\[5\]\[11\] CPU.registerFile\[4\]\[11\] _08864_ VGND VGND
+ VPWR VPWR _02869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16537_ _03847_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16468_ CPU.registerFile\[10\]\[11\] CPU.registerFile\[11\]\[11\] _03931_ VGND VGND
+ VPWR VPWR _04184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15419_ CPU.registerFile\[24\]\[27\] _08582_ _03473_ _03175_ VGND VGND VPWR VPWR
+ _03474_ sky130_fd_sc_hd__o211a_1
X_18207_ net1218 _01735_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[8\] sky130_fd_sc_hd__dfxtp_1
X_19187_ clknet_leaf_3_clk _02705_ VGND VGND VPWR VPWR per_uart.d_in_uart\[2\] sky130_fd_sc_hd__dfxtp_1
X_16399_ _06140_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_115_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18138_ net1149 _01666_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold103 _08244_ VGND VGND VPWR VPWR net1400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold114 _08218_ VGND VGND VPWR VPWR net1411 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18069_ net1080 _01597_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[11\] sky130_fd_sc_hd__dfxtp_1
Xhold125 _06506_ VGND VGND VPWR VPWR net1422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 mapped_spi_flash.rcv_bitcount\[2\] VGND VGND VPWR VPWR net1433 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_16
Xhold147 mapped_spi_flash.rcv_bitcount\[3\] VGND VGND VPWR VPWR net1444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 _01697_ VGND VGND VPWR VPWR net1455 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _06244_ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__buf_4
Xhold169 mapped_spi_ram.cmd_addr\[13\] VGND VGND VPWR VPWR net1466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09842_ _05556_ _06173_ _06174_ _06175_ _06177_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__o221a_1
Xclkbuf_0__03689_ _03689_ VGND VGND VPWR VPWR clknet_0__03689_ sky130_fd_sc_hd__clkbuf_16
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _05357_ _06094_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__xnor2_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09207_ CPU.aluIn1\[21\] _05545_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09138_ _05362_ CPU.aluIn1\[20\] VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09069_ _05253_ _05415_ _05420_ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__o21ai_1
X_14257__385 clknet_1_1__leaf__08510_ VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__inv_2
X_11100_ _07124_ _07114_ mapped_spi_flash.snd_bitcount\[0\] VGND VGND VPWR VPWR _07125_
+ sky130_fd_sc_hd__mux2_1
X_12080_ _06992_ _07678_ VGND VGND VPWR VPWR _07679_ sky130_fd_sc_hd__and2_1
Xhold670 CPU.registerFile\[15\]\[14\] VGND VGND VPWR VPWR net1967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 CPU.registerFile\[18\]\[5\] VGND VGND VPWR VPWR net1978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 CPU.registerFile\[30\]\[29\] VGND VGND VPWR VPWR net1989 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ _05604_ _07070_ VGND VGND VPWR VPWR _07071_ sky130_fd_sc_hd__nor2_1
X_12982_ _08194_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__clkbuf_1
Xhold1370 CPU.aluReg\[26\] VGND VGND VPWR VPWR net2667 sky130_fd_sc_hd__dlygate4sd3_1
X_14721_ _08574_ _02788_ _02793_ _02746_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__o211a_1
X_13517__909 clknet_1_1__leaf__08436_ VGND VGND VPWR VPWR net965 sky130_fd_sc_hd__inv_2
XFILLER_0_99_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11933_ _07596_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17440_ _08255_ net1707 _06973_ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__o21ai_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _08722_ _02721_ _02725_ _08851_ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__o211a_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11864_ net2093 _07376_ _07525_ VGND VGND VPWR VPWR _07560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03678_ clknet_0__03678_ VGND VGND VPWR VPWR clknet_1_0__leaf__03678_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ CPU.aluReg\[23\] CPU.aluReg\[21\] _06872_ VGND VGND VPWR VPWR _06900_ sky130_fd_sc_hd__mux2_1
X_17371_ _04996_ _04999_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__and2_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ CPU.registerFile\[6\]\[6\] CPU.registerFile\[7\]\[6\] _08740_ VGND VGND VPWR
+ VPWR _08823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11795_ _07523_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__clkbuf_1
X_16322_ _08403_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__clkbuf_4
X_19110_ net93 _02630_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_13943__102 clknet_1_1__leaf__08479_ VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__inv_2
X_10746_ _06846_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19041_ net783 _02561_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_16253_ _08398_ _03971_ _03973_ _08401_ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__a211o_1
X_13465_ _08422_ VGND VGND VPWR VPWR _08423_ sky130_fd_sc_hd__buf_4
XFILLER_0_125_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10677_ _06808_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15204_ _03263_ _03264_ _02937_ VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12416_ net1722 _07328_ _07884_ VGND VGND VPWR VPWR _07893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16184_ CPU.registerFile\[0\]\[4\] _03828_ _03725_ _03906_ VGND VGND VPWR VPWR _03907_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13396_ _05856_ _08376_ _08372_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15739__530 clknet_1_1__leaf__03651_ VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__inv_2
X_15135_ _02826_ _03192_ _03197_ _03151_ VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__o211a_1
X_12347_ _07856_ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15891__634 clknet_1_1__leaf__03684_ VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__inv_2
XFILLER_0_105_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13915__77 clknet_1_0__leaf__08476_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__inv_2
X_15066_ _03006_ _03127_ _03129_ _02814_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__a211o_1
X_12278_ mapped_spi_ram.rcv_data\[11\] _07813_ VGND VGND VPWR VPWR _07814_ sky130_fd_sc_hd__or2_1
X_11229_ _06607_ net1865 _07201_ VGND VGND VPWR VPWR _07207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18825_ net614 _02349_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_18756_ net545 _02280_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[18\] sky130_fd_sc_hd__dfxtp_1
X_15968_ CPU.registerFile\[10\]\[0\] CPU.registerFile\[11\]\[0\] _03694_ VGND VGND
+ VPWR VPWR _03695_ sky130_fd_sc_hd__mux2_1
X_17707_ CPU.mem_wdata\[5\] per_uart.d_in_uart\[5\] _05218_ VGND VGND VPWR VPWR _05229_
+ sky130_fd_sc_hd__mux2_1
X_14919_ _02831_ _02832_ CPU.registerFile\[1\]\[14\] VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18687_ net476 _02211_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_15899_ clknet_1_1__leaf__03654_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__buf_1
X_13751__1120 clknet_1_1__leaf__08459_ VGND VGND VPWR VPWR net1176 sky130_fd_sc_hd__inv_2
X_17638_ per_uart.uart0.rx_ack VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17569_ per_uart.tx_busy per_uart.uart0.tx_wr VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_147_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09825_ _05341_ _05747_ VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__nor2_1
X_09756_ _05351_ _06095_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__xnor2_1
X_17415__37 clknet_1_0__leaf__05014_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__inv_2
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09687_ _05912_ _06029_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__nor2_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17718__49 clknet_1_0__leaf__05015_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__inv_2
X_10600_ net2151 _06413_ _06761_ VGND VGND VPWR VPWR _06767_ sky130_fd_sc_hd__mux2_1
X_11580_ _07408_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__clkbuf_1
X_13254__774 clknet_1_1__leaf__08344_ VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__inv_2
XFILLER_0_153_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10531_ net1941 _06413_ _06724_ VGND VGND VPWR VPWR _06730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15840__588 clknet_1_1__leaf__03679_ VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__inv_2
XFILLER_0_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10462_ _06649_ net2493 _06687_ VGND VGND VPWR VPWR _06693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12201_ _07670_ net1301 net1312 _07762_ _05703_ VGND VGND VPWR VPWR _07763_ sky130_fd_sc_hd__o311a_1
XFILLER_0_150_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13181_ CPU.cycles\[25\] CPU.cycles\[26\] _08299_ VGND VGND VPWR VPWR _08301_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10393_ _06653_ net1975 _06639_ VGND VGND VPWR VPWR _06654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12132_ mapped_spi_ram.cmd_addr\[20\] _07033_ _07704_ VGND VGND VPWR VPWR _07716_
+ sky130_fd_sc_hd__mux2_1
X_14190__325 clknet_1_1__leaf__08503_ VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__inv_2
XFILLER_0_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12063_ CPU.registerFile\[24\]\[3\] _07370_ _07657_ VGND VGND VPWR VPWR _07666_ sky130_fd_sc_hd__mux2_1
X_16940_ _04643_ _04644_ _04279_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__mux2_1
X_11014_ _05619_ _07055_ _05602_ VGND VGND VPWR VPWR _07056_ sky130_fd_sc_hd__o21a_1
X_16871_ CPU.registerFile\[19\]\[20\] CPU.registerFile\[18\]\[20\] _04327_ VGND VGND
+ VPWR VPWR _04578_ sky130_fd_sc_hd__mux2_1
X_18610_ net431 _02134_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_15822_ clknet_1_0__leaf__03654_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__buf_1
XFILLER_0_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15769__556 clknet_1_1__leaf__03655_ VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__inv_2
X_18541_ net362 _02065_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_12965_ _08185_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__clkbuf_1
X_14704_ CPU.registerFile\[13\]\[9\] CPU.registerFile\[12\]\[9\] _08693_ VGND VGND
+ VPWR VPWR _02777_ sky130_fd_sc_hd__mux2_1
X_11916_ _06645_ net1995 _07584_ VGND VGND VPWR VPWR _07588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18472_ net293 _01996_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_14010__162 clknet_1_1__leaf__08486_ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__inv_2
X_14084__230 clknet_1_0__leaf__08492_ VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__inv_2
X_12896_ _05805_ net2027 _08145_ VGND VGND VPWR VPWR _08149_ sky130_fd_sc_hd__mux2_1
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _08425_ _08853_ _08873_ _08597_ VGND VGND VPWR VPWR _08874_ sky130_fd_sc_hd__a211o_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ _07551_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__clkbuf_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _08804_ _08805_ _08609_ VGND VGND VPWR VPWR _08806_ sky130_fd_sc_hd__mux2_1
X_11778_ _06643_ net1879 _07512_ VGND VGND VPWR VPWR _07515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16305_ CPU.registerFile\[5\]\[7\] CPU.registerFile\[4\]\[7\] _04024_ VGND VGND VPWR
+ VPWR _04025_ sky130_fd_sc_hd__mux2_1
X_17285_ clknet_1_0__leaf__03686_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__buf_1
X_10729_ _06837_ VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__clkbuf_1
X_14497_ _08557_ _08734_ _08738_ _08423_ VGND VGND VPWR VPWR _08739_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19024_ net766 _02544_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_16236_ _03736_ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__buf_4
Xclkbuf_1_1__f__08450_ clknet_0__08450_ VGND VGND VPWR VPWR clknet_1_1__leaf__08450_
+ sky130_fd_sc_hd__clkbuf_16
X_13448_ _08408_ VGND VGND VPWR VPWR _08409_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_153_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__08481_ _08481_ VGND VGND VPWR VPWR clknet_0__08481_ sky130_fd_sc_hd__clkbuf_16
X_16167_ _03881_ _03890_ _08406_ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15118_ CPU.registerFile\[13\]\[19\] CPU.registerFile\[12\]\[19\] _02935_ VGND VGND
+ VPWR VPWR _03181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16098_ _03703_ _03820_ _03822_ _03714_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__a211o_1
X_15049_ _03103_ _03113_ _02837_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__o21a_2
XFILLER_0_48_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09610_ CPU.instr\[3\] CPU.instr\[4\] _05738_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__or3b_1
X_18808_ net597 _02332_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_13320__820 clknet_1_1__leaf__08363_ VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__inv_2
X_09541_ CPU.PC\[8\] _05884_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__and2_1
X_18739_ net528 _02263_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09472_ _05393_ _05769_ _05770_ CPU.aluReg\[27\] _05819_ VGND VGND VPWR VPWR _05820_
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_148_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13546__935 clknet_1_0__leaf__08439_ VGND VGND VPWR VPWR net991 sky130_fd_sc_hd__inv_2
XFILLER_0_15_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09808_ net2295 _06145_ _06055_ VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__08470_ clknet_0__08470_ VGND VGND VPWR VPWR clknet_1_0__leaf__08470_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09739_ _06079_ _05999_ VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__xnor2_1
X_12750_ _08070_ VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _07473_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__clkbuf_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _06605_ net2524 _08029_ VGND VGND VPWR VPWR _08034_ sky130_fd_sc_hd__mux2_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ CPU.registerFile\[6\]\[2\] CPU.registerFile\[7\]\[2\] _08522_ VGND VGND VPWR
+ VPWR _08664_ sky130_fd_sc_hd__mux2_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _07436_ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__clkbuf_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14351_ _08596_ VGND VGND VPWR VPWR _08597_ sky130_fd_sc_hd__buf_2
X_11563_ _07399_ VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17070_ CPU.registerFile\[8\]\[26\] _04505_ _04506_ _04770_ VGND VGND VPWR VPWR _04771_
+ sky130_fd_sc_hd__o211a_1
X_10514_ net2098 _06224_ _06713_ VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__mux2_1
X_14282_ _06062_ VGND VGND VPWR VPWR _08528_ sky130_fd_sc_hd__buf_2
X_11494_ net1717 _07358_ _07354_ VGND VGND VPWR VPWR _07359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16021_ _05689_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__buf_4
X_10445_ _06632_ net2336 _06676_ VGND VGND VPWR VPWR _06684_ sky130_fd_sc_hd__mux2_1
X_13629__1010 clknet_1_1__leaf__08447_ VGND VGND VPWR VPWR net1066 sky130_fd_sc_hd__inv_2
X_13164_ net1608 _08289_ VGND VGND VPWR VPWR _08292_ sky130_fd_sc_hd__nor2_1
X_10376_ _06642_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__clkbuf_1
X_12115_ net1312 VGND VGND VPWR VPWR _07703_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17972_ net983 _01500_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_13095_ CPU.state\[1\] VGND VGND VPWR VPWR _08255_ sky130_fd_sc_hd__clkbuf_4
X_16923_ _04503_ _04625_ _04627_ _04509_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__a211o_1
X_12046_ _07634_ VGND VGND VPWR VPWR _07657_ sky130_fd_sc_hd__clkbuf_4
X_16854_ CPU.registerFile\[0\]\[20\] _04233_ _04472_ _04560_ VGND VGND VPWR VPWR _04561_
+ sky130_fd_sc_hd__o211a_1
X_15805_ net1526 _08353_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__nand2_1
X_13997_ clknet_1_0__leaf__08339_ VGND VGND VPWR VPWR _08484_ sky130_fd_sc_hd__buf_1
X_16785_ _06534_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18524_ net345 _02048_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_12948_ _06486_ net2233 _08167_ VGND VGND VPWR VPWR _08176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18455_ net276 _01983_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_12879_ _08139_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__clkbuf_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14618_ _06418_ VGND VGND VPWR VPWR _08857_ sky130_fd_sc_hd__clkbuf_4
X_18386_ net207 _01914_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15823__572 clknet_1_0__leaf__03678_ VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__inv_2
XFILLER_0_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13350__846 clknet_1_1__leaf__08367_ VGND VGND VPWR VPWR net902 sky130_fd_sc_hd__inv_2
XFILLER_0_161_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14549_ _08574_ _08784_ _08789_ _08592_ VGND VGND VPWR VPWR _08790_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15897__640 clknet_1_0__leaf__03684_ VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__inv_2
XFILLER_0_154_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__08502_ clknet_0__08502_ VGND VGND VPWR VPWR clknet_1_1__leaf__08502_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17268_ CPU.registerFile\[27\]\[31\] CPU.registerFile\[26\]\[31\] _04646_ VGND VGND
+ VPWR VPWR _04964_ sky130_fd_sc_hd__mux2_1
X_19007_ clknet_leaf_11_clk _02527_ VGND VGND VPWR VPWR CPU.aluIn1\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15596__401 clknet_1_1__leaf__08511_ VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__inv_2
XFILLER_0_24_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16219_ CPU.registerFile\[5\]\[5\] CPU.registerFile\[4\]\[5\] _03704_ VGND VGND VPWR
+ VPWR _03941_ sky130_fd_sc_hd__mux2_1
X_17199_ _03722_ _04894_ _04896_ _04612_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__a211o_1
XFILLER_0_51_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__08464_ _08464_ VGND VGND VPWR VPWR clknet_0__08464_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__08364_ clknet_0__08364_ VGND VGND VPWR VPWR clknet_1_1__leaf__08364_
+ sky130_fd_sc_hd__clkbuf_16
X_13995__150 clknet_1_1__leaf__08483_ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__inv_2
X_08972_ _05316_ _05323_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__or2_1
Xhold18 _01728_ VGND VGND VPWR VPWR net1315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 mapped_spi_ram.cmd_addr\[27\] VGND VGND VPWR VPWR net1326 sky130_fd_sc_hd__dlygate4sd3_1
X_09524_ _05391_ _05523_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__nor2_1
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09455_ _05789_ _05803_ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__or2_4
XFILLER_0_78_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09386_ CPU.Bimm\[2\] VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10230_ _06549_ _06550_ VGND VGND VPWR VPWR _06551_ sky130_fd_sc_hd__nor2_1
X_13327__826 clknet_1_1__leaf__08364_ VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__inv_2
X_10161_ _06470_ net1439 VGND VGND VPWR VPWR _06485_ sky130_fd_sc_hd__or2_2
X_15952__689 clknet_1_1__leaf__03690_ VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__inv_2
X_10092_ mapped_spi_flash.rcv_data\[13\] _05859_ _06034_ VGND VGND VPWR VPWR _06418_
+ sky130_fd_sc_hd__a21o_4
X_13920_ clknet_1_1__leaf__08473_ VGND VGND VPWR VPWR _08477_ sky130_fd_sc_hd__buf_1
Xclkbuf_1_0__f__08453_ clknet_0__08453_ VGND VGND VPWR VPWR clknet_1_0__leaf__08453_
+ sky130_fd_sc_hd__clkbuf_16
X_12802_ _08097_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__clkbuf_1
X_16570_ _04037_ _04281_ _04283_ _04208_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__a211o_1
X_10994_ _06976_ VGND VGND VPWR VPWR _07039_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _06657_ net2615 _08051_ VGND VGND VPWR VPWR _08061_ sky130_fd_sc_hd__mux2_1
X_15521_ CPU.registerFile\[20\]\[30\] _08523_ _03572_ _08578_ VGND VGND VPWR VPWR
+ _03573_ sky130_fd_sc_hd__o211a_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18240_ net1251 _01768_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_15452_ _03504_ _03505_ _03255_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _08024_ VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__clkbuf_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14403_ CPU.registerFile\[28\]\[2\] CPU.registerFile\[29\]\[2\] _08538_ VGND VGND
+ VPWR VPWR _08647_ sky130_fd_sc_hd__mux2_1
X_11615_ net2000 _07332_ _07427_ VGND VGND VPWR VPWR _07428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18171_ net1182 _01699_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[10\] sky130_fd_sc_hd__dfxtp_1
X_15383_ CPU.registerFile\[24\]\[26\] _08582_ _03438_ _03175_ VGND VGND VPWR VPWR
+ _03439_ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12595_ net2595 _07370_ _07979_ VGND VGND VPWR VPWR _07988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14334_ _06418_ VGND VGND VPWR VPWR _08580_ sky130_fd_sc_hd__buf_4
X_17122_ CPU.registerFile\[28\]\[27\] CPU.registerFile\[29\]\[27\] _04526_ VGND VGND
+ VPWR VPWR _04822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14122__263 clknet_1_1__leaf__08497_ VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__inv_2
X_11546_ net2095 _07332_ _07390_ VGND VGND VPWR VPWR _07391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_918 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14196__331 clknet_1_0__leaf__08503_ VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__inv_2
XFILLER_0_151_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17053_ _04484_ _04485_ CPU.registerFile\[25\]\[25\] VGND VGND VPWR VPWR _04755_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03691_ clknet_0__03691_ VGND VGND VPWR VPWR clknet_1_1__leaf__03691_
+ sky130_fd_sc_hd__clkbuf_16
X_11477_ _06223_ VGND VGND VPWR VPWR _07347_ sky130_fd_sc_hd__clkbuf_4
X_16004_ _03722_ _03723_ _03729_ _03730_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__a211o_1
XFILLER_0_110_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13216_ _08325_ _08327_ _08329_ _05241_ CPU.instr\[2\] VGND VGND VPWR VPWR _08330_
+ sky130_fd_sc_hd__a311oi_4
X_10428_ _06615_ net2250 _06665_ VGND VGND VPWR VPWR _06675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ CPU.cycles\[10\] _08279_ net1528 VGND VGND VPWR VPWR _08282_ sky130_fd_sc_hd__a21oi_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _06630_ net1858 _06618_ VGND VGND VPWR VPWR _06631_ sky130_fd_sc_hd__mux2_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955_ net966 _01483_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_13078_ CPU.registerFile\[4\]\[6\] net1377 _08239_ VGND VGND VPWR VPWR _08245_ sky130_fd_sc_hd__mux2_1
X_12029_ _07648_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__clkbuf_1
X_16906_ _06141_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__clkbuf_4
X_17886_ clknet_leaf_21_clk _00036_ VGND VGND VPWR VPWR CPU.cycles\[29\] sky130_fd_sc_hd__dfxtp_1
X_15710__503 clknet_1_0__leaf__03649_ VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__inv_2
XFILLER_0_79_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16837_ CPU.aluIn1\[19\] _04458_ _04544_ _04259_ VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__o211a_1
X_13575__961 clknet_1_1__leaf__08442_ VGND VGND VPWR VPWR net1017 sky130_fd_sc_hd__inv_2
X_16768_ _04305_ _04470_ _04475_ _04476_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18507_ net328 _02031_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_15719_ clknet_1_1__leaf__03643_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__buf_1
X_13849__1208 clknet_1_1__leaf__08469_ VGND VGND VPWR VPWR net1264 sky130_fd_sc_hd__inv_2
XFILLER_0_119_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16699_ _06141_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__clkbuf_4
X_09240_ _05571_ _05590_ _05591_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__o21a_1
X_18438_ net259 _01966_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09171_ _05522_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__clkbuf_4
X_18369_ net190 _01897_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__08447_ _08447_ VGND VGND VPWR VPWR clknet_0__08447_ sky130_fd_sc_hd__clkbuf_16
X_08955_ _05267_ _05306_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__nor2_2
X_08886_ _05236_ net1480 net1320 _05238_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15650__450 clknet_1_1__leaf__03642_ VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__inv_2
X_09507_ _05852_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__clkbuf_4
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09438_ _05787_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__clkbuf_1
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09369_ net1611 VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11400_ net1785 _06316_ _07296_ VGND VGND VPWR VPWR _07298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12380_ _06645_ net1822 _07870_ VGND VGND VPWR VPWR _07874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_70 _06123_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_81 clknet_1_0__leaf__08341_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11331_ _07261_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11262_ _07224_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13001_ _08204_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__clkbuf_1
X_10213_ _06148_ VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__buf_6
X_11193_ mapped_spi_flash.state\[1\] mapped_spi_flash.state\[0\] _07130_ VGND VGND
+ VPWR VPWR _07184_ sky130_fd_sc_hd__o21ai_1
X_10144_ _05957_ _05959_ VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17740_ net825 _01306_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_14952_ _02733_ _02734_ CPU.registerFile\[9\]\[15\] VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__a21o_1
X_10075_ CPU.cycles\[6\] _05553_ _06197_ _06401_ VGND VGND VPWR VPWR _06402_ sky130_fd_sc_hd__o2bb2a_1
X_17671_ per_uart.uart0.rx_bitcount\[2\] per_uart.uart0.rx_bitcount\[1\] per_uart.uart0.rx_bitcount\[0\]
+ _05194_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__and4_1
X_14883_ _02826_ _02946_ _02951_ _02746_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_0__f__08505_ clknet_0__08505_ VGND VGND VPWR VPWR clknet_1_0__leaf__08505_
+ sky130_fd_sc_hd__clkbuf_16
X_16622_ CPU.aluIn1\[14\] _04054_ _04334_ _04259_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__08436_ clknet_0__08436_ VGND VGND VPWR VPWR clknet_1_0__leaf__08436_
+ sky130_fd_sc_hd__clkbuf_16
X_13297__799 clknet_1_1__leaf__08361_ VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__inv_2
X_16553_ _04015_ _04264_ _04266_ _03979_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__a211o_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10977_ _05558_ VGND VGND VPWR VPWR _07023_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__08367_ clknet_0__08367_ VGND VGND VPWR VPWR clknet_1_0__leaf__08367_
+ sky130_fd_sc_hd__clkbuf_16
X_15504_ CPU.registerFile\[5\]\[29\] CPU.registerFile\[4\]\[29\] _08558_ VGND VGND
+ VPWR VPWR _03557_ sky130_fd_sc_hd__mux2_1
X_12716_ _08052_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__clkbuf_1
X_16484_ _04098_ _04187_ _04191_ _04199_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__a31o_2
XFILLER_0_128_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18223_ net1234 _01751_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15435_ _03235_ _03236_ CPU.registerFile\[1\]\[27\] VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12647_ _06638_ net1950 _08015_ VGND VGND VPWR VPWR _08016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18154_ net1165 _01682_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_bitcount\[0\] sky130_fd_sc_hd__dfxtp_1
X_15366_ _03230_ _03418_ _03422_ _03151_ VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__o211a_1
X_12578_ _07956_ VGND VGND VPWR VPWR _07979_ sky130_fd_sc_hd__buf_4
XFILLER_0_136_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17105_ CPU.registerFile\[9\]\[27\] _04460_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__or2_1
X_11529_ net1708 _07316_ _07379_ VGND VGND VPWR VPWR _07382_ sky130_fd_sc_hd__mux2_1
X_14317_ _08559_ _08561_ _08562_ VGND VGND VPWR VPWR _08563_ sky130_fd_sc_hd__mux2_1
X_18085_ net1096 _01613_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_15297_ CPU.registerFile\[19\]\[24\] CPU.registerFile\[18\]\[24\] _03157_ VGND VGND
+ VPWR VPWR _03355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold307 CPU.cycles\[4\] VGND VGND VPWR VPWR net1604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold318 CPU.cycles\[3\] VGND VGND VPWR VPWR net1615 sky130_fd_sc_hd__dlygate4sd3_1
X_17036_ CPU.registerFile\[15\]\[25\] CPU.registerFile\[14\]\[25\] _04550_ VGND VGND
+ VPWR VPWR _04738_ sky130_fd_sc_hd__mux2_1
Xhold329 _02327_ VGND VGND VPWR VPWR net1626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15935__673 clknet_1_1__leaf__03689_ VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__inv_2
XFILLER_0_21_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ clknet_leaf_17_clk _02507_ VGND VGND VPWR VPWR CPU.aluIn1\[4\] sky130_fd_sc_hd__dfxtp_4
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1007 CPU.registerFile\[13\]\[11\] VGND VGND VPWR VPWR net2304 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1018 CPU.registerFile\[3\]\[23\] VGND VGND VPWR VPWR net2315 sky130_fd_sc_hd__dlygate4sd3_1
X_17938_ net949 _01466_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xhold1029 CPU.registerFile\[11\]\[25\] VGND VGND VPWR VPWR net2326 sky130_fd_sc_hd__dlygate4sd3_1
X_13499__892 clknet_1_0__leaf__08435_ VGND VGND VPWR VPWR net948 sky130_fd_sc_hd__inv_2
X_17869_ clknet_leaf_24_clk _00018_ VGND VGND VPWR VPWR CPU.cycles\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09223_ CPU.aluIn1\[2\] _05574_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_555 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15680__476 clknet_1_0__leaf__03646_ VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__inv_2
X_17322__735 clknet_1_0__leaf__04982_ VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__inv_2
XFILLER_0_16_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09154_ _05396_ _05497_ _05498_ _05505_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__a31o_1
XFILLER_0_115_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09085_ CPU.aluIn1\[0\] VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold830 CPU.registerFile\[23\]\[30\] VGND VGND VPWR VPWR net2127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 CPU.registerFile\[22\]\[16\] VGND VGND VPWR VPWR net2138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold852 CPU.registerFile\[13\]\[15\] VGND VGND VPWR VPWR net2149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold863 CPU.registerFile\[14\]\[27\] VGND VGND VPWR VPWR net2160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 CPU.registerFile\[15\]\[11\] VGND VGND VPWR VPWR net2171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 CPU.registerFile\[28\]\[2\] VGND VGND VPWR VPWR net2182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 CPU.registerFile\[9\]\[12\] VGND VGND VPWR VPWR net2193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09987_ _06317_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__clkbuf_1
X_08938_ _05288_ _05289_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__nor2_2
X_10900_ CPU.aluIn1\[2\] _06964_ _06880_ VGND VGND VPWR VPWR _06965_ sky130_fd_sc_hd__mux2_1
X_11880_ _06609_ net1969 _07562_ VGND VGND VPWR VPWR _07569_ sky130_fd_sc_hd__mux2_1
X_10831_ _06912_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10762_ net9 VGND VGND VPWR VPWR _06857_ sky130_fd_sc_hd__inv_2
X_12501_ net2069 _07345_ _07931_ VGND VGND VPWR VPWR _07938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13481_ CPU.Bimm\[10\] _05763_ _08416_ VGND VGND VPWR VPWR _08432_ sky130_fd_sc_hd__mux2_1
X_10693_ net1997 _05786_ _06816_ VGND VGND VPWR VPWR _06819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15220_ _03271_ _03280_ _03241_ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__o21a_2
X_12432_ _07901_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17297__712 clknet_1_0__leaf__04980_ VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__inv_2
XFILLER_0_63_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15151_ CPU.registerFile\[28\]\[20\] CPU.registerFile\[29\]\[20\] _03212_ VGND VGND
+ VPWR VPWR _03213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12363_ _06628_ net1902 _07859_ VGND VGND VPWR VPWR _07865_ sky130_fd_sc_hd__mux2_1
X_11314_ _07252_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__clkbuf_1
X_15082_ _03144_ _03145_ _03025_ VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__mux2_1
X_12294_ net1468 _07812_ _07821_ _07822_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18910_ net684 _02430_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_11245_ _07215_ VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__clkbuf_1
X_13848__1207 clknet_1_1__leaf__08469_ VGND VGND VPWR VPWR net1263 sky130_fd_sc_hd__inv_2
XFILLER_0_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18841_ clknet_leaf_7_clk net1509 VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_14234__364 clknet_1_1__leaf__08508_ VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__inv_2
X_11176_ net1592 _07160_ _07171_ _07164_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__o211a_1
X_10127_ CPU.PC\[3\] CPU.PC\[2\] CPU.PC\[4\] VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__a21oi_1
X_18772_ net561 _02296_ VGND VGND VPWR VPWR CPU.aluReg\[2\] sky130_fd_sc_hd__dfxtp_1
X_15984_ CPU.registerFile\[12\]\[0\] _03707_ _03708_ _03710_ VGND VGND VPWR VPWR _03711_
+ sky130_fd_sc_hd__o211a_1
X_17723_ net808 _01289_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_10058_ _06385_ VGND VGND VPWR VPWR _06386_ sky130_fd_sc_hd__buf_4
X_14935_ _08837_ _02999_ _03001_ _08802_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17654_ _04986_ _05185_ _05189_ _05190_ VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_159_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14866_ _06061_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__buf_4
X_16605_ CPU.registerFile\[27\]\[14\] CPU.registerFile\[26\]\[14\] _04242_ VGND VGND
+ VPWR VPWR _04318_ sky130_fd_sc_hd__mux2_1
X_17585_ per_uart.uart0.tx_bitcount\[0\] _05145_ _06854_ VGND VGND VPWR VPWR _05146_
+ sky130_fd_sc_hd__mux2_1
X_14797_ CPU.registerFile\[6\]\[11\] CPU.registerFile\[7\]\[11\] _08740_ VGND VGND
+ VPWR VPWR _02868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16536_ CPU.registerFile\[19\]\[12\] CPU.registerFile\[18\]\[12\] _03923_ VGND VGND
+ VPWR VPWR _04251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13689__1063 clknet_1_0__leaf__08454_ VGND VGND VPWR VPWR net1119 sky130_fd_sc_hd__inv_2
XFILLER_0_73_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16467_ CPU.aluIn1\[10\] _04054_ _04183_ _03855_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18206_ net1217 net1342 VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[7\] sky130_fd_sc_hd__dfxtp_1
X_15418_ _08566_ _08568_ CPU.registerFile\[25\]\[27\] VGND VGND VPWR VPWR _03473_
+ sky130_fd_sc_hd__a21o_1
X_19186_ clknet_leaf_3_clk _02704_ VGND VGND VPWR VPWR per_uart.d_in_uart\[1\] sky130_fd_sc_hd__dfxtp_1
X_16398_ CPU.registerFile\[0\]\[9\] _03828_ _04068_ _04115_ VGND VGND VPWR VPWR _04116_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18137_ net1148 _01665_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_15349_ _06013_ _03401_ _03405_ _03092_ VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold104 mapped_spi_flash.rcv_data\[4\] VGND VGND VPWR VPWR net1401 sky130_fd_sc_hd__buf_1
Xhold115 mapped_spi_ram.cmd_addr\[18\] VGND VGND VPWR VPWR net1412 sky130_fd_sc_hd__dlygate4sd3_1
X_18068_ net1079 _01596_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold126 _08249_ VGND VGND VPWR VPWR net1423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold137 _07194_ VGND VGND VPWR VPWR net1434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold148 _02220_ VGND VGND VPWR VPWR net1445 sky130_fd_sc_hd__dlygate4sd3_1
X_17019_ _04441_ _04719_ _04721_ _04612_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__a211o_1
X_09910_ _05745_ _06234_ _06239_ _06243_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__a211o_2
Xhold159 mapped_spi_flash.snd_bitcount\[3\] VGND VGND VPWR VPWR net1456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09841_ _05520_ _05728_ _06176_ VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__a21boi_4
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__03688_ _03688_ VGND VGND VPWR VPWR clknet_0__03688_ sky130_fd_sc_hd__clkbuf_16
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ CPU.PC\[18\] _05891_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__xnor2_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18234__18 VGND VGND VPWR VPWR _18234__18/HI net18 sky130_fd_sc_hd__conb_1
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15762__551 clknet_1_1__leaf__03653_ VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__inv_2
XFILLER_0_147_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09206_ _05557_ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09137_ _05374_ _05379_ _05488_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__and3_1
XFILLER_0_161_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09068_ _05418_ _05419_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__nor2_2
XFILLER_0_4_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold660 CPU.registerFile\[15\]\[12\] VGND VGND VPWR VPWR net1957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 CPU.registerFile\[27\]\[17\] VGND VGND VPWR VPWR net1968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 CPU.registerFile\[2\]\[22\] VGND VGND VPWR VPWR net1979 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ CPU.aluIn1\[8\] CPU.Bimm\[8\] _07055_ VGND VGND VPWR VPWR _07070_ sky130_fd_sc_hd__a21oi_1
Xhold693 CPU.registerFile\[13\]\[0\] VGND VGND VPWR VPWR net1990 sky130_fd_sc_hd__dlygate4sd3_1
X_12981_ net2043 _07335_ _08192_ VGND VGND VPWR VPWR _08194_ sky130_fd_sc_hd__mux2_1
Xhold1360 CPU.Jimm\[19\] VGND VGND VPWR VPWR net2657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1371 CPU.aluReg\[17\] VGND VGND VPWR VPWR net2668 sky130_fd_sc_hd__dlygate4sd3_1
X_14720_ _08785_ _02789_ _02792_ _08870_ VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__a211o_1
X_11932_ _06661_ net1731 _07561_ VGND VGND VPWR VPWR _07596_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ _07559_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__clkbuf_1
X_14651_ _08764_ _02722_ _02724_ _08552_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__a211o_1
XFILLER_0_86_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _06899_ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__clkbuf_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ per_uart.uart0.rxd_reg\[4\] _04992_ _04993_ per_uart.uart0.rxd_reg\[3\] VGND
+ VGND VPWR VPWR _04999_ sky130_fd_sc_hd__a22o_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14582_ _08557_ _08817_ _08821_ _08423_ VGND VGND VPWR VPWR _08822_ sky130_fd_sc_hd__o211a_1
X_11794_ _06659_ net2189 _07489_ VGND VGND VPWR VPWR _07523_ sky130_fd_sc_hd__mux2_1
X_16321_ _04037_ _04038_ _04040_ _03803_ VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__a211o_1
X_10745_ net2437 _06465_ _06838_ VGND VGND VPWR VPWR _06846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19040_ net782 _02560_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_16252_ CPU.registerFile\[8\]\[6\] _08394_ _06150_ _03972_ VGND VGND VPWR VPWR _03973_
+ sky130_fd_sc_hd__o211a_1
X_13464_ _06363_ VGND VGND VPWR VPWR _08422_ sky130_fd_sc_hd__buf_6
X_10676_ net2640 _06486_ _06799_ VGND VGND VPWR VPWR _06808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15203_ CPU.registerFile\[13\]\[21\] CPU.registerFile\[12\]\[21\] _02935_ VGND VGND
+ VPWR VPWR _03264_ sky130_fd_sc_hd__mux2_1
X_12415_ _07892_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__clkbuf_1
X_13231__753 clknet_1_1__leaf__08342_ VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__inv_2
XFILLER_0_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16183_ _03726_ _03727_ CPU.registerFile\[1\]\[4\] VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__a21o_1
X_13395_ _05530_ _05696_ _06203_ VGND VGND VPWR VPWR _08376_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12346_ _06611_ net2005 _07848_ VGND VGND VPWR VPWR _07856_ sky130_fd_sc_hd__mux2_1
X_15134_ _03027_ _03193_ _03196_ _03111_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__a211o_1
XFILLER_0_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15065_ CPU.registerFile\[24\]\[18\] _02928_ _03128_ _02771_ VGND VGND VPWR VPWR
+ _03129_ sky130_fd_sc_hd__o211a_1
X_12277_ _07786_ VGND VGND VPWR VPWR _07813_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11228_ _07206_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18824_ net613 _02348_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_11159_ net2613 _07149_ VGND VGND VPWR VPWR _07162_ sky130_fd_sc_hd__or2_1
X_18755_ net544 _02279_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[17\] sky130_fd_sc_hd__dfxtp_1
X_15967_ _03693_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__buf_4
X_17706_ _05228_ VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__clkbuf_1
X_14918_ CPU.registerFile\[2\]\[14\] CPU.registerFile\[3\]\[14\] _02871_ VGND VGND
+ VPWR VPWR _02986_ sky130_fd_sc_hd__mux2_1
X_18686_ net475 _02210_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17637_ net2632 VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__clkbuf_1
X_14849_ CPU.registerFile\[16\]\[13\] _02755_ _02917_ _02757_ VGND VGND VPWR VPWR
+ _02918_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17568_ _08360_ _05118_ _05131_ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16519_ _03985_ _03986_ CPU.registerFile\[1\]\[12\] VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17499_ _05055_ _06221_ _05061_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19169_ clknet_leaf_0_clk _02689_ VGND VGND VPWR VPWR per_uart.rx_avail sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09824_ _05424_ _06157_ _06160_ _05516_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__o211a_1
X_09755_ _05356_ _06094_ _05482_ VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__a21oi_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09686_ _06028_ _06004_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__xnor2_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17346__7 clknet_1_0__leaf__04984_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__inv_2
XFILLER_0_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17328__741 clknet_1_1__leaf__04982_ VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__inv_2
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13847__1206 clknet_1_0__leaf__08469_ VGND VGND VPWR VPWR net1262 sky130_fd_sc_hd__inv_2
XFILLER_0_107_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10530_ _06729_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10461_ _06692_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12200_ _07703_ _07761_ VGND VGND VPWR VPWR _07762_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13180_ net1645 _08299_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__xor2_1
X_10392_ _06464_ VGND VGND VPWR VPWR _06653_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12131_ _07695_ VGND VGND VPWR VPWR _07715_ sky130_fd_sc_hd__clkbuf_2
X_13523__914 clknet_1_1__leaf__08437_ VGND VGND VPWR VPWR net970 sky130_fd_sc_hd__inv_2
X_12062_ _07665_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__clkbuf_1
Xhold490 CPU.registerFile\[28\]\[3\] VGND VGND VPWR VPWR net1787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11013_ _07025_ _05601_ VGND VGND VPWR VPWR _07055_ sky130_fd_sc_hd__nor2_1
X_13688__1062 clknet_1_0__leaf__08454_ VGND VGND VPWR VPWR net1118 sky130_fd_sc_hd__inv_2
X_16870_ _04575_ _04576_ _04365_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18540_ net361 _02064_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_15752_ clknet_1_1__leaf__03643_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__buf_1
X_12964_ net1891 _07318_ _08181_ VGND VGND VPWR VPWR _08185_ sky130_fd_sc_hd__mux2_1
Xhold1190 CPU.registerFile\[31\]\[18\] VGND VGND VPWR VPWR net2487 sky130_fd_sc_hd__dlygate4sd3_1
X_14703_ CPU.registerFile\[15\]\[9\] CPU.registerFile\[14\]\[9\] _08771_ VGND VGND
+ VPWR VPWR _02776_ sky130_fd_sc_hd__mux2_1
X_18471_ net292 _01995_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_11915_ _07587_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__clkbuf_1
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _08148_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__clkbuf_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ _08862_ _08872_ _08594_ VGND VGND VPWR VPWR _08873_ sky130_fd_sc_hd__o21a_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ net2578 _07358_ _07548_ VGND VGND VPWR VPWR _07551_ sky130_fd_sc_hd__mux2_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14565_ CPU.registerFile\[28\]\[6\] CPU.registerFile\[29\]\[6\] _08538_ VGND VGND
+ VPWR VPWR _08805_ sky130_fd_sc_hd__mux2_1
X_11777_ _07514_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _03744_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__buf_4
XFILLER_0_71_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10728_ net2066 _06267_ _06827_ VGND VGND VPWR VPWR _06837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14496_ _08520_ _08735_ _08737_ _08661_ VGND VGND VPWR VPWR _08738_ sky130_fd_sc_hd__a211o_1
XFILLER_0_83_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19023_ net765 _02543_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16235_ _03735_ _03952_ _03956_ _03755_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__o211a_1
X_13447_ _06058_ _06059_ VGND VGND VPWR VPWR _08408_ sky130_fd_sc_hd__nand2_1
X_10659_ _06776_ VGND VGND VPWR VPWR _06799_ sky130_fd_sc_hd__buf_4
XFILLER_0_23_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__08480_ _08480_ VGND VGND VPWR VPWR clknet_0__08480_ sky130_fd_sc_hd__clkbuf_16
X_13378_ clknet_1_0__leaf__08366_ VGND VGND VPWR VPWR _08370_ sky130_fd_sc_hd__buf_1
X_16166_ _03758_ _03885_ _03889_ _03775_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15117_ CPU.registerFile\[15\]\[19\] CPU.registerFile\[14\]\[19\] _03013_ VGND VGND
+ VPWR VPWR _03180_ sky130_fd_sc_hd__mux2_1
X_12329_ _07846_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__clkbuf_1
X_16097_ CPU.registerFile\[12\]\[2\] _03707_ _03708_ _03821_ VGND VGND VPWR VPWR _03822_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15048_ _02826_ _03107_ _03112_ _02746_ VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__o211a_1
X_13769__1136 clknet_1_1__leaf__08461_ VGND VGND VPWR VPWR net1192 sky130_fd_sc_hd__inv_2
X_18807_ net596 _02331_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_16999_ _04503_ _04699_ _04701_ _04509_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__a211o_1
X_09540_ CPU.PC\[7\] CPU.PC\[6\] _05883_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__and3_1
X_18738_ net527 _02262_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[0\] sky130_fd_sc_hd__dfxtp_1
X_09471_ _05394_ _05807_ _05817_ _05818_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__a2bb2o_1
X_18669_ net458 _02193_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09807_ _06144_ VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__buf_4
X_09738_ _05925_ _05995_ _06000_ VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__a21bo_1
X_14068__215 clknet_1_0__leaf__08491_ VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__inv_2
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ mapped_spi_ram.rcv_data\[14\] _05858_ _05860_ net1600 VGND VGND VPWR VPWR
+ _06012_ sky130_fd_sc_hd__a22oi_4
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ net2508 _07349_ _07464_ VGND VGND VPWR VPWR _07473_ sky130_fd_sc_hd__mux2_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _08033_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__clkbuf_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11631_ net1991 _07349_ _07427_ VGND VGND VPWR VPWR _07436_ sky130_fd_sc_hd__mux2_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11562_ net2085 _07349_ _07390_ VGND VGND VPWR VPWR _07399_ sky130_fd_sc_hd__mux2_1
X_14350_ _08264_ VGND VGND VPWR VPWR _08596_ sky130_fd_sc_hd__buf_4
XFILLER_0_64_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10513_ _06720_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__clkbuf_1
X_14281_ _08526_ VGND VGND VPWR VPWR _08527_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_162_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11493_ net1332 VGND VGND VPWR VPWR _07358_ sky130_fd_sc_hd__buf_4
X_16020_ _06534_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__buf_2
XFILLER_0_107_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10444_ _06683_ VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13163_ CPU.cycles\[18\] _08289_ VGND VGND VPWR VPWR _08291_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10375_ _06641_ net1896 _06639_ VGND VGND VPWR VPWR _06642_ sky130_fd_sc_hd__mux2_1
X_12114_ net1325 _07693_ _07702_ _07175_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__o211a_1
X_17971_ net982 _01499_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_13094_ _05538_ _06175_ _05729_ VGND VGND VPWR VPWR _08254_ sky130_fd_sc_hd__a21oi_2
X_16922_ CPU.registerFile\[8\]\[22\] _04505_ _04506_ _04626_ VGND VGND VPWR VPWR _04627_
+ sky130_fd_sc_hd__o211a_1
X_12045_ _07656_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__clkbuf_1
X_13304__805 clknet_1_0__leaf__08362_ VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__inv_2
X_16853_ _04389_ _04390_ CPU.registerFile\[1\]\[20\] VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__a21o_1
X_15804_ _08353_ _03670_ _03661_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__a21oi_1
X_16784_ CPU.registerFile\[19\]\[18\] CPU.registerFile\[18\]\[18\] _04327_ VGND VGND
+ VPWR VPWR _04493_ sky130_fd_sc_hd__mux2_1
X_18523_ net344 _02047_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12947_ _08175_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13493__887 clknet_1_0__leaf__08434_ VGND VGND VPWR VPWR net943 sky130_fd_sc_hd__inv_2
X_18454_ net275 _01982_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _06465_ net2462 _08131_ VGND VGND VPWR VPWR _08139_ sky130_fd_sc_hd__mux2_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ _08854_ _08855_ _08695_ VGND VGND VPWR VPWR _08856_ sky130_fd_sc_hd__mux2_1
X_11829_ net2581 _07341_ _07537_ VGND VGND VPWR VPWR _07542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18385_ net206 _01913_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15597_ clknet_1_1__leaf__08506_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__buf_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14548_ _08785_ _08786_ _08788_ _08590_ VGND VGND VPWR VPWR _08789_ sky130_fd_sc_hd__a211o_1
XFILLER_0_44_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__08501_ clknet_0__08501_ VGND VGND VPWR VPWR clknet_1_1__leaf__08501_
+ sky130_fd_sc_hd__clkbuf_16
X_17267_ _04961_ _04962_ _06535_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__mux2_1
X_14479_ _08521_ _08717_ _08720_ _08533_ VGND VGND VPWR VPWR _08721_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19006_ clknet_leaf_12_clk _02526_ VGND VGND VPWR VPWR CPU.aluIn1\[23\] sky130_fd_sc_hd__dfxtp_2
X_16218_ CPU.registerFile\[6\]\[5\] CPU.registerFile\[7\]\[5\] _03717_ VGND VGND VPWR
+ VPWR _03940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17198_ CPU.registerFile\[24\]\[29\] _03724_ _04569_ _04895_ VGND VGND VPWR VPWR
+ _04896_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__08463_ _08463_ VGND VGND VPWR VPWR clknet_0__08463_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__08363_ clknet_0__08363_ VGND VGND VPWR VPWR clknet_1_1__leaf__08363_
+ sky130_fd_sc_hd__clkbuf_16
X_16149_ CPU.registerFile\[30\]\[3\] CPU.registerFile\[31\]\[3\] _03796_ VGND VGND
+ VPWR VPWR _03873_ sky130_fd_sc_hd__mux2_1
X_14173__310 clknet_1_1__leaf__08501_ VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__inv_2
XFILLER_0_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08971_ CPU.aluIn1\[13\] _05322_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__and2_1
X_13846__1205 clknet_1_0__leaf__08469_ VGND VGND VPWR VPWR net1261 sky130_fd_sc_hd__inv_2
Xhold19 mapped_spi_ram.cmd_addr\[25\] VGND VGND VPWR VPWR net1316 sky130_fd_sc_hd__dlygate4sd3_1
X_14017__169 clknet_1_0__leaf__08486_ VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__inv_2
X_18579__36 VGND VGND VPWR VPWR _18579__36/HI net36 sky130_fd_sc_hd__conb_1
XFILLER_0_97_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09523_ _05388_ _05532_ _05535_ CPU.aluReg\[24\] _05867_ VGND VGND VPWR VPWR _05868_
+ sky130_fd_sc_hd__a221o_1
X_09454_ CPU.Bimm\[8\] _05550_ _05790_ CPU.cycles\[28\] _05802_ VGND VGND VPWR VPWR
+ _05803_ sky130_fd_sc_hd__a221o_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15906__648 clknet_1_1__leaf__03685_ VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__inv_2
XFILLER_0_149_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09385_ CPU.Bimm\[3\] VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15605__409 clknet_1_1__leaf__03638_ VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__inv_2
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_862 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17291__707 clknet_1_1__leaf__04979_ VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__inv_2
XFILLER_0_30_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10160_ _06176_ _06476_ _06483_ _05541_ VGND VGND VPWR VPWR _06484_ sky130_fd_sc_hd__a22o_1
X_10091_ _05691_ _06240_ VGND VGND VPWR VPWR _06417_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__08452_ clknet_0__08452_ VGND VGND VPWR VPWR clknet_1_0__leaf__08452_
+ sky130_fd_sc_hd__clkbuf_16
X_12801_ _06657_ net2571 _08087_ VGND VGND VPWR VPWR _08097_ sky130_fd_sc_hd__mux2_1
X_10993_ _07023_ _07036_ _07037_ _06853_ VGND VGND VPWR VPWR _07038_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15520_ CPU.registerFile\[21\]\[30\] _02752_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__or2_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _08060_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18593__50 VGND VGND VPWR VPWR _18593__50/HI net50 sky130_fd_sc_hd__conb_1
X_15451_ CPU.registerFile\[28\]\[28\] CPU.registerFile\[29\]\[28\] _03212_ VGND VGND
+ VPWR VPWR _03505_ sky130_fd_sc_hd__mux2_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _06655_ net2121 _08015_ VGND VGND VPWR VPWR _08024_ sky130_fd_sc_hd__mux2_1
X_13768__1135 clknet_1_1__leaf__08461_ VGND VGND VPWR VPWR net1191 sky130_fd_sc_hd__inv_2
XFILLER_0_139_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ CPU.registerFile\[30\]\[2\] CPU.registerFile\[31\]\[2\] _08645_ VGND VGND
+ VPWR VPWR _08646_ sky130_fd_sc_hd__mux2_1
X_11614_ _07415_ VGND VGND VPWR VPWR _07427_ sky130_fd_sc_hd__buf_4
X_18170_ net1181 _01698_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[9\] sky130_fd_sc_hd__dfxtp_2
X_15382_ _08566_ _08568_ CPU.registerFile\[25\]\[26\] VGND VGND VPWR VPWR _03438_
+ sky130_fd_sc_hd__a21o_1
X_12594_ _07987_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17121_ CPU.registerFile\[30\]\[27\] CPU.registerFile\[31\]\[27\] _04605_ VGND VGND
+ VPWR VPWR _04821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14333_ _08575_ _08577_ _08578_ VGND VGND VPWR VPWR _08579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11545_ _07378_ VGND VGND VPWR VPWR _07390_ sky130_fd_sc_hd__buf_4
XFILLER_0_107_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13529__920 clknet_1_0__leaf__08437_ VGND VGND VPWR VPWR net976 sky130_fd_sc_hd__inv_2
XFILLER_0_108_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17052_ CPU.registerFile\[27\]\[25\] CPU.registerFile\[26\]\[25\] _04646_ VGND VGND
+ VPWR VPWR _04754_ sky130_fd_sc_hd__mux2_1
X_11476_ _07346_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14264_ clknet_1_0__leaf__08506_ VGND VGND VPWR VPWR _08511_ sky130_fd_sc_hd__buf_1
Xclkbuf_1_1__f__03690_ clknet_0__03690_ VGND VGND VPWR VPWR clknet_1_1__leaf__03690_
+ sky130_fd_sc_hd__clkbuf_16
X_13979__135 clknet_1_0__leaf__08482_ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__inv_2
X_16003_ _06140_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__buf_4
X_10427_ _06674_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__clkbuf_1
X_13215_ _05527_ _08328_ VGND VGND VPWR VPWR _08329_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10358_ _06199_ VGND VGND VPWR VPWR _06630_ sky130_fd_sc_hd__buf_4
X_13146_ CPU.cycles\[10\] CPU.cycles\[11\] _08279_ VGND VGND VPWR VPWR _08281_ sky130_fd_sc_hd__and3_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ net1400 VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__clkbuf_1
X_17954_ net965 _01482_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_10289_ net1939 _06386_ _06580_ VGND VGND VPWR VPWR _06585_ sky130_fd_sc_hd__mux2_1
X_12028_ CPU.registerFile\[24\]\[20\] _07335_ _07646_ VGND VGND VPWR VPWR _07648_
+ sky130_fd_sc_hd__mux2_1
X_16905_ CPU.registerFile\[24\]\[21\] _04319_ _04569_ _04610_ VGND VGND VPWR VPWR
+ _04611_ sky130_fd_sc_hd__o211a_1
X_17885_ clknet_leaf_23_clk _00035_ VGND VGND VPWR VPWR CPU.cycles\[28\] sky130_fd_sc_hd__dfxtp_1
X_16836_ _04141_ _04524_ _04543_ _04500_ VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__a211o_1
X_13501__894 clknet_1_0__leaf__08435_ VGND VGND VPWR VPWR net950 sky130_fd_sc_hd__inv_2
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16767_ _06108_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__buf_4
X_18506_ net327 _02030_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16698_ CPU.registerFile\[16\]\[16\] _04252_ _04090_ _04408_ VGND VGND VPWR VPWR
+ _04409_ sky130_fd_sc_hd__o211a_1
X_18437_ net258 _01965_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14205__339 clknet_1_1__leaf__08504_ VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__inv_2
XFILLER_0_91_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09170_ _05521_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__clkbuf_4
X_18368_ net189 _01896_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18299_ net120 _01827_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__08446_ _08446_ VGND VGND VPWR VPWR clknet_0__08446_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08954_ _05292_ _05301_ _05305_ _05295_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__o2bb2a_1
X_15912__652 clknet_1_1__leaf__03687_ VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__inv_2
X_08885_ _05237_ _05238_ net1480 net1320 VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_98_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13828__1189 clknet_1_0__leaf__08467_ VGND VGND VPWR VPWR net1245 sky130_fd_sc_hd__inv_2
X_09506_ CPU.Bimm\[5\] _05758_ _05759_ CPU.cycles\[25\] net1641 VGND VGND VPWR VPWR
+ _05852_ sky130_fd_sc_hd__a221o_4
XFILLER_0_66_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09437_ net2178 _05786_ _05742_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__mux2_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09368_ per_uart.rx_error _05717_ _05719_ per_uart.rx_data\[7\] VGND VGND VPWR VPWR
+ _05720_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_93_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09299_ CPU.PC\[22\] _05643_ _05650_ _05235_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__o211a_1
XANTENNA_60 clknet_1_1__leaf__08448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_71 _06142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 _06053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11330_ net2374 _06292_ _07260_ VGND VGND VPWR VPWR _07261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11261_ _06638_ net2231 _07223_ VGND VGND VPWR VPWR _07224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13000_ net2366 _07353_ _08203_ VGND VGND VPWR VPWR _08204_ sky130_fd_sc_hd__mux2_1
X_10212_ mapped_spi_ram.rcv_data\[24\] _05858_ _05860_ net1356 _06462_ VGND VGND VPWR
+ VPWR _06533_ sky130_fd_sc_hd__a221o_1
X_11192_ net1393 mapped_spi_flash.state\[3\] VGND VGND VPWR VPWR _07183_ sky130_fd_sc_hd__nand2_1
X_10143_ CPU.PC\[3\] CPU.PC\[2\] VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__xor2_1
XFILLER_0_101_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14951_ _08410_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__clkbuf_4
X_10074_ CPU.PC\[6\] _05883_ VGND VGND VPWR VPWR _06401_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13559__946 clknet_1_1__leaf__08441_ VGND VGND VPWR VPWR net1002 sky130_fd_sc_hd__inv_2
X_17670_ _05201_ _05199_ _05202_ _05194_ _05237_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__a221oi_1
X_14882_ _08785_ _02947_ _02950_ _08870_ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_0__f__08504_ clknet_0__08504_ VGND VGND VPWR VPWR clknet_1_0__leaf__08504_
+ sky130_fd_sc_hd__clkbuf_16
X_16621_ _04141_ _04314_ _04333_ _04096_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_0__f__08435_ clknet_0__08435_ VGND VGND VPWR VPWR clknet_1_0__leaf__08435_
+ sky130_fd_sc_hd__clkbuf_16
X_16552_ CPU.registerFile\[12\]\[13\] _04017_ _04018_ _04265_ VGND VGND VPWR VPWR
+ _04266_ sky130_fd_sc_hd__o211a_1
X_13764_ clknet_1_0__leaf__08451_ VGND VGND VPWR VPWR _08461_ sky130_fd_sc_hd__buf_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10976_ net1525 _07007_ _07022_ _07014_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_0__f__08366_ clknet_0__08366_ VGND VGND VPWR VPWR clknet_1_0__leaf__08366_
+ sky130_fd_sc_hd__clkbuf_16
X_15503_ CPU.registerFile\[6\]\[29\] CPU.registerFile\[7\]\[29\] _08536_ VGND VGND
+ VPWR VPWR _03556_ sky130_fd_sc_hd__mux2_1
X_12715_ _06638_ net2546 _08051_ VGND VGND VPWR VPWR _08052_ sky130_fd_sc_hd__mux2_1
X_16483_ _03901_ _04194_ _04198_ _04072_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__o211a_1
X_18222_ net1233 _01750_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[23\] sky130_fd_sc_hd__dfxtp_1
X_15434_ CPU.registerFile\[2\]\[27\] CPU.registerFile\[3\]\[27\] _03275_ VGND VGND
+ VPWR VPWR _03489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13845__1204 clknet_1_0__leaf__08469_ VGND VGND VPWR VPWR net1260 sky130_fd_sc_hd__inv_2
X_12646_ _07992_ VGND VGND VPWR VPWR _08015_ sky130_fd_sc_hd__buf_4
XFILLER_0_109_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14046__195 clknet_1_1__leaf__08489_ VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__inv_2
XFILLER_0_109_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18153_ net1164 _01681_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15365_ _08414_ _03419_ _03421_ _03111_ VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__a211o_1
X_12577_ _07978_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17104_ CPU.registerFile\[10\]\[27\] CPU.registerFile\[11\]\[27\] _06173_ VGND VGND
+ VPWR VPWR _04804_ sky130_fd_sc_hd__mux2_1
X_14316_ _08540_ VGND VGND VPWR VPWR _08562_ sky130_fd_sc_hd__buf_4
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11528_ _07381_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18084_ net1095 _01612_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15296_ net1574 _03201_ _03354_ _02993_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold308 mapped_spi_flash.rcv_data\[8\] VGND VGND VPWR VPWR net1605 sky130_fd_sc_hd__dlygate4sd3_1
X_17035_ _04503_ _04734_ _04736_ _04509_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__a211o_1
Xhold319 CPU.cycles\[28\] VGND VGND VPWR VPWR net1616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11459_ _06082_ VGND VGND VPWR VPWR _07335_ sky130_fd_sc_hd__buf_4
XFILLER_0_123_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ net1615 _08269_ VGND VGND VPWR VPWR _08272_ sky130_fd_sc_hd__nor2_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ clknet_leaf_17_clk _02506_ VGND VGND VPWR VPWR CPU.aluIn1\[3\] sky130_fd_sc_hd__dfxtp_2
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15634__435 clknet_1_0__leaf__03641_ VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__inv_2
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1008 CPU.registerFile\[12\]\[8\] VGND VGND VPWR VPWR net2305 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17937_ net948 _01465_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold1019 CPU.registerFile\[22\]\[17\] VGND VGND VPWR VPWR net2316 sky130_fd_sc_hd__dlygate4sd3_1
X_17868_ clknet_leaf_24_clk _00017_ VGND VGND VPWR VPWR CPU.cycles\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16819_ CPU.registerFile\[28\]\[19\] CPU.registerFile\[29\]\[19\] _04526_ VGND VGND
+ VPWR VPWR _04527_ sky130_fd_sc_hd__mux2_1
X_17799_ net879 _01361_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09222_ CPU.Iimm\[2\] CPU.Bimm\[2\] CPU.instr\[5\] VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09153_ _05396_ _05503_ _05504_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09084_ _05277_ _05244_ _05278_ _05279_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold820 CPU.registerFile\[17\]\[22\] VGND VGND VPWR VPWR net2117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold831 CPU.registerFile\[23\]\[18\] VGND VGND VPWR VPWR net2128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 CPU.registerFile\[26\]\[29\] VGND VGND VPWR VPWR net2139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 CPU.registerFile\[5\]\[25\] VGND VGND VPWR VPWR net2150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold864 CPU.registerFile\[18\]\[1\] VGND VGND VPWR VPWR net2161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 CPU.registerFile\[15\]\[19\] VGND VGND VPWR VPWR net2172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold886 CPU.registerFile\[8\]\[30\] VGND VGND VPWR VPWR net2183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold897 mapped_spi_flash.rcv_data\[1\] VGND VGND VPWR VPWR net2194 sky130_fd_sc_hd__dlygate4sd3_1
X_09986_ net2333 _06316_ _06293_ VGND VGND VPWR VPWR _06317_ sky130_fd_sc_hd__mux2_1
X_13767__1134 clknet_1_1__leaf__08461_ VGND VGND VPWR VPWR net1190 sky130_fd_sc_hd__inv_2
X_08937_ CPU.aluIn1\[4\] _05287_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__nor2_1
X_14151__290 clknet_1_1__leaf__08499_ VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__inv_2
XFILLER_0_98_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10830_ CPU.aluReg\[19\] _06911_ _06889_ VGND VGND VPWR VPWR _06912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10761_ net1625 _06851_ _06852_ _06856_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12500_ _07937_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13480_ _08431_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__clkbuf_1
X_10692_ _06818_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12431_ net1925 _07343_ _07895_ VGND VGND VPWR VPWR _07901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15150_ _08409_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__buf_4
XFILLER_0_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12362_ _07864_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__clkbuf_1
X_11313_ net1903 _06106_ _07249_ VGND VGND VPWR VPWR _07252_ sky130_fd_sc_hd__mux2_1
X_15081_ CPU.registerFile\[5\]\[18\] CPU.registerFile\[4\]\[18\] _03105_ VGND VGND
+ VPWR VPWR _03145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12293_ _07163_ VGND VGND VPWR VPWR _07822_ sky130_fd_sc_hd__buf_4
XFILLER_0_160_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11244_ _06622_ net2130 _07212_ VGND VGND VPWR VPWR _07215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18840_ clknet_leaf_7_clk _02364_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11175_ net1338 _07134_ VGND VGND VPWR VPWR _07171_ sky130_fd_sc_hd__or2_1
X_10126_ _06450_ _05961_ VGND VGND VPWR VPWR _06451_ sky130_fd_sc_hd__xnor2_1
X_18771_ net560 _02295_ VGND VGND VPWR VPWR CPU.aluReg\[1\] sky130_fd_sc_hd__dfxtp_1
X_15983_ CPU.registerFile\[13\]\[0\] _03709_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__or2_1
X_17722_ clknet_leaf_2_clk _01288_ VGND VGND VPWR VPWR CPU.PC\[1\] sky130_fd_sc_hd__dfxtp_1
X_10057_ _06176_ _06367_ _06384_ VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__a21o_2
X_14934_ CPU.registerFile\[20\]\[15\] _08839_ _03000_ _08841_ VGND VGND VPWR VPWR
+ _03001_ sky130_fd_sc_hd__o211a_1
X_17653_ per_uart.uart0.rx_count16\[1\] per_uart.uart0.rx_count16\[0\] _05185_ per_uart.uart0.rx_count16\[2\]
+ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__a31oi_1
X_14865_ CPU.registerFile\[15\]\[13\] CPU.registerFile\[14\]\[13\] _08771_ VGND VGND
+ VPWR VPWR _02934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16604_ _04315_ _04316_ _04279_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__mux2_1
X_17584_ _05120_ _05125_ _05144_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__mux2_1
X_14796_ _02728_ _02861_ _02866_ _02784_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16535_ _04248_ _04249_ _03961_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__mux2_1
X_10959_ _07008_ _07010_ VGND VGND VPWR VPWR _07011_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16466_ _04141_ _04160_ _04182_ _04096_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__a211o_1
X_13613__995 clknet_1_0__leaf__08446_ VGND VGND VPWR VPWR net1051 sky130_fd_sc_hd__inv_2
XFILLER_0_6_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18205_ net1216 net1350 VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[6\] sky130_fd_sc_hd__dfxtp_1
X_15417_ CPU.registerFile\[27\]\[27\] CPU.registerFile\[26\]\[27\] _03172_ VGND VGND
+ VPWR VPWR _03472_ sky130_fd_sc_hd__mux2_1
X_12629_ _08006_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__clkbuf_1
X_19185_ clknet_leaf_3_clk _02703_ VGND VGND VPWR VPWR per_uart.d_in_uart\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16397_ _03985_ _03986_ CPU.registerFile\[1\]\[9\] VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18136_ net1147 _01664_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_15348_ _08580_ _03402_ _03404_ _03218_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__a211o_1
XFILLER_0_130_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13827__1188 clknet_1_0__leaf__08467_ VGND VGND VPWR VPWR net1244 sky130_fd_sc_hd__inv_2
X_18067_ net1078 _01595_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[9\] sky130_fd_sc_hd__dfxtp_1
Xhold105 _05804_ VGND VGND VPWR VPWR net1402 sky130_fd_sc_hd__buf_1
X_15279_ CPU.registerFile\[13\]\[23\] CPU.registerFile\[12\]\[23\] _08794_ VGND VGND
+ VPWR VPWR _03338_ sky130_fd_sc_hd__mux2_1
X_13386__879 clknet_1_0__leaf__08370_ VGND VGND VPWR VPWR net935 sky130_fd_sc_hd__inv_2
Xhold116 _01745_ VGND VGND VPWR VPWR net1413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 mapped_spi_ram.cmd_addr\[22\] VGND VGND VPWR VPWR net1424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 mapped_spi_ram.rcv_data\[28\] VGND VGND VPWR VPWR net1435 sky130_fd_sc_hd__dlygate4sd3_1
X_17018_ CPU.registerFile\[24\]\[24\] _03724_ _04569_ _04720_ VGND VGND VPWR VPWR
+ _04721_ sky130_fd_sc_hd__o211a_1
Xhold149 mapped_spi_flash.rcv_bitcount\[4\] VGND VGND VPWR VPWR net1446 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__03656_ clknet_0__03656_ VGND VGND VPWR VPWR clknet_1_1__leaf__03656_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ _05730_ VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__clkbuf_4
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__03687_ _03687_ VGND VGND VPWR VPWR clknet_0__03687_ sky130_fd_sc_hd__clkbuf_16
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _05856_ _06109_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18969_ net743 _02489_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09205_ CPU.state\[3\] CPU.state\[2\] VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13588__972 clknet_1_0__leaf__08444_ VGND VGND VPWR VPWR net1028 sky130_fd_sc_hd__inv_2
XFILLER_0_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09136_ _05487_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09067_ CPU.aluIn1\[31\] _05416_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold650 CPU.registerFile\[11\]\[9\] VGND VGND VPWR VPWR net1947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 CPU.registerFile\[15\]\[9\] VGND VGND VPWR VPWR net1958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 CPU.registerFile\[22\]\[25\] VGND VGND VPWR VPWR net1969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 CPU.registerFile\[15\]\[1\] VGND VGND VPWR VPWR net1980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 CPU.registerFile\[7\]\[13\] VGND VGND VPWR VPWR net1991 sky130_fd_sc_hd__dlygate4sd3_1
X_09969_ _05794_ _06299_ VGND VGND VPWR VPWR _06300_ sky130_fd_sc_hd__or2_1
X_13844__1203 clknet_1_0__leaf__08469_ VGND VGND VPWR VPWR net1259 sky130_fd_sc_hd__inv_2
X_12980_ _08193_ VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__clkbuf_1
Xhold1350 CPU.aluReg\[3\] VGND VGND VPWR VPWR net2647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1361 CPU.aluIn1\[4\] VGND VGND VPWR VPWR net2658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1372 CPU.aluReg\[12\] VGND VGND VPWR VPWR net2669 sky130_fd_sc_hd__dlygate4sd3_1
X_11931_ _07595_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__clkbuf_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ CPU.registerFile\[24\]\[8\] _08686_ _02723_ _08550_ VGND VGND VPWR VPWR _02724_
+ sky130_fd_sc_hd__o211a_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ net1931 _07374_ _07525_ VGND VGND VPWR VPWR _07559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10813_ CPU.aluReg\[23\] _06898_ _06889_ VGND VGND VPWR VPWR _06899_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _08520_ _08818_ _08820_ _08661_ VGND VGND VPWR VPWR _08821_ sky130_fd_sc_hd__a211o_1
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _07522_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__clkbuf_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_914 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16320_ CPU.registerFile\[24\]\[7\] _03915_ _03747_ _04039_ VGND VGND VPWR VPWR _04040_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10744_ _06845_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__clkbuf_1
X_17305__720 clknet_1_1__leaf__04980_ VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__inv_2
X_15663__461 clknet_1_0__leaf__03644_ VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__inv_2
X_16251_ CPU.registerFile\[9\]\[6\] _03698_ VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__or2_1
X_13463_ _08421_ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__clkbuf_1
X_10675_ _06807_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__clkbuf_1
X_15202_ CPU.registerFile\[15\]\[21\] CPU.registerFile\[14\]\[21\] _03013_ VGND VGND
+ VPWR VPWR _03263_ sky130_fd_sc_hd__mux2_1
X_12414_ net1823 _07326_ _07884_ VGND VGND VPWR VPWR _07892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16182_ CPU.registerFile\[2\]\[4\] CPU.registerFile\[3\]\[4\] _03693_ VGND VGND VPWR
+ VPWR _03905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13394_ _05856_ _06395_ _08372_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__o21a_1
XFILLER_0_152_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15133_ CPU.registerFile\[0\]\[19\] _02948_ _03194_ _03195_ VGND VGND VPWR VPWR _03196_
+ sky130_fd_sc_hd__o211a_1
X_12345_ _07855_ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__clkbuf_1
X_15064_ _03049_ _03050_ CPU.registerFile\[25\]\[18\] VGND VGND VPWR VPWR _03128_
+ sky130_fd_sc_hd__a21o_1
X_12276_ _07784_ VGND VGND VPWR VPWR _07812_ sky130_fd_sc_hd__buf_2
XFILLER_0_120_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14158__296 clknet_1_0__leaf__08500_ VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__inv_2
XFILLER_0_120_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11227_ _06605_ net1788 _07201_ VGND VGND VPWR VPWR _07206_ sky130_fd_sc_hd__mux2_1
X_18823_ net612 _02347_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11158_ net1419 _07160_ _07161_ _07151_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__o211a_1
X_10109_ _05284_ _05285_ _05769_ _05770_ net1862 VGND VGND VPWR VPWR _06435_ sky130_fd_sc_hd__a32o_1
X_15966_ _06172_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__clkbuf_8
X_11089_ _06973_ _06985_ _07117_ _07114_ net1588 VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__a32o_1
X_18754_ net543 _02278_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[16\] sky130_fd_sc_hd__dfxtp_1
X_14917_ _02983_ _02984_ _08783_ VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__mux2_1
X_17705_ _05207_ _05227_ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__and2_1
X_18685_ net474 _02209_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17636_ per_uart.rx_data\[7\] net2631 _05170_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__mux2_1
X_14848_ CPU.registerFile\[17\]\[13\] _08795_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15746__536 clknet_1_0__leaf__03652_ VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__inv_2
X_17567_ per_uart.uart0.tx_count16\[1\] per_uart.uart0.tx_count16\[0\] VGND VGND VPWR
+ VPWR _05131_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14779_ CPU.registerFile\[28\]\[11\] CPU.registerFile\[29\]\[11\] _02808_ VGND VGND
+ VPWR VPWR _02850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16518_ _06172_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17498_ _05075_ _05017_ _06219_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_74_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13766__1133 clknet_1_1__leaf__08461_ VGND VGND VPWR VPWR net1189 sky130_fd_sc_hd__inv_2
X_16449_ _04080_ _04081_ CPU.registerFile\[25\]\[10\] VGND VGND VPWR VPWR _04166_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19168_ clknet_leaf_0_clk _02688_ VGND VGND VPWR VPWR per_uart.rx_data\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18119_ net1130 _01647_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19099_ net82 _02619_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03639_ clknet_0__03639_ VGND VGND VPWR VPWR clknet_1_1__leaf__03639_
+ sky130_fd_sc_hd__clkbuf_16
X_09823_ _06017_ _06159_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__nand2_1
X_09754_ _05477_ _06093_ _05480_ VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__a21o_1
X_09685_ _06005_ _05918_ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__and2b_1
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14263__391 clknet_1_0__leaf__08510_ VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__inv_2
XFILLER_0_92_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10460_ _06647_ net2002 _06687_ VGND VGND VPWR VPWR _06692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13369__863 clknet_1_0__leaf__08369_ VGND VGND VPWR VPWR net919 sky130_fd_sc_hd__inv_2
X_09119_ _05333_ _05469_ _05470_ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_150_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10391_ _06652_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__clkbuf_1
X_12130_ _07692_ VGND VGND VPWR VPWR _07714_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12061_ CPU.registerFile\[24\]\[4\] _07368_ _07657_ VGND VGND VPWR VPWR _07665_ sky130_fd_sc_hd__mux2_1
Xhold480 CPU.registerFile\[15\]\[22\] VGND VGND VPWR VPWR net1777 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold491 CPU.registerFile\[30\]\[27\] VGND VGND VPWR VPWR net1788 sky130_fd_sc_hd__dlygate4sd3_1
X_11012_ _06999_ VGND VGND VPWR VPWR _07054_ sky130_fd_sc_hd__buf_2
XFILLER_0_35_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12963_ _08184_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__clkbuf_1
Xhold1180 CPU.registerFile\[20\]\[0\] VGND VGND VPWR VPWR net2477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 CPU.registerFile\[1\]\[11\] VGND VGND VPWR VPWR net2488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14702_ _08515_ _02760_ _02764_ _02774_ VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__a31o_1
X_18470_ net291 _01994_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11914_ _06643_ net2125 _07584_ VGND VGND VPWR VPWR _07587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13826__1187 clknet_1_0__leaf__08467_ VGND VGND VPWR VPWR net1243 sky130_fd_sc_hd__inv_2
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _05786_ net2114 _08145_ VGND VGND VPWR VPWR _08148_ sky130_fd_sc_hd__mux2_1
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _08574_ _08866_ _08871_ _08592_ VGND VGND VPWR VPWR _08872_ sky130_fd_sc_hd__o211a_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11845_ _07550_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__clkbuf_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ CPU.registerFile\[30\]\[6\] CPU.registerFile\[31\]\[6\] _08645_ VGND VGND
+ VPWR VPWR _08804_ sky130_fd_sc_hd__mux2_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _06641_ net1916 _07512_ VGND VGND VPWR VPWR _07514_ sky130_fd_sc_hd__mux2_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16303_ CPU.registerFile\[6\]\[7\] CPU.registerFile\[7\]\[7\] _04022_ VGND VGND VPWR
+ VPWR _04023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10727_ _06836_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__clkbuf_1
X_17283_ CPU.aluIn1\[31\] _08513_ _04978_ _04663_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__o211a_1
X_14495_ CPU.registerFile\[8\]\[4\] _08526_ _08736_ _08622_ VGND VGND VPWR VPWR _08737_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19022_ net764 _02542_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_16234_ _03702_ _03953_ _03955_ _03803_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13446_ _08407_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__clkbuf_1
X_10658_ _06798_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16165_ _03766_ _03886_ _03888_ _06142_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10589_ _06738_ VGND VGND VPWR VPWR _06761_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15116_ _02798_ _03164_ _03168_ _03178_ VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__a31o_1
X_12328_ _07838_ net1303 mapped_spi_ram.rcv_bitcount\[0\] VGND VGND VPWR VPWR _07846_
+ sky130_fd_sc_hd__mux2_1
X_16096_ CPU.registerFile\[13\]\[2\] _03709_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__or2_1
X_15047_ _03027_ _03108_ _03110_ _03111_ VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__a211o_1
X_14091__236 clknet_1_1__leaf__08493_ VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__inv_2
X_12259_ mapped_spi_ram.rcv_data\[19\] _07800_ VGND VGND VPWR VPWR _07803_ sky130_fd_sc_hd__or2_1
X_18806_ net595 _02330_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_16998_ CPU.registerFile\[8\]\[24\] _04505_ _04506_ _04700_ VGND VGND VPWR VPWR _04701_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18737_ net526 _02261_ VGND VGND VPWR VPWR mapped_spi_flash.snd_bitcount\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09470_ _05517_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__clkbuf_4
X_18668_ net457 _02192_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_17619_ _03659_ _04989_ _04990_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__nor3_2
X_18599_ net420 _02123_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13843__1202 clknet_1_0__leaf__08469_ VGND VGND VPWR VPWR net1258 sky130_fd_sc_hd__inv_2
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09806_ _05745_ _06134_ _06139_ _06143_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__a211o_2
XFILLER_0_157_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13260__780 clknet_1_0__leaf__08344_ VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__inv_2
X_09737_ CPU.Iimm\[0\] _05550_ _05790_ CPU.cycles\[20\] _06077_ VGND VGND VPWR VPWR
+ _06078_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09668_ _06011_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__clkbuf_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ CPU.PC\[11\] _05942_ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__or2_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _07435_ VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__clkbuf_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11561_ _07398_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13300_ clknet_1_1__leaf__08341_ VGND VGND VPWR VPWR _08362_ sky130_fd_sc_hd__buf_1
X_10512_ net1905 _06200_ _06713_ VGND VGND VPWR VPWR _06720_ sky130_fd_sc_hd__mux2_1
X_14280_ _08525_ VGND VGND VPWR VPWR _08526_ sky130_fd_sc_hd__clkbuf_8
X_11492_ _07357_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10443_ _06630_ net2555 _06676_ VGND VGND VPWR VPWR _06683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13162_ _08289_ net1539 VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__nor2_1
X_10374_ _06315_ VGND VGND VPWR VPWR _06641_ sky130_fd_sc_hd__buf_4
X_12113_ net1316 _07694_ _07696_ VGND VGND VPWR VPWR _07702_ sky130_fd_sc_hd__a21o_1
X_17970_ net981 _01498_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_13093_ CPU.mem_wbusy _06861_ _08252_ VGND VGND VPWR VPWR _08253_ sky130_fd_sc_hd__or3b_1
X_16921_ CPU.registerFile\[9\]\[22\] _04460_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__or2_1
X_12044_ CPU.registerFile\[24\]\[12\] _07351_ _07646_ VGND VGND VPWR VPWR _07656_
+ sky130_fd_sc_hd__mux2_1
X_16852_ CPU.registerFile\[2\]\[20\] CPU.registerFile\[3\]\[20\] _04431_ VGND VGND
+ VPWR VPWR _04559_ sky130_fd_sc_hd__mux2_1
X_13765__1132 clknet_1_0__leaf__08461_ VGND VGND VPWR VPWR net1188 sky130_fd_sc_hd__inv_2
X_15803_ net1596 _08351_ net1610 VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__o21ai_1
X_16783_ _04490_ _04491_ _04365_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__mux2_1
X_18522_ net343 _02046_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_12946_ _06465_ net2334 _08167_ VGND VGND VPWR VPWR _08175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18453_ net274 _01981_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12877_ _08138_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__clkbuf_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14616_ CPU.registerFile\[13\]\[7\] CPU.registerFile\[12\]\[7\] _08693_ VGND VGND
+ VPWR VPWR _08855_ sky130_fd_sc_hd__mux2_1
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _07541_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__clkbuf_1
X_18384_ net205 _01912_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ CPU.registerFile\[0\]\[5\] _08706_ _08787_ _08588_ VGND VGND VPWR VPWR _08788_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11759_ _06624_ net2539 _07501_ VGND VGND VPWR VPWR _07505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15858__604 clknet_1_0__leaf__03681_ VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__08500_ clknet_0__08500_ VGND VGND VPWR VPWR clknet_1_1__leaf__08500_
+ sky130_fd_sc_hd__clkbuf_16
X_17266_ CPU.registerFile\[28\]\[31\] CPU.registerFile\[29\]\[31\] _03717_ VGND VGND
+ VPWR VPWR _04962_ sky130_fd_sc_hd__mux2_1
X_14478_ CPU.registerFile\[20\]\[4\] _08527_ _08719_ _08530_ VGND VGND VPWR VPWR _08720_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16217_ _03703_ _03936_ _03938_ _03714_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19005_ clknet_leaf_12_clk _02525_ VGND VGND VPWR VPWR CPU.aluIn1\[22\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_52_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13429_ CPU.Jimm\[15\] _08394_ _08388_ VGND VGND VPWR VPWR _08395_ sky130_fd_sc_hd__mux2_1
X_17197_ _03726_ _03727_ CPU.registerFile\[25\]\[29\] VGND VGND VPWR VPWR _04895_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__08462_ _08462_ VGND VGND VPWR VPWR clknet_0__08462_ sky130_fd_sc_hd__clkbuf_16
X_16148_ _08404_ _03859_ _03863_ _03871_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__a31o_2
Xclkbuf_1_1__f__08362_ clknet_0__08362_ VGND VGND VPWR VPWR clknet_1_1__leaf__08362_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13956__114 clknet_1_0__leaf__08480_ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__inv_2
XFILLER_0_121_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16079_ _03735_ _03799_ _03804_ _03755_ VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__o211a_1
X_08970_ CPU.rs2\[13\] _05245_ _05249_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__o21a_1
Xinput1 RXD VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09522_ _05389_ _05748_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09453_ _05792_ _05801_ _05744_ VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__o21a_1
X_13552__941 clknet_1_1__leaf__08439_ VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__inv_2
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09384_ CPU.Bimm\[11\] VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__buf_4
XFILLER_0_74_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13825__1186 clknet_1_0__leaf__08467_ VGND VGND VPWR VPWR net1242 sky130_fd_sc_hd__inv_2
XFILLER_0_100_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10090_ net1366 _05860_ _05719_ per_uart.rx_data\[5\] _06415_ VGND VGND VPWR VPWR
+ _06416_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__08451_ clknet_0__08451_ VGND VGND VPWR VPWR clknet_1_0__leaf__08451_
+ sky130_fd_sc_hd__clkbuf_16
X_12800_ _08096_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__clkbuf_1
X_10992_ CPU.PC\[14\] _07031_ VGND VGND VPWR VPWR _07037_ sky130_fd_sc_hd__or2_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _06655_ net2646 _08051_ VGND VGND VPWR VPWR _08060_ sky130_fd_sc_hd__mux2_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ CPU.registerFile\[30\]\[28\] CPU.registerFile\[31\]\[28\] _03291_ VGND VGND
+ VPWR VPWR _03504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _08023_ VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__clkbuf_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _08409_ VGND VGND VPWR VPWR _08645_ sky130_fd_sc_hd__buf_4
XFILLER_0_38_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11613_ _07426_ VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__clkbuf_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15381_ CPU.registerFile\[27\]\[26\] CPU.registerFile\[26\]\[26\] _03172_ VGND VGND
+ VPWR VPWR _03437_ sky130_fd_sc_hd__mux2_1
X_12593_ net2600 _07368_ _07979_ VGND VGND VPWR VPWR _07987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17120_ _04502_ _04807_ _04811_ _04819_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__a31o_2
X_14332_ _08540_ VGND VGND VPWR VPWR _08578_ sky130_fd_sc_hd__clkbuf_8
X_11544_ _07389_ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17051_ _04751_ _04752_ _06535_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11475_ net1808 _07345_ _07333_ VGND VGND VPWR VPWR _07346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16002_ CPU.registerFile\[0\]\[0\] _03724_ _03725_ _03728_ VGND VGND VPWR VPWR _03729_
+ sky130_fd_sc_hd__o211a_1
X_15699__493 clknet_1_0__leaf__03648_ VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__inv_2
X_13214_ _05526_ _06544_ VGND VGND VPWR VPWR _08328_ sky130_fd_sc_hd__xnor2_1
X_10426_ _06613_ net2455 _06665_ VGND VGND VPWR VPWR _06674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13145_ net1613 _08279_ VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__xor2_1
X_10357_ _06629_ VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__clkbuf_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ CPU.registerFile\[4\]\[7\] net1399 _08239_ VGND VGND VPWR VPWR _08244_ sky130_fd_sc_hd__mux2_1
X_17953_ net964 _01481_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_10288_ _06584_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__clkbuf_1
X_12027_ _07647_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__clkbuf_1
X_16904_ _04484_ _04485_ CPU.registerFile\[25\]\[21\] VGND VGND VPWR VPWR _04610_
+ sky130_fd_sc_hd__a21o_1
X_17884_ clknet_leaf_20_clk _00034_ VGND VGND VPWR VPWR CPU.cycles\[27\] sky130_fd_sc_hd__dfxtp_1
X_16835_ _04533_ _04541_ _04542_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__o21a_1
X_16766_ _04347_ _04471_ _04474_ _04117_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__a211o_1
XFILLER_0_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18505_ net326 _02029_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_12929_ _06267_ net2265 _08156_ VGND VGND VPWR VPWR _08166_ sky130_fd_sc_hd__mux2_1
X_16697_ _04175_ _04176_ CPU.registerFile\[17\]\[16\] VGND VGND VPWR VPWR _04408_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18436_ net257 _01964_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18367_ net188 _01895_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_15579_ _03628_ _03629_ _08562_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17318_ clknet_1_1__leaf__03686_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__buf_1
X_18298_ net119 _01826_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17249_ CPU.registerFile\[9\]\[31\] _03709_ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__or2_1
X_14023__174 clknet_1_0__leaf__08487_ VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__inv_2
XFILLER_0_113_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13582__967 clknet_1_1__leaf__08443_ VGND VGND VPWR VPWR net1023 sky130_fd_sc_hd__inv_2
XFILLER_0_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__08445_ _08445_ VGND VGND VPWR VPWR clknet_0__08445_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__08345_ clknet_0__08345_ VGND VGND VPWR VPWR clknet_1_1__leaf__08345_
+ sky130_fd_sc_hd__clkbuf_16
X_08953_ _05299_ _05303_ _05304_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08884_ mapped_spi_ram.div_counter\[3\] mapped_spi_ram.div_counter\[2\] mapped_spi_ram.div_counter\[5\]
+ mapped_spi_ram.div_counter\[4\] VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__or4_2
XFILLER_0_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15611__414 clknet_1_1__leaf__03639_ VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__inv_2
XFILLER_0_154_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09505_ _05731_ _05842_ _05850_ _05541_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09436_ _05785_ VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__clkbuf_4
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09367_ _05718_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_50 clknet_1_1__leaf__03640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09298_ _05643_ _05649_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_61 clknet_1_0__leaf__08341_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _07464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_83 _06123_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11260_ _07200_ VGND VGND VPWR VPWR _07223_ sky130_fd_sc_hd__buf_4
XFILLER_0_31_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10211_ per_uart.rx_data\[0\] _05719_ VGND VGND VPWR VPWR _06532_ sky130_fd_sc_hd__and2_1
X_11191_ _07009_ _07181_ VGND VGND VPWR VPWR _07182_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10142_ _06466_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__clkbuf_1
X_14950_ CPU.registerFile\[10\]\[15\] CPU.registerFile\[11\]\[15\] _02779_ VGND VGND
+ VPWR VPWR _03017_ sky130_fd_sc_hd__mux2_1
X_10073_ _06399_ _05965_ VGND VGND VPWR VPWR _06400_ sky130_fd_sc_hd__xnor2_1
X_14881_ CPU.registerFile\[0\]\[13\] _02948_ _02949_ _02791_ VGND VGND VPWR VPWR _02950_
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_0__f__08503_ clknet_0__08503_ VGND VGND VPWR VPWR clknet_1_0__leaf__08503_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16620_ _04323_ _04332_ _04138_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__o21a_1
Xclkbuf_1_0__f__08434_ clknet_0__08434_ VGND VGND VPWR VPWR clknet_1_0__leaf__08434_
+ sky130_fd_sc_hd__clkbuf_16
X_16551_ CPU.registerFile\[13\]\[13\] _03976_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13890__54 clknet_1_0__leaf__08474_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__inv_2
X_10975_ _07008_ _07021_ VGND VGND VPWR VPWR _07022_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_0__f__08365_ clknet_0__08365_ VGND VGND VPWR VPWR clknet_1_0__leaf__08365_
+ sky130_fd_sc_hd__clkbuf_16
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15502_ _08533_ _03550_ _03554_ _08554_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__o211a_1
X_12714_ _08028_ VGND VGND VPWR VPWR _08051_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16482_ _03943_ _04195_ _04197_ _04117_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15433_ _03486_ _03487_ _08562_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__mux2_1
X_18221_ net1232 _01749_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12645_ _08014_ VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18152_ net1163 _01680_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_15364_ CPU.registerFile\[0\]\[25\] _08411_ _03420_ _03195_ VGND VGND VPWR VPWR _03421_
+ sky130_fd_sc_hd__o211a_1
X_12576_ net2597 _07351_ _07968_ VGND VGND VPWR VPWR _07978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14315_ CPU.registerFile\[13\]\[0\] CPU.registerFile\[12\]\[0\] _08560_ VGND VGND
+ VPWR VPWR _08561_ sky130_fd_sc_hd__mux2_1
X_17103_ net2617 _04458_ _04803_ _04663_ VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__o211a_1
X_11527_ net1676 _07314_ _07379_ VGND VGND VPWR VPWR _07381_ sky130_fd_sc_hd__mux2_1
X_18083_ net1094 _01611_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_15295_ _03155_ _03336_ _03353_ _03243_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__a211o_2
XFILLER_0_151_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17034_ CPU.registerFile\[8\]\[25\] _04505_ _04506_ _04735_ VGND VGND VPWR VPWR _04736_
+ sky130_fd_sc_hd__o211a_1
Xhold309 CPU.cycles\[26\] VGND VGND VPWR VPWR net1606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11458_ _07334_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10409_ _06664_ VGND VGND VPWR VPWR _06665_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11389_ net1814 _06200_ _07285_ VGND VGND VPWR VPWR _07292_ sky130_fd_sc_hd__mux2_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ CPU.cycles\[3\] _08269_ VGND VGND VPWR VPWR _08271_ sky130_fd_sc_hd__and2_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ clknet_leaf_18_clk _02505_ VGND VGND VPWR VPWR CPU.aluIn1\[2\] sky130_fd_sc_hd__dfxtp_4
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ CPU.registerFile\[4\]\[15\] _06199_ _08228_ VGND VGND VPWR VPWR _08235_ sky130_fd_sc_hd__mux2_1
X_17936_ net947 _01464_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold1009 CPU.registerFile\[3\]\[12\] VGND VGND VPWR VPWR net2306 sky130_fd_sc_hd__dlygate4sd3_1
X_13686__1061 clknet_1_1__leaf__08453_ VGND VGND VPWR VPWR net1117 sky130_fd_sc_hd__inv_2
X_14211__344 clknet_1_0__leaf__08505_ VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__inv_2
XFILLER_0_84_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17867_ clknet_leaf_24_clk _00016_ VGND VGND VPWR VPWR CPU.cycles\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16818_ _06171_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__buf_4
X_17798_ net878 _01360_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16749_ _08513_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13824__1185 clknet_1_1__leaf__08467_ VGND VGND VPWR VPWR net1241 sky130_fd_sc_hd__inv_2
XFILLER_0_124_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09221_ CPU.aluIn1\[3\] _05572_ VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__or2_1
X_18419_ net240 _01947_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09152_ _05392_ CPU.aluIn1\[27\] VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__and2b_1
XFILLER_0_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09083_ _05279_ _05434_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold810 CPU.registerFile\[13\]\[22\] VGND VGND VPWR VPWR net2107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold821 CPU.registerFile\[26\]\[26\] VGND VGND VPWR VPWR net2118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 CPU.registerFile\[27\]\[2\] VGND VGND VPWR VPWR net2129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 CPU.registerFile\[8\]\[16\] VGND VGND VPWR VPWR net2140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 CPU.registerFile\[18\]\[6\] VGND VGND VPWR VPWR net2151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 CPU.registerFile\[11\]\[3\] VGND VGND VPWR VPWR net2162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold876 CPU.registerFile\[16\]\[14\] VGND VGND VPWR VPWR net2173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 CPU.registerFile\[15\]\[0\] VGND VGND VPWR VPWR net2184 sky130_fd_sc_hd__dlygate4sd3_1
X_15836__584 clknet_1_0__leaf__03679_ VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__inv_2
X_13363__858 clknet_1_1__leaf__08368_ VGND VGND VPWR VPWR net914 sky130_fd_sc_hd__inv_2
Xhold898 CPU.registerFile\[14\]\[24\] VGND VGND VPWR VPWR net2195 sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ _06315_ VGND VGND VPWR VPWR _06316_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08936_ CPU.aluIn1\[4\] _05287_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10760_ _06855_ VGND VGND VPWR VPWR _06856_ sky130_fd_sc_hd__buf_4
XFILLER_0_137_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09419_ _05532_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10691_ net1988 _05767_ _06816_ VGND VGND VPWR VPWR _06818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12430_ _07900_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12361_ _06626_ net1897 _07859_ VGND VGND VPWR VPWR _07864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11312_ _07251_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15080_ CPU.registerFile\[6\]\[18\] CPU.registerFile\[7\]\[18\] _02982_ VGND VGND
+ VPWR VPWR _03144_ sky130_fd_sc_hd__mux2_1
X_15919__659 clknet_1_0__leaf__03687_ VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__inv_2
X_12292_ mapped_spi_ram.rcv_data\[4\] _07813_ VGND VGND VPWR VPWR _07821_ sky130_fd_sc_hd__or2_1
X_13927__88 clknet_1_1__leaf__08477_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__inv_2
XFILLER_0_105_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14031_ clknet_1_1__leaf__08484_ VGND VGND VPWR VPWR _08488_ sky130_fd_sc_hd__buf_1
X_11243_ _07214_ VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11174_ net1338 _07160_ _07170_ _07164_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10125_ _05962_ _05951_ VGND VGND VPWR VPWR _06450_ sky130_fd_sc_hd__and2b_1
X_18770_ net559 _02294_ VGND VGND VPWR VPWR CPU.aluReg\[0\] sky130_fd_sc_hd__dfxtp_1
X_15982_ _03697_ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__buf_2
X_10056_ CPU.cycles\[7\] _05759_ _06368_ _06370_ _06383_ VGND VGND VPWR VPWR _06384_
+ sky130_fd_sc_hd__a221o_1
X_14933_ CPU.registerFile\[21\]\[15\] _02960_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17652_ per_uart.uart0.rx_count16\[2\] per_uart.uart0.rx_count16\[1\] per_uart.uart0.rx_count16\[0\]
+ _05185_ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__and4_1
X_14864_ _02798_ _02919_ _02923_ _02932_ VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__a31o_1
X_16603_ CPU.registerFile\[28\]\[14\] CPU.registerFile\[29\]\[14\] _04122_ VGND VGND
+ VPWR VPWR _04316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14795_ _08857_ _02862_ _02865_ _08661_ VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__a211o_1
X_17583_ per_uart.uart0.tx_bitcount\[0\] _05133_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16534_ CPU.registerFile\[20\]\[12\] CPU.registerFile\[21\]\[12\] _03883_ VGND VGND
+ VPWR VPWR _04249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10958_ net1520 _05638_ _07009_ VGND VGND VPWR VPWR _07010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16465_ _04169_ _04181_ _04138_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10889_ net1862 _06956_ _06868_ VGND VGND VPWR VPWR _06957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18204_ net1215 _01732_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[5\] sky130_fd_sc_hd__dfxtp_1
X_12628_ _06620_ net2012 _08004_ VGND VGND VPWR VPWR _08006_ sky130_fd_sc_hd__mux2_1
X_15416_ _03469_ _03470_ _03255_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16396_ CPU.registerFile\[2\]\[9\] CPU.registerFile\[3\]\[9\] _04027_ VGND VGND VPWR
+ VPWR _04114_ sky130_fd_sc_hd__mux2_1
X_19184_ clknet_leaf_3_clk _02702_ VGND VGND VPWR VPWR per_uart.uart0.tx_wr sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18135_ net1146 _01663_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15347_ CPU.registerFile\[24\]\[25\] _08582_ _03403_ _03175_ VGND VGND VPWR VPWR
+ _03404_ sky130_fd_sc_hd__o211a_1
X_12559_ _07969_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15278_ CPU.registerFile\[15\]\[23\] CPU.registerFile\[14\]\[23\] _03013_ VGND VGND
+ VPWR VPWR _03337_ sky130_fd_sc_hd__mux2_1
X_18066_ net1077 _01594_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xhold106 _08221_ VGND VGND VPWR VPWR net1403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold117 CPU.aluReg\[15\] VGND VGND VPWR VPWR net1414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 mapped_spi_ram.cmd_addr\[23\] VGND VGND VPWR VPWR net1425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold139 _01718_ VGND VGND VPWR VPWR net1436 sky130_fd_sc_hd__dlygate4sd3_1
X_17017_ _04484_ _04485_ CPU.registerFile\[25\]\[24\] VGND VGND VPWR VPWR _04720_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03655_ clknet_0__03655_ VGND VGND VPWR VPWR clknet_1_1__leaf__03655_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__03686_ _03686_ VGND VGND VPWR VPWR clknet_0__03686_ sky130_fd_sc_hd__clkbuf_16
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14135__275 clknet_1_0__leaf__08498_ VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__inv_2
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _06108_ VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__clkbuf_8
X_18968_ net742 _02488_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ clknet_leaf_26_clk _01447_ VGND VGND VPWR VPWR CPU.Bimm\[6\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18899_ net673 _02419_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15723__515 clknet_1_0__leaf__03650_ VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__inv_2
X_14029__180 clknet_1_1__leaf__08487_ VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__inv_2
XFILLER_0_17_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09204_ _05555_ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09135_ _05380_ _05369_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__or2_1
XFILLER_0_162_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09066_ _05417_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold640 CPU.registerFile\[13\]\[28\] VGND VGND VPWR VPWR net1937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold651 CPU.registerFile\[2\]\[4\] VGND VGND VPWR VPWR net1948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold662 per_uart.rx_data\[4\] VGND VGND VPWR VPWR net1959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 CPU.registerFile\[17\]\[4\] VGND VGND VPWR VPWR net1970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 CPU.registerFile\[2\]\[29\] VGND VGND VPWR VPWR net1981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold695 CPU.registerFile\[21\]\[5\] VGND VGND VPWR VPWR net1992 sky130_fd_sc_hd__dlygate4sd3_1
X_15617__420 clknet_1_0__leaf__03639_ VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__inv_2
X_09968_ _05311_ _06298_ VGND VGND VPWR VPWR _06299_ sky130_fd_sc_hd__nor2_1
X_08919_ CPU.aluIn1\[2\] _05270_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09899_ _05818_ _06228_ _06231_ _06232_ _05335_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__a32o_1
Xhold1340 CPU.registerFile\[1\]\[5\] VGND VGND VPWR VPWR net2637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1351 CPU.registerFile\[1\]\[23\] VGND VGND VPWR VPWR net2648 sky130_fd_sc_hd__dlygate4sd3_1
X_11930_ _06659_ net2391 _07561_ VGND VGND VPWR VPWR _07595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1362 CPU.PC\[1\] VGND VGND VPWR VPWR net2659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1373 CPU.aluReg\[15\] VGND VGND VPWR VPWR net2670 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _07558_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__clkbuf_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ CPU.aluIn1\[23\] _06897_ _06881_ VGND VGND VPWR VPWR _06898_ sky130_fd_sc_hd__mux2_1
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14580_ CPU.registerFile\[8\]\[6\] _08776_ _08819_ _08622_ VGND VGND VPWR VPWR _08820_
+ sky130_fd_sc_hd__o211a_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _06657_ net2067 _07512_ VGND VGND VPWR VPWR _07522_ sky130_fd_sc_hd__mux2_1
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ clknet_1_0__leaf__08366_ VGND VGND VPWR VPWR _08438_ sky130_fd_sc_hd__buf_1
X_10743_ net2463 _06440_ _06838_ VGND VGND VPWR VPWR _06845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16250_ CPU.registerFile\[10\]\[6\] CPU.registerFile\[11\]\[6\] _03931_ VGND VGND
+ VPWR VPWR _03971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13462_ CPU.Iimm\[2\] _08420_ _08416_ VGND VGND VPWR VPWR _08421_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10674_ net2606 _06465_ _06799_ VGND VGND VPWR VPWR _06807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14240__370 clknet_1_0__leaf__08508_ VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__inv_2
X_17354__14 clknet_1_0__leaf__04985_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__inv_2
X_15201_ _03202_ _03248_ _03252_ _03261_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__a31o_1
X_12413_ _07891_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__clkbuf_1
X_16181_ _03902_ _03903_ _03720_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__mux2_1
X_13685__1060 clknet_1_1__leaf__08453_ VGND VGND VPWR VPWR net1116 sky130_fd_sc_hd__inv_2
XFILLER_0_3_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13393_ _08375_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15132_ _08549_ VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__clkbuf_4
X_12344_ _06609_ net1806 _07848_ VGND VGND VPWR VPWR _07855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15063_ CPU.registerFile\[27\]\[18\] CPU.registerFile\[26\]\[18\] _02768_ VGND VGND
+ VPWR VPWR _03127_ sky130_fd_sc_hd__mux2_1
X_12275_ net1486 _07799_ _07811_ _07809_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__o211a_1
X_13346__842 clknet_1_1__leaf__08367_ VGND VGND VPWR VPWR net898 sky130_fd_sc_hd__inv_2
X_13823__1184 clknet_1_1__leaf__08467_ VGND VGND VPWR VPWR net1240 sky130_fd_sc_hd__inv_2
X_11226_ _07205_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18822_ net611 _02346_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11157_ net1812 _07149_ VGND VGND VPWR VPWR _07161_ sky130_fd_sc_hd__or2_1
X_10108_ _06428_ _06433_ _05800_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__a21oi_1
X_13950__109 clknet_1_0__leaf__08479_ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__inv_2
X_18753_ net542 _02277_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[15\] sky130_fd_sc_hd__dfxtp_1
X_11088_ _07112_ _07116_ VGND VGND VPWR VPWR _07117_ sky130_fd_sc_hd__or2_1
X_15965_ _06085_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__clkbuf_4
X_17704_ CPU.mem_wdata\[4\] per_uart.d_in_uart\[4\] _05218_ VGND VGND VPWR VPWR _05227_
+ sky130_fd_sc_hd__mux2_1
X_14916_ CPU.registerFile\[5\]\[14\] CPU.registerFile\[4\]\[14\] _08864_ VGND VGND
+ VPWR VPWR _02984_ sky130_fd_sc_hd__mux2_1
X_10039_ _06202_ _06365_ _06366_ VGND VGND VPWR VPWR _06367_ sky130_fd_sc_hd__o21ba_1
X_18684_ net473 _02208_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_17635_ net2574 VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__clkbuf_1
X_14847_ CPU.registerFile\[19\]\[13\] CPU.registerFile\[18\]\[13\] _02753_ VGND VGND
+ VPWR VPWR _02916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17566_ net2393 _08360_ _05130_ _07002_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14778_ CPU.registerFile\[30\]\[11\] CPU.registerFile\[31\]\[11\] _08645_ VGND VGND
+ VPWR VPWR _02849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16517_ CPU.registerFile\[2\]\[12\] CPU.registerFile\[3\]\[12\] _04027_ VGND VGND
+ VPWR VPWR _04232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17497_ _08310_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16448_ _06534_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19167_ clknet_leaf_0_clk _02687_ VGND VGND VPWR VPWR per_uart.rx_data\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16379_ CPU.aluIn1\[8\] _04054_ _04097_ _03855_ VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18118_ net1129 _01646_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19098_ net81 _02618_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18049_ net1060 _01577_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_13906__69 clknet_1_0__leaf__08475_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__inv_2
X_14217__350 clknet_1_1__leaf__08505_ VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__inv_2
XFILLER_0_112_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__03638_ clknet_0__03638_ VGND VGND VPWR VPWR clknet_1_1__leaf__03638_
+ sky130_fd_sc_hd__clkbuf_16
X_09822_ _05344_ _06158_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__or2_1
X_09753_ _05343_ _05474_ _05479_ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__a21o_1
X_09684_ CPU.Iimm\[2\] _05758_ _05790_ CPU.cycles\[22\] _06026_ VGND VGND VPWR VPWR
+ _06027_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15948__685 clknet_1_0__leaf__03690_ VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__inv_2
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13650__1029 clknet_1_1__leaf__08449_ VGND VGND VPWR VPWR net1085 sky130_fd_sc_hd__inv_2
XFILLER_0_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_858 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09118_ _05330_ CPU.aluIn1\[14\] VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__or2b_1
XFILLER_0_103_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10390_ _06651_ net2020 _06639_ VGND VGND VPWR VPWR _06652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09049_ _05386_ _05391_ _05396_ _05400_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__or4_1
XFILLER_0_102_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12060_ _07664_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold470 CPU.registerFile\[6\]\[14\] VGND VGND VPWR VPWR net1767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 CPU.registerFile\[28\]\[4\] VGND VGND VPWR VPWR net1778 sky130_fd_sc_hd__dlygate4sd3_1
X_15693__488 clknet_1_1__leaf__03647_ VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__inv_2
X_17335__747 clknet_1_0__leaf__04983_ VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__inv_2
Xhold492 CPU.registerFile\[19\]\[1\] VGND VGND VPWR VPWR net1789 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ net1494 _07007_ _07053_ _07014_ VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__o211a_1
X_12962_ net2181 _07316_ _08181_ VGND VGND VPWR VPWR _08184_ sky130_fd_sc_hd__mux2_1
X_17406__29 clknet_1_1__leaf__05013_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__inv_2
XFILLER_0_99_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1170 CPU.registerFile\[23\]\[6\] VGND VGND VPWR VPWR net2467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1181 CPU.registerFile\[16\]\[28\] VGND VGND VPWR VPWR net2478 sky130_fd_sc_hd__dlygate4sd3_1
X_11913_ _07586_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__clkbuf_1
X_14701_ _08722_ _02767_ _02773_ _08851_ VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__o211a_1
Xhold1192 CPU.registerFile\[1\]\[21\] VGND VGND VPWR VPWR net2489 sky130_fd_sc_hd__dlygate4sd3_1
X_12893_ _08147_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ clknet_1_0__leaf__08340_ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__buf_1
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ net2585 _07356_ _07548_ VGND VGND VPWR VPWR _07550_ sky130_fd_sc_hd__mux2_1
X_14632_ _08785_ _08867_ _08869_ _08870_ VGND VGND VPWR VPWR _08871_ sky130_fd_sc_hd__a211o_1
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _08521_ _08799_ _08801_ _08802_ VGND VGND VPWR VPWR _08803_ sky130_fd_sc_hd__a211o_1
X_17351_ clknet_1_1__leaf__08340_ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__buf_1
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11775_ _07513_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _06171_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__buf_4
XFILLER_0_67_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10726_ net2224 _06245_ _06827_ VGND VGND VPWR VPWR _06836_ sky130_fd_sc_hd__mux2_1
X_14494_ _08567_ _08569_ CPU.registerFile\[9\]\[4\] VGND VGND VPWR VPWR _08736_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17282_ _06085_ _04960_ _04977_ _08596_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__a211o_2
X_19021_ net763 _02541_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16233_ CPU.registerFile\[24\]\[5\] _03915_ _03747_ _03954_ VGND VGND VPWR VPWR _03955_
+ sky130_fd_sc_hd__o211a_1
X_13445_ net2657 _08406_ _08388_ VGND VGND VPWR VPWR _08407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10657_ CPU.registerFile\[1\]\[12\] _06267_ _06788_ VGND VGND VPWR VPWR _06798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16164_ CPU.registerFile\[16\]\[3\] _03848_ _03769_ _03887_ VGND VGND VPWR VPWR _03888_
+ sky130_fd_sc_hd__o211a_1
X_10588_ _06760_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__clkbuf_1
X_12327_ _07843_ _07838_ net1299 mapped_spi_ram.rcv_bitcount\[1\] VGND VGND VPWR VPWR
+ _01683_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15115_ _02964_ _03171_ _03177_ _03092_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16095_ CPU.registerFile\[15\]\[2\] CPU.registerFile\[14\]\[2\] _03705_ VGND VGND
+ VPWR VPWR _03820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15046_ _08418_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__clkbuf_4
X_12258_ net1558 _07799_ _07802_ _07796_ VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11209_ net1630 _07190_ VGND VGND VPWR VPWR _07195_ sky130_fd_sc_hd__nor2_1
X_12189_ net1314 _07749_ _07706_ CPU.mem_wdata\[2\] _07739_ VGND VGND VPWR VPWR _07754_
+ sky130_fd_sc_hd__a221o_1
X_18805_ net594 _02329_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_16997_ CPU.registerFile\[9\]\[24\] _04460_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__or2_1
X_18736_ net525 _02260_ VGND VGND VPWR VPWR mapped_spi_flash.snd_bitcount\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18667_ net456 _02191_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14247__376 clknet_1_0__leaf__08509_ VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__inv_2
X_17618_ _05159_ _05166_ _05167_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__a21oi_1
X_18598_ net419 _02122_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17549_ per_uart.uart0.tx_bitcount\[0\] _05116_ per_uart.uart0.tx_bitcount\[1\] VGND
+ VGND VPWR VPWR _05117_ sky130_fd_sc_hd__and3b_1
XFILLER_0_157_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09805_ _05556_ _06142_ _05731_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__o21a_1
XFILLER_0_157_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09736_ _05881_ _06067_ _06076_ _05744_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__a2bb2o_1
X_09667_ net2072 _06010_ _05742_ VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__mux2_1
X_15729__521 clknet_1_1__leaf__03650_ VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__inv_2
XFILLER_0_69_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15881__625 clknet_1_1__leaf__03683_ VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__inv_2
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ CPU.Iimm\[0\] _05547_ _05922_ CPU.Bimm\[11\] VGND VGND VPWR VPWR _05942_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13822__1183 clknet_1_1__leaf__08467_ VGND VGND VPWR VPWR net1239 sky130_fd_sc_hd__inv_2
XFILLER_0_148_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11560_ net1767 _07347_ _07390_ VGND VGND VPWR VPWR _07398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10511_ _06719_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11491_ net1772 _07356_ _07354_ VGND VGND VPWR VPWR _07357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10442_ _06682_ VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13161_ CPU.cycles\[16\] _08287_ net1538 VGND VGND VPWR VPWR _08290_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10373_ _06640_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__clkbuf_1
X_15701__495 clknet_1_0__leaf__03648_ VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__inv_2
XFILLER_0_20_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12112_ net1326 _07693_ _07701_ _07175_ VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__o211a_1
X_13092_ mapped_spi_flash.rbusy mapped_spi_ram.rbusy VGND VGND VPWR VPWR _08252_ sky130_fd_sc_hd__nor2_1
X_16920_ CPU.registerFile\[10\]\[22\] CPU.registerFile\[11\]\[22\] _04335_ VGND VGND
+ VPWR VPWR _04625_ sky130_fd_sc_hd__mux2_1
X_12043_ _07655_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__clkbuf_1
X_16851_ _04555_ _04556_ _04557_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__mux2_1
X_15802_ _08352_ _03669_ _03661_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__a21oi_1
X_16782_ CPU.registerFile\[20\]\[18\] CPU.registerFile\[21\]\[18\] _04287_ VGND VGND
+ VPWR VPWR _04491_ sky130_fd_sc_hd__mux2_1
X_18521_ net342 _02045_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12945_ net1705 VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18452_ net273 _01980_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_15664_ clknet_1_0__leaf__03643_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__buf_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _06440_ net2213 _08131_ VGND VGND VPWR VPWR _08138_ sky130_fd_sc_hd__mux2_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14615_ CPU.registerFile\[15\]\[7\] CPU.registerFile\[14\]\[7\] _08771_ VGND VGND
+ VPWR VPWR _08854_ sky130_fd_sc_hd__mux2_1
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ net1982 _07339_ _07537_ VGND VGND VPWR VPWR _07541_ sky130_fd_sc_hd__mux2_1
X_18383_ net204 _01911_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14546_ _08585_ _08586_ CPU.registerFile\[1\]\[5\] VGND VGND VPWR VPWR _08787_ sky130_fd_sc_hd__a21o_1
X_11758_ _07504_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10709_ _06815_ VGND VGND VPWR VPWR _06827_ sky130_fd_sc_hd__buf_4
X_17265_ CPU.registerFile\[30\]\[31\] CPU.registerFile\[31\]\[31\] _03739_ VGND VGND
+ VPWR VPWR _04961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11689_ _07467_ VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__clkbuf_1
X_14477_ CPU.registerFile\[21\]\[4\] _08718_ VGND VGND VPWR VPWR _08719_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19004_ clknet_leaf_12_clk _02524_ VGND VGND VPWR VPWR CPU.aluIn1\[21\] sky130_fd_sc_hd__dfxtp_2
X_16216_ CPU.registerFile\[12\]\[5\] _03707_ _03708_ _03937_ VGND VGND VPWR VPWR _03938_
+ sky130_fd_sc_hd__o211a_1
X_13428_ _08393_ VGND VGND VPWR VPWR _08394_ sky130_fd_sc_hd__buf_4
XFILLER_0_125_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17196_ CPU.registerFile\[27\]\[29\] CPU.registerFile\[26\]\[29\] _04646_ VGND VGND
+ VPWR VPWR _04894_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__08461_ _08461_ VGND VGND VPWR VPWR clknet_0__08461_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__08361_ clknet_0__08361_ VGND VGND VPWR VPWR clknet_1_1__leaf__08361_
+ sky130_fd_sc_hd__clkbuf_16
X_16147_ _03716_ _03866_ _03870_ _03732_ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16078_ _03702_ _03800_ _03802_ _03803_ VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__a211o_1
X_15676__472 clknet_1_0__leaf__03646_ VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__inv_2
XFILLER_0_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15029_ _02798_ _03077_ _03084_ _03093_ VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__a31o_1
X_13244__765 clknet_1_0__leaf__08343_ VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__inv_2
X_13896__60 clknet_1_1__leaf__08474_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__inv_2
X_15830__579 clknet_1_1__leaf__03678_ VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__inv_2
Xinput2 resetn VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_2
X_09521_ _05427_ _05863_ _05865_ _05517_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__o211a_1
X_18719_ net508 _02243_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09452_ _05410_ _05522_ _05798_ _05800_ VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__o22ai_1
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14180__316 clknet_1_1__leaf__08502_ VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__inv_2
XFILLER_0_137_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09383_ CPU.Bimm\[1\] VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__buf_4
XFILLER_0_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14000__153 clknet_1_1__leaf__08485_ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__inv_2
XFILLER_0_113_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14074__221 clknet_1_1__leaf__08491_ VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__inv_2
XFILLER_0_100_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__08450_ clknet_0__08450_ VGND VGND VPWR VPWR clknet_1_0__leaf__08450_
+ sky130_fd_sc_hd__clkbuf_16
X_09719_ _06058_ _06059_ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__and2_1
X_10991_ _05615_ _07028_ VGND VGND VPWR VPWR _07036_ sky130_fd_sc_hd__xnor2_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _08059_ VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__clkbuf_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17396__20 clknet_1_1__leaf__04985_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__inv_2
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12661_ _06653_ net1867 _08015_ VGND VGND VPWR VPWR _08023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ net1833 _07330_ _07416_ VGND VGND VPWR VPWR _07426_ sky130_fd_sc_hd__mux2_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _08521_ _08641_ _08643_ _08533_ VGND VGND VPWR VPWR _08644_ sky130_fd_sc_hd__a211o_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _07986_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__clkbuf_1
X_15380_ _03434_ _03435_ _03255_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11543_ net1908 _07330_ _07379_ VGND VGND VPWR VPWR _07389_ sky130_fd_sc_hd__mux2_1
X_14331_ CPU.registerFile\[5\]\[0\] CPU.registerFile\[4\]\[0\] _08576_ VGND VGND VPWR
+ VPWR _08577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13310__811 clknet_1_1__leaf__08362_ VGND VGND VPWR VPWR net867 sky130_fd_sc_hd__inv_2
X_17050_ CPU.registerFile\[28\]\[25\] CPU.registerFile\[29\]\[25\] _04526_ VGND VGND
+ VPWR VPWR _04752_ sky130_fd_sc_hd__mux2_1
X_11474_ _06199_ VGND VGND VPWR VPWR _07345_ sky130_fd_sc_hd__buf_4
XFILLER_0_151_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16001_ _03726_ _03727_ CPU.registerFile\[1\]\[0\] VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__a21o_1
X_13213_ _05522_ _08326_ _06545_ VGND VGND VPWR VPWR _08327_ sky130_fd_sc_hd__mux2_1
X_10425_ _06673_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13144_ _08279_ _08280_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__nor2_1
X_10356_ _06628_ net1944 _06618_ VGND VGND VPWR VPWR _06629_ sky130_fd_sc_hd__mux2_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ net1386 VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__clkbuf_1
X_17952_ net963 _01480_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_10287_ net2133 _06361_ _06580_ VGND VGND VPWR VPWR _06584_ sky130_fd_sc_hd__mux2_1
X_12026_ CPU.registerFile\[24\]\[21\] _07332_ _07646_ VGND VGND VPWR VPWR _07647_
+ sky130_fd_sc_hd__mux2_1
X_16903_ CPU.registerFile\[27\]\[21\] CPU.registerFile\[26\]\[21\] _04242_ VGND VGND
+ VPWR VPWR _04609_ sky130_fd_sc_hd__mux2_1
X_17883_ clknet_leaf_20_clk _00033_ VGND VGND VPWR VPWR CPU.cycles\[26\] sky130_fd_sc_hd__dfxtp_1
X_16834_ _06474_ VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__clkbuf_4
X_16765_ CPU.registerFile\[0\]\[18\] _04233_ _04472_ _04473_ VGND VGND VPWR VPWR _04474_
+ sky130_fd_sc_hd__o211a_1
X_13536__926 clknet_1_0__leaf__08438_ VGND VGND VPWR VPWR net982 sky130_fd_sc_hd__inv_2
X_18504_ net325 _02028_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_12928_ _08165_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__clkbuf_1
X_16696_ CPU.registerFile\[19\]\[16\] CPU.registerFile\[18\]\[16\] _04327_ VGND VGND
+ VPWR VPWR _04407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18435_ net256 _01963_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18584__41 VGND VGND VPWR VPWR _18584__41/HI net41 sky130_fd_sc_hd__conb_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _06245_ net2004 _08120_ VGND VGND VPWR VPWR _08129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18366_ net187 _01894_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15578_ CPU.registerFile\[5\]\[31\] CPU.registerFile\[4\]\[31\] _08558_ VGND VGND
+ VPWR VPWR _03629_ sky130_fd_sc_hd__mux2_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14529_ _08515_ _08755_ _08760_ _08769_ VGND VGND VPWR VPWR _08770_ sky130_fd_sc_hd__a31o_1
X_18297_ net118 _01825_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17248_ CPU.registerFile\[10\]\[31\] CPU.registerFile\[11\]\[31\] _06173_ VGND VGND
+ VPWR VPWR _04944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17179_ _03703_ _04874_ _04876_ _06142_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__08444_ _08444_ VGND VGND VPWR VPWR clknet_0__08444_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__08344_ clknet_0__08344_ VGND VGND VPWR VPWR clknet_1_1__leaf__08344_
+ sky130_fd_sc_hd__clkbuf_16
X_08952_ _05294_ _05298_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__nor2_1
X_13821__1182 clknet_1_1__leaf__08467_ VGND VGND VPWR VPWR net1238 sky130_fd_sc_hd__inv_2
X_08883_ _05236_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09504_ _05403_ _05843_ _05844_ _05849_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__a211o_2
X_09435_ _05745_ _05781_ _05782_ _05784_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__a211o_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09366_ _05708_ _05704_ _05659_ _05716_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__and4b_1
XFILLER_0_90_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09297_ _05645_ _05648_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__xnor2_1
XANTENNA_40 _08419_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 clknet_1_0__leaf__08473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 net1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _08520_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 _07464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10210_ _06531_ VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11190_ _07129_ _07180_ _07130_ VGND VGND VPWR VPWR _07181_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10141_ net2322 _06465_ _06293_ VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10072_ _05966_ _05948_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__and2b_1
X_15887__631 clknet_1_0__leaf__03683_ VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__inv_2
X_14880_ _02831_ _02832_ CPU.registerFile\[1\]\[13\] VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__a21o_1
Xclkbuf_1_0__f__08502_ clknet_0__08502_ VGND VGND VPWR VPWR clknet_1_0__leaf__08502_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13831_ clknet_1_0__leaf__08462_ VGND VGND VPWR VPWR _08468_ sky130_fd_sc_hd__buf_1
XFILLER_0_97_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16550_ CPU.registerFile\[15\]\[13\] CPU.registerFile\[14\]\[13\] _04146_ VGND VGND
+ VPWR VPWR _04264_ sky130_fd_sc_hd__mux2_1
X_10974_ mapped_spi_flash.cmd_addr\[15\] _05667_ _07009_ VGND VGND VPWR VPWR _07021_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__08364_ clknet_0__08364_ VGND VGND VPWR VPWR clknet_1_0__leaf__08364_
+ sky130_fd_sc_hd__clkbuf_16
X_15501_ _08543_ _03551_ _03553_ _03307_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__a211o_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12713_ _08050_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13985__141 clknet_1_1__leaf__08482_ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__inv_2
X_16481_ CPU.registerFile\[0\]\[11\] _03828_ _04068_ _04196_ VGND VGND VPWR VPWR _04197_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18220_ net1231 _01748_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[21\] sky130_fd_sc_hd__dfxtp_1
X_15432_ CPU.registerFile\[5\]\[27\] CPU.registerFile\[4\]\[27\] _08558_ VGND VGND
+ VPWR VPWR _03487_ sky130_fd_sc_hd__mux2_1
X_12644_ _06636_ net1971 _08004_ VGND VGND VPWR VPWR _08014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18151_ net1162 _01679_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_12575_ _07977_ VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__clkbuf_1
X_15363_ _03235_ _03236_ CPU.registerFile\[1\]\[25\] VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__a21o_1
X_17102_ _04545_ _04785_ _04802_ _04500_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__a211o_2
X_14314_ _06061_ VGND VGND VPWR VPWR _08560_ sky130_fd_sc_hd__buf_4
X_11526_ _07380_ VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__clkbuf_1
X_18082_ net1093 _01610_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_15294_ _03344_ _03352_ _03241_ VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__o21a_2
XFILLER_0_151_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17033_ CPU.registerFile\[9\]\[25\] _04460_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__or2_1
X_11457_ net1721 _07332_ _07333_ VGND VGND VPWR VPWR _07334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10408_ _06594_ _06663_ VGND VGND VPWR VPWR _06664_ sky130_fd_sc_hd__nand2_4
X_11388_ _07291_ VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__clkbuf_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _06053_ VGND VGND VPWR VPWR _06617_ sky130_fd_sc_hd__buf_4
X_13127_ _08269_ net1570 VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__nor2_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ clknet_leaf_18_clk _02504_ VGND VGND VPWR VPWR CPU.aluIn1\[1\] sky130_fd_sc_hd__dfxtp_4
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _08234_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__clkbuf_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17935_ net946 _01463_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_12009_ net2423 _07316_ _07635_ VGND VGND VPWR VPWR _07638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17866_ clknet_leaf_25_clk _00046_ VGND VGND VPWR VPWR CPU.cycles\[9\] sky130_fd_sc_hd__dfxtp_1
X_16817_ CPU.registerFile\[30\]\[19\] CPU.registerFile\[31\]\[19\] _04201_ VGND VGND
+ VPWR VPWR _04525_ sky130_fd_sc_hd__mux2_1
X_17797_ net877 _01359_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16748_ CPU.aluIn1\[17\] _04054_ _04457_ _04259_ VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13317__817 clknet_1_1__leaf__08363_ VGND VGND VPWR VPWR net873 sky130_fd_sc_hd__inv_2
X_16679_ _05690_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09220_ CPU.Iimm\[3\] CPU.Bimm\[3\] CPU.instr\[5\] VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18418_ net239 _01946_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09151_ _05400_ _05501_ _05502_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__a21o_1
X_18349_ net170 _01877_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09082_ _05277_ _05244_ _05278_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold800 CPU.registerFile\[11\]\[30\] VGND VGND VPWR VPWR net2097 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold811 CPU.registerFile\[30\]\[24\] VGND VGND VPWR VPWR net2108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold822 CPU.registerFile\[14\]\[28\] VGND VGND VPWR VPWR net2119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold833 CPU.registerFile\[30\]\[19\] VGND VGND VPWR VPWR net2130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 CPU.registerFile\[23\]\[19\] VGND VGND VPWR VPWR net2141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold855 CPU.registerFile\[23\]\[16\] VGND VGND VPWR VPWR net2152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 CPU.registerFile\[18\]\[31\] VGND VGND VPWR VPWR net2163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold877 CPU.registerFile\[21\]\[17\] VGND VGND VPWR VPWR net2174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 CPU.registerFile\[11\]\[16\] VGND VGND VPWR VPWR net2185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 CPU.registerFile\[26\]\[25\] VGND VGND VPWR VPWR net2196 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ _05745_ _06304_ _06310_ _06314_ VGND VGND VPWR VPWR _06315_ sky130_fd_sc_hd__a211o_2
XFILLER_0_0_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08935_ CPU.mem_wdata\[4\] CPU.Iimm\[4\] _05244_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__mux2_2
XFILLER_0_99_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14112__254 clknet_1_0__leaf__08496_ VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__03691_ clknet_0__03691_ VGND VGND VPWR VPWR clknet_1_0__leaf__03691_
+ sky130_fd_sc_hd__clkbuf_16
X_09418_ _05768_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10690_ _06817_ VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09349_ _05700_ _05583_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12360_ _07863_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13841__1201 clknet_1_1__leaf__08468_ VGND VGND VPWR VPWR net1257 sky130_fd_sc_hd__inv_2
X_11311_ net1868 _06083_ _07249_ VGND VGND VPWR VPWR _07251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12291_ net1473 _07812_ _07820_ _07809_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11242_ _06620_ net1928 _07212_ VGND VGND VPWR VPWR _07214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11173_ net1401 _07134_ VGND VGND VPWR VPWR _07170_ sky130_fd_sc_hd__or2_1
X_10124_ _05514_ _05290_ _06202_ _06446_ _06448_ VGND VGND VPWR VPWR _06449_ sky130_fd_sc_hd__a311o_2
X_15981_ _06149_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__clkbuf_4
X_10055_ _05744_ _06379_ _06381_ _06382_ VGND VGND VPWR VPWR _06383_ sky130_fd_sc_hd__a22o_1
X_14932_ CPU.registerFile\[22\]\[15\] CPU.registerFile\[23\]\[15\] _02998_ VGND VGND
+ VPWR VPWR _02999_ sky130_fd_sc_hd__mux2_1
X_17651_ net1766 _05185_ _05188_ _07002_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__o211a_1
X_14863_ _08722_ _02926_ _02931_ _08851_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16602_ CPU.registerFile\[30\]\[14\] CPU.registerFile\[31\]\[14\] _04201_ VGND VGND
+ VPWR VPWR _04315_ sky130_fd_sc_hd__mux2_1
X_17582_ _05143_ VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__clkbuf_1
X_14794_ CPU.registerFile\[8\]\[11\] _08776_ _02863_ _02864_ VGND VGND VPWR VPWR _02865_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16533_ CPU.registerFile\[22\]\[12\] CPU.registerFile\[23\]\[12\] _03958_ VGND VGND
+ VPWR VPWR _04248_ sky130_fd_sc_hd__mux2_1
X_10957_ _06976_ VGND VGND VPWR VPWR _07009_ sky130_fd_sc_hd__buf_4
XFILLER_0_85_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16464_ _04170_ _04173_ _04179_ _04180_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__o211a_1
X_13676_ clknet_1_0__leaf__08451_ VGND VGND VPWR VPWR _08453_ sky130_fd_sc_hd__buf_1
X_10888_ _05284_ _06955_ _06880_ VGND VGND VPWR VPWR _06956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18203_ net1214 _01731_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[4\] sky130_fd_sc_hd__dfxtp_1
X_15415_ CPU.registerFile\[28\]\[27\] CPU.registerFile\[29\]\[27\] _03212_ VGND VGND
+ VPWR VPWR _03470_ sky130_fd_sc_hd__mux2_1
X_12627_ _08005_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__clkbuf_1
X_19183_ clknet_leaf_0_clk _02701_ VGND VGND VPWR VPWR per_uart.uart_ctrl\[2\] sky130_fd_sc_hd__dfxtp_1
X_16395_ _04111_ _04112_ _03720_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18134_ net1145 _01662_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15346_ _03049_ _03050_ CPU.registerFile\[25\]\[25\] VGND VGND VPWR VPWR _03403_
+ sky130_fd_sc_hd__a21o_1
X_12558_ net2058 _07332_ _07968_ VGND VGND VPWR VPWR _07969_ sky130_fd_sc_hd__mux2_1
X_15640__441 clknet_1_1__leaf__03641_ VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__inv_2
XFILLER_0_53_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18065_ net1076 _01593_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11509_ net1856 _07368_ _07354_ VGND VGND VPWR VPWR _07369_ sky130_fd_sc_hd__mux2_1
X_15277_ _03202_ _03323_ _03327_ _03335_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__a31o_1
X_12489_ net2053 _07332_ _07931_ VGND VGND VPWR VPWR _07932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold107 mapped_spi_ram.cmd_addr\[21\] VGND VGND VPWR VPWR net1404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold118 _08235_ VGND VGND VPWR VPWR net1415 sky130_fd_sc_hd__dlygate4sd3_1
X_17016_ CPU.registerFile\[27\]\[24\] CPU.registerFile\[26\]\[24\] _04646_ VGND VGND
+ VPWR VPWR _04719_ sky130_fd_sc_hd__mux2_1
Xhold129 mapped_spi_ram.cmd_addr\[19\] VGND VGND VPWR VPWR net1426 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__03654_ clknet_0__03654_ VGND VGND VPWR VPWR clknet_1_1__leaf__03654_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__03685_ _03685_ VGND VGND VPWR VPWR clknet_0__03685_ sky130_fd_sc_hd__clkbuf_16
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18967_ net741 _02487_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17918_ clknet_leaf_26_clk _01446_ VGND VGND VPWR VPWR CPU.Bimm\[5\] sky130_fd_sc_hd__dfxtp_4
X_18898_ net672 _02418_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_13763__1131 clknet_1_1__leaf__08460_ VGND VGND VPWR VPWR net1187 sky130_fd_sc_hd__inv_2
X_17849_ net929 _01411_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09203_ CPU.Jimm\[13\] VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__inv_4
XFILLER_0_17_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09134_ _05356_ _05474_ _05478_ _05485_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__a31o_1
XFILLER_0_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09065_ CPU.aluIn1\[31\] _05416_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__or2_2
XFILLER_0_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold630 CPU.registerFile\[18\]\[19\] VGND VGND VPWR VPWR net1927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold641 CPU.registerFile\[17\]\[24\] VGND VGND VPWR VPWR net1938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 CPU.registerFile\[15\]\[24\] VGND VGND VPWR VPWR net1949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 _05175_ VGND VGND VPWR VPWR net1960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 CPU.registerFile\[27\]\[12\] VGND VGND VPWR VPWR net1971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 CPU.registerFile\[9\]\[18\] VGND VGND VPWR VPWR net1982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 CPU.registerFile\[11\]\[2\] VGND VGND VPWR VPWR net1993 sky130_fd_sc_hd__dlygate4sd3_1
X_13932__92 clknet_1_1__leaf__08478_ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__inv_2
X_09967_ _05310_ _06297_ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__nor2_1
X_08918_ CPU.mem_wdata\[2\] CPU.Iimm\[2\] _05244_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__mux2_2
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _05323_ _05522_ _05749_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__o21ai_1
Xhold1330 CPU.registerFile\[12\]\[14\] VGND VGND VPWR VPWR net2627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1341 CPU.registerFile\[25\]\[19\] VGND VGND VPWR VPWR net2638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1352 mapped_spi_flash.div_counter\[0\] VGND VGND VPWR VPWR net2649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1363 CPU.aluReg\[22\] VGND VGND VPWR VPWR net2660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1374 CPU.aluReg\[2\] VGND VGND VPWR VPWR net2671 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ net2443 _07372_ _07548_ VGND VGND VPWR VPWR _07558_ sky130_fd_sc_hd__mux2_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ CPU.aluReg\[24\] CPU.aluReg\[22\] _06872_ VGND VGND VPWR VPWR _06897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11791_ _07521_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__clkbuf_1
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15925__664 clknet_1_1__leaf__03688_ VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__inv_2
XFILLER_0_95_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10742_ _06844_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10673_ _06806_ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__clkbuf_1
X_13461_ _08419_ VGND VGND VPWR VPWR _08420_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15200_ _02964_ _03256_ _03260_ _03092_ VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__o211a_1
X_12412_ net1886 _07324_ _07884_ VGND VGND VPWR VPWR _07891_ sky130_fd_sc_hd__mux2_1
X_16180_ CPU.registerFile\[5\]\[4\] CPU.registerFile\[4\]\[4\] _03704_ VGND VGND VPWR
+ VPWR _03903_ sky130_fd_sc_hd__mux2_1
X_13392_ _06390_ _08372_ _08374_ VGND VGND VPWR VPWR _08375_ sky130_fd_sc_hd__and3_1
X_13489__883 clknet_1_1__leaf__08434_ VGND VGND VPWR VPWR net939 sky130_fd_sc_hd__inv_2
XFILLER_0_51_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15131_ _02831_ _02832_ CPU.registerFile\[1\]\[19\] VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__a21o_1
X_12343_ _07854_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12274_ mapped_spi_ram.rcv_data\[12\] _07800_ VGND VGND VPWR VPWR _07811_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15062_ _03124_ _03125_ _02851_ VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__mux2_1
X_11225_ _06603_ net1952 _07201_ VGND VGND VPWR VPWR _07205_ sky130_fd_sc_hd__mux2_1
X_11156_ _07132_ VGND VGND VPWR VPWR _07160_ sky130_fd_sc_hd__buf_2
X_18821_ net610 _02345_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10107_ _05794_ _06432_ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__or2_1
X_18752_ net541 _02276_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[14\] sky130_fd_sc_hd__dfxtp_1
X_11087_ mapped_spi_flash.snd_bitcount\[1\] mapped_spi_flash.snd_bitcount\[0\] _06978_
+ mapped_spi_flash.snd_bitcount\[4\] VGND VGND VPWR VPWR _07116_ sky130_fd_sc_hd__o31a_1
X_15670__467 clknet_1_1__leaf__03645_ VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__inv_2
X_17312__726 clknet_1_0__leaf__04981_ VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__inv_2
X_17703_ _05226_ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__clkbuf_1
X_14915_ CPU.registerFile\[6\]\[14\] CPU.registerFile\[7\]\[14\] _02982_ VGND VGND
+ VPWR VPWR _02983_ sky130_fd_sc_hd__mux2_1
X_10038_ _05520_ _05697_ _05726_ VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__and3_1
X_18683_ net472 _02207_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_17634_ net2573 per_uart.uart0.rxd_reg\[7\] _05170_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__mux2_1
X_14846_ net1665 _02797_ _02915_ _08751_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17565_ _08360_ _05129_ net2393 VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__o21ai_1
X_14777_ _08837_ _02845_ _02847_ _08802_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__a211o_1
XFILLER_0_58_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11989_ _07626_ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16516_ _04229_ _04230_ _04153_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17496_ _05069_ net2630 _05072_ _05074_ _05053_ VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16447_ CPU.registerFile\[27\]\[10\] CPU.registerFile\[26\]\[10\] _03837_ VGND VGND
+ VPWR VPWR _04164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19166_ clknet_leaf_0_clk _02686_ VGND VGND VPWR VPWR per_uart.rx_data\[5\] sky130_fd_sc_hd__dfxtp_1
X_16378_ _03692_ _04074_ _04095_ _04096_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__a211o_1
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18117_ net1128 _01645_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15329_ _03230_ _03382_ _03386_ _03151_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19097_ net80 _02617_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18048_ net1059 _01576_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09821_ _05343_ _05336_ _05338_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09752_ _05351_ _06091_ VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__xnor2_2
X_17287__703 clknet_1_1__leaf__04979_ VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__inv_2
X_09683_ _05881_ _06016_ _06025_ _05744_ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__a2bb2o_1
X_13840__1200 clknet_1_1__leaf__08468_ VGND VGND VPWR VPWR net1256 sky130_fd_sc_hd__inv_2
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15647__447 clknet_1_1__leaf__03642_ VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__inv_2
XFILLER_0_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14224__355 clknet_1_1__leaf__08507_ VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__inv_2
XFILLER_0_91_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09117_ CPU.aluIn1\[12\] _05317_ _05457_ _05468_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09048_ _05398_ _05399_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__or2_2
XFILLER_0_103_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold460 CPU.registerFile\[30\]\[25\] VGND VGND VPWR VPWR net1757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 CPU.registerFile\[28\]\[20\] VGND VGND VPWR VPWR net1768 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ _07048_ _07052_ VGND VGND VPWR VPWR _07053_ sky130_fd_sc_hd__or2_1
Xhold482 CPU.registerFile\[19\]\[2\] VGND VGND VPWR VPWR net1779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold493 CPU.registerFile\[13\]\[13\] VGND VGND VPWR VPWR net1790 sky130_fd_sc_hd__dlygate4sd3_1
X_14118__260 clknet_1_1__leaf__08496_ VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__inv_2
X_12961_ _08183_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__clkbuf_1
Xhold1160 CPU.registerFile\[23\]\[7\] VGND VGND VPWR VPWR net2457 sky130_fd_sc_hd__dlygate4sd3_1
X_14700_ _08764_ _02769_ _02772_ _08552_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__a211o_1
Xhold1171 CPU.registerFile\[29\]\[9\] VGND VGND VPWR VPWR net2468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 CPU.registerFile\[6\]\[27\] VGND VGND VPWR VPWR net2479 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11912_ _06641_ net2278 _07584_ VGND VGND VPWR VPWR _07586_ sky130_fd_sc_hd__mux2_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1193 CPU.registerFile\[13\]\[2\] VGND VGND VPWR VPWR net2490 sky130_fd_sc_hd__dlygate4sd3_1
X_12892_ _05767_ net2377 _08145_ VGND VGND VPWR VPWR _08147_ sky130_fd_sc_hd__mux2_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _08418_ VGND VGND VPWR VPWR _08870_ sky130_fd_sc_hd__clkbuf_4
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _07549_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__clkbuf_1
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _08532_ VGND VGND VPWR VPWR _08802_ sky130_fd_sc_hd__clkbuf_4
X_15706__500 clknet_1_1__leaf__03648_ VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__inv_2
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _06638_ net2491 _07512_ VGND VGND VPWR VPWR _07513_ sky130_fd_sc_hd__mux2_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _04015_ _04016_ _04020_ _03979_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__a211o_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17281_ _04968_ _04976_ _06474_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__o21a_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ _06835_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__clkbuf_1
X_14493_ CPU.registerFile\[10\]\[4\] CPU.registerFile\[11\]\[4\] _08564_ VGND VGND
+ VPWR VPWR _08735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19020_ net762 _02540_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16232_ _03749_ _03751_ CPU.registerFile\[25\]\[5\] VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__a21o_1
X_13444_ _06474_ VGND VGND VPWR VPWR _08406_ sky130_fd_sc_hd__clkbuf_4
X_10656_ _06797_ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16163_ _03770_ _03771_ CPU.registerFile\[17\]\[3\] VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__a21o_1
XFILLER_0_141_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13762__1130 clknet_1_1__leaf__08460_ VGND VGND VPWR VPWR net1186 sky130_fd_sc_hd__inv_2
X_10587_ net2180 _06267_ _06750_ VGND VGND VPWR VPWR _06760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15114_ _03006_ _03173_ _03176_ _02814_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__a211o_1
X_12326_ mapped_spi_ram.rcv_bitcount\[0\] net1298 _07835_ VGND VGND VPWR VPWR _07845_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16094_ _08398_ _03816_ _03818_ _08401_ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__a211o_1
XFILLER_0_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15045_ CPU.registerFile\[0\]\[17\] _02948_ _03109_ _02791_ VGND VGND VPWR VPWR _03110_
+ sky130_fd_sc_hd__o211a_1
X_12257_ net1524 _07800_ VGND VGND VPWR VPWR _07802_ sky130_fd_sc_hd__or2_1
X_11208_ _07126_ _07190_ net1434 VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__o21ai_1
X_12188_ net1343 _07738_ _07753_ _07737_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__o211a_1
X_18804_ net593 _02328_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11139_ net1370 _07147_ _07150_ _07151_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__o211a_1
X_13911__73 clknet_1_1__leaf__08476_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__inv_2
X_16996_ CPU.registerFile\[10\]\[24\] CPU.registerFile\[11\]\[24\] _04335_ VGND VGND
+ VPWR VPWR _04699_ sky130_fd_sc_hd__mux2_1
X_18735_ net524 net1457 VGND VGND VPWR VPWR mapped_spi_flash.snd_bitcount\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18666_ net455 _02190_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14829_ _02897_ _02898_ _08695_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__mux2_1
X_17617_ _06973_ _05129_ net1449 VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__a21oi_1
X_18597_ net418 _02121_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17548_ per_uart.uart0.tx_bitcount\[2\] per_uart.uart0.tx_bitcount\[3\] VGND VGND
+ VPWR VPWR _05116_ sky130_fd_sc_hd__and2b_1
XFILLER_0_157_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17479_ _08379_ _05017_ _06282_ VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_144_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19149_ clknet_leaf_6_clk _02669_ VGND VGND VPWR VPWR per_uart.uart0.tx_bitcount\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_125_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09804_ _06141_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__clkbuf_8
X_09735_ _06072_ _06074_ _06075_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__or3_1
X_09666_ _06009_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__buf_4
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ CPU.PC\[12\] _05923_ _05940_ VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__or3_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411__33 clknet_1_1__leaf__05014_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__inv_2
XFILLER_0_65_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10510_ net2060 _06169_ _06713_ VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11490_ _06315_ VGND VGND VPWR VPWR _07356_ sky130_fd_sc_hd__buf_4
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10441_ _06628_ net2422 _06676_ VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10372_ _06638_ net2171 _06639_ VGND VGND VPWR VPWR _06640_ sky130_fd_sc_hd__mux2_1
X_13160_ CPU.cycles\[16\] CPU.cycles\[17\] _08287_ VGND VGND VPWR VPWR _08289_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12111_ net1325 _07694_ _07696_ VGND VGND VPWR VPWR _07701_ sky130_fd_sc_hd__a21o_1
X_13091_ net1359 VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12042_ CPU.registerFile\[24\]\[13\] _07349_ _07646_ VGND VGND VPWR VPWR _07655_
+ sky130_fd_sc_hd__mux2_1
Xhold290 per_uart.uart0.enable16_counter\[10\] VGND VGND VPWR VPWR net1587 sky130_fd_sc_hd__dlygate4sd3_1
X_14051__200 clknet_1_0__leaf__08489_ VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__inv_2
X_16850_ _06534_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__buf_4
X_15801_ net1596 _08351_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__nand2_1
X_16781_ CPU.registerFile\[22\]\[18\] CPU.registerFile\[23\]\[18\] _04362_ VGND VGND
+ VPWR VPWR _04490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18520_ net341 _02044_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12944_ _06440_ net1704 _08167_ VGND VGND VPWR VPWR _08174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18451_ net272 _01979_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _08137_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14614_ _08515_ _08836_ _08843_ _08852_ VGND VGND VPWR VPWR _08853_ sky130_fd_sc_hd__a31o_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _07540_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__clkbuf_1
X_18382_ net203 _01910_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15782__568 clknet_1_1__leaf__03656_ VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__inv_2
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ CPU.registerFile\[2\]\[5\] CPU.registerFile\[3\]\[5\] _08629_ VGND VGND VPWR
+ VPWR _08786_ sky130_fd_sc_hd__mux2_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _06622_ net2109 _07501_ VGND VGND VPWR VPWR _07504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17264_ _03755_ _04947_ _04951_ _04959_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__a31o_1
X_10708_ _06826_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14476_ _06062_ VGND VGND VPWR VPWR _08718_ sky130_fd_sc_hd__buf_2
X_11688_ net2604 _07337_ _07464_ VGND VGND VPWR VPWR _07467_ sky130_fd_sc_hd__mux2_1
X_19003_ clknet_leaf_12_clk _02523_ VGND VGND VPWR VPWR CPU.aluIn1\[20\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_153_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16215_ CPU.registerFile\[13\]\[5\] _03709_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__or2_1
X_13427_ _06172_ VGND VGND VPWR VPWR _08393_ sky130_fd_sc_hd__buf_4
X_10639_ net2489 _06054_ _06788_ VGND VGND VPWR VPWR _06789_ sky130_fd_sc_hd__mux2_1
X_17195_ _04891_ _04892_ _06535_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__08460_ _08460_ VGND VGND VPWR VPWR clknet_0__08460_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16146_ _03722_ _03867_ _03869_ _03730_ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__a211o_1
XFILLER_0_140_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12309_ _07782_ _07831_ VGND VGND VPWR VPWR _07832_ sky130_fd_sc_hd__nand2_1
X_16077_ _06141_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__clkbuf_4
X_13289_ clknet_1_0__leaf__08341_ VGND VGND VPWR VPWR _08361_ sky130_fd_sc_hd__buf_1
X_15028_ _02964_ _03087_ _03091_ _03092_ VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput3 spi_miso VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
X_16979_ _04681_ _04682_ _06535_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09520_ _05808_ _05864_ _05425_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__o21ai_1
X_18718_ net507 _02242_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[18\] sky130_fd_sc_hd__dfxtp_1
X_09451_ _05799_ _05520_ VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__nand2_4
X_18649_ clknet_leaf_11_clk _02173_ VGND VGND VPWR VPWR CPU.rs2\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13513__905 clknet_1_0__leaf__08436_ VGND VGND VPWR VPWR net961 sky130_fd_sc_hd__inv_2
X_09382_ _05733_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15759__548 clknet_1_1__leaf__03653_ VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__inv_2
XFILLER_0_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08489_ clknet_0__08489_ VGND VGND VPWR VPWR clknet_1_1__leaf__08489_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09718_ mapped_spi_ram.rcv_data\[12\] _05683_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__nand2_8
X_10990_ net1493 _07007_ _07035_ _07014_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09649_ _05937_ _05986_ _05990_ _05992_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__a31o_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _08022_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__clkbuf_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11611_ _07425_ VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__clkbuf_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12591_ net2465 _07366_ _07979_ VGND VGND VPWR VPWR _07986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14330_ _06062_ VGND VGND VPWR VPWR _08576_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_135_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11542_ _07388_ VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11473_ _07344_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__clkbuf_1
X_16000_ _05690_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__buf_4
X_13212_ _05514_ _05534_ VGND VGND VPWR VPWR _08326_ sky130_fd_sc_hd__nand2_1
X_10424_ _06611_ net2195 _06665_ VGND VGND VPWR VPWR _06673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13143_ net1559 _08277_ VGND VGND VPWR VPWR _08280_ sky130_fd_sc_hd__nor2_1
X_10355_ _06168_ VGND VGND VPWR VPWR _06628_ sky130_fd_sc_hd__buf_4
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _06583_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__clkbuf_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ CPU.registerFile\[4\]\[8\] net1385 _08239_ VGND VGND VPWR VPWR _08243_ sky130_fd_sc_hd__mux2_1
X_17951_ net962 _01479_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12025_ _07634_ VGND VGND VPWR VPWR _07646_ sky130_fd_sc_hd__buf_4
X_16902_ _04606_ _04607_ _04279_ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__mux2_1
X_17882_ clknet_leaf_20_clk _00032_ VGND VGND VPWR VPWR CPU.cycles\[25\] sky130_fd_sc_hd__dfxtp_1
X_16833_ _04170_ _04536_ _04540_ _04180_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__o211a_1
X_16764_ _04389_ _04390_ CPU.registerFile\[1\]\[18\] VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__a21o_1
X_15864__610 clknet_1_1__leaf__03681_ VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__inv_2
X_18503_ net324 _02027_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12927_ _06245_ net2186 _08156_ VGND VGND VPWR VPWR _08165_ sky130_fd_sc_hd__mux2_1
X_16695_ _04404_ _04405_ _04365_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18434_ net255 _01962_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12858_ _08128_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__clkbuf_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18365_ net186 _01893_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_11809_ _07531_ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__clkbuf_1
X_15577_ CPU.registerFile\[6\]\[31\] CPU.registerFile\[7\]\[31\] _08536_ VGND VGND
+ VPWR VPWR _03628_ sky130_fd_sc_hd__mux2_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12789_ _06645_ net2164 _08087_ VGND VGND VPWR VPWR _08091_ sky130_fd_sc_hd__mux2_1
X_13962__120 clknet_1_1__leaf__08480_ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__inv_2
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14528_ _08722_ _08763_ _08768_ _08554_ VGND VGND VPWR VPWR _08769_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18296_ net117 _01824_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17247_ net2420 _08513_ _04943_ _04663_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__o211a_1
X_14459_ CPU.registerFile\[6\]\[3\] CPU.registerFile\[7\]\[3\] _08522_ VGND VGND VPWR
+ VPWR _08702_ sky130_fd_sc_hd__mux2_1
X_14058__206 clknet_1_0__leaf__08490_ VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__inv_2
X_17178_ CPU.registerFile\[8\]\[29\] _03707_ _03708_ _04875_ VGND VGND VPWR VPWR _04876_
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_0__08443_ _08443_ VGND VGND VPWR VPWR clknet_0__08443_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16129_ _03692_ _03833_ _03853_ _03601_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_1__f__08343_ clknet_0__08343_ VGND VGND VPWR VPWR clknet_1_1__leaf__08343_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08951_ _05284_ _05285_ _05302_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__o21ai_1
X_08882_ _05235_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__inv_6
XFILLER_0_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09503_ _05427_ _05845_ _05848_ _05517_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09434_ _05556_ _05783_ _05764_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__o21a_1
X_15765__552 clknet_1_0__leaf__03655_ VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__inv_2
XFILLER_0_149_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09365_ _05704_ _05708_ _05716_ _05659_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__and4b_2
XANTENNA_30 _06062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09296_ _05646_ _05647_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__nor2_1
XANTENNA_41 _08419_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_52 clknet_1_1__leaf__08473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 CPU.mem_wdata\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_74 _08520_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10140_ _06464_ VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__buf_4
X_13779__1144 clknet_1_1__leaf__08463_ VGND VGND VPWR VPWR net1200 sky130_fd_sc_hd__inv_2
XFILLER_0_11_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10071_ _06389_ _06392_ _06397_ _05556_ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__a22o_1
X_13340__838 clknet_1_1__leaf__08365_ VGND VGND VPWR VPWR net894 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__08501_ clknet_0__08501_ VGND VGND VPWR VPWR clknet_1_0__leaf__08501_
+ sky130_fd_sc_hd__clkbuf_16
X_10973_ net1552 _07007_ _07020_ _07014_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_0__f__08363_ clknet_0__08363_ VGND VGND VPWR VPWR clknet_1_0__leaf__08363_
+ sky130_fd_sc_hd__clkbuf_16
X_15500_ CPU.registerFile\[8\]\[29\] _08545_ _03552_ _03268_ VGND VGND VPWR VPWR _03553_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14163__301 clknet_1_1__leaf__08500_ VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__inv_2
X_12712_ _06636_ net2471 _08040_ VGND VGND VPWR VPWR _08050_ sky130_fd_sc_hd__mux2_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16480_ _03985_ _03986_ CPU.registerFile\[1\]\[11\] VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15431_ CPU.registerFile\[6\]\[27\] CPU.registerFile\[7\]\[27\] _08536_ VGND VGND
+ VPWR VPWR _03486_ sky130_fd_sc_hd__mux2_1
X_12643_ _08013_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18150_ net1161 _01678_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15362_ CPU.registerFile\[2\]\[25\] CPU.registerFile\[3\]\[25\] _03275_ VGND VGND
+ VPWR VPWR _03419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12574_ net2620 _07349_ _07968_ VGND VGND VPWR VPWR _07977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17101_ _04793_ _04801_ _04542_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__o21a_1
XFILLER_0_142_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14313_ CPU.registerFile\[15\]\[0\] CPU.registerFile\[14\]\[0\] _08558_ VGND VGND
+ VPWR VPWR _08559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11525_ net1900 _07309_ _07379_ VGND VGND VPWR VPWR _07380_ sky130_fd_sc_hd__mux2_1
X_18081_ net1092 _01609_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15293_ _03230_ _03347_ _03351_ _03151_ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__o211a_1
X_17032_ CPU.registerFile\[10\]\[25\] CPU.registerFile\[11\]\[25\] _06173_ VGND VGND
+ VPWR VPWR _04734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11456_ _07311_ VGND VGND VPWR VPWR _07333_ sky130_fd_sc_hd__buf_4
XFILLER_0_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10407_ _05736_ CPU.writeBack _05735_ VGND VGND VPWR VPWR _06663_ sky130_fd_sc_hd__and3b_4
X_14175_ clknet_1_1__leaf__08495_ VGND VGND VPWR VPWR _08502_ sky130_fd_sc_hd__buf_1
X_11387_ net2050 _06169_ _07285_ VGND VGND VPWR VPWR _07291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13126_ net1448 CPU.cycles\[1\] net1569 VGND VGND VPWR VPWR _08270_ sky130_fd_sc_hd__a21oi_1
X_10338_ _06616_ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__clkbuf_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ clknet_leaf_18_clk _02503_ VGND VGND VPWR VPWR CPU.aluIn1\[0\] sky130_fd_sc_hd__dfxtp_4
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ net1973 _06168_ _08228_ VGND VGND VPWR VPWR _08234_ sky130_fd_sc_hd__mux2_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ net945 _01462_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_10269_ _06574_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__clkbuf_1
X_12008_ _07637_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17865_ clknet_leaf_25_clk _00045_ VGND VGND VPWR VPWR CPU.cycles\[8\] sky130_fd_sc_hd__dfxtp_1
X_16816_ _04502_ _04510_ _04514_ _04523_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__a31o_2
XFILLER_0_88_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17796_ net876 _01358_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16747_ _04141_ _04437_ _04456_ _04096_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__a211o_1
XFILLER_0_159_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16678_ _05689_ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18417_ net238 _01945_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09150_ _05397_ CPU.aluIn1\[26\] VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__and2b_1
X_18348_ net169 _01876_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18279_ net1290 _01807_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_09081_ _05270_ CPU.aluIn1\[2\] VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold801 CPU.registerFile\[17\]\[14\] VGND VGND VPWR VPWR net2098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold812 CPU.registerFile\[21\]\[19\] VGND VGND VPWR VPWR net2109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 CPU.registerFile\[31\]\[27\] VGND VGND VPWR VPWR net2120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold834 CPU.registerFile\[3\]\[16\] VGND VGND VPWR VPWR net2131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold845 CPU.registerFile\[26\]\[10\] VGND VGND VPWR VPWR net2142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 CPU.registerFile\[9\]\[28\] VGND VGND VPWR VPWR net2153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 CPU.registerFile\[26\]\[8\] VGND VGND VPWR VPWR net2164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 CPU.registerFile\[18\]\[9\] VGND VGND VPWR VPWR net2175 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ _06202_ net1352 _06177_ VGND VGND VPWR VPWR _06314_ sky130_fd_sc_hd__o21a_1
Xhold889 CPU.registerFile\[31\]\[13\] VGND VGND VPWR VPWR net2186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08934_ _05284_ _05285_ VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__xor2_2
XFILLER_0_98_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13519__911 clknet_1_1__leaf__08436_ VGND VGND VPWR VPWR net967 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__03690_ clknet_0__03690_ VGND VGND VPWR VPWR clknet_1_0__leaf__03690_
+ sky130_fd_sc_hd__clkbuf_16
X_13969__126 clknet_1_1__leaf__08481_ VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__inv_2
XFILLER_0_79_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09417_ net2396 _05767_ _05742_ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09348_ _05584_ _05573_ VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__or2b_1
XFILLER_0_81_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09279_ CPU.aluIn1\[20\] _05544_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11310_ _07250_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12290_ mapped_spi_ram.rcv_data\[5\] _07813_ VGND VGND VPWR VPWR _07820_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11241_ _07213_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11172_ net1401 _07160_ _07169_ _07164_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__o211a_1
X_10123_ CPU.aluIn1\[4\] _05287_ _05769_ _06447_ VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__a31o_1
X_15980_ _08393_ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__clkbuf_4
X_14931_ _08522_ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__buf_4
X_10054_ _05910_ VGND VGND VPWR VPWR _06382_ sky130_fd_sc_hd__inv_2
X_14862_ _08764_ _02927_ _02930_ _02814_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__a211o_2
X_17650_ _04987_ _05187_ _04986_ _03659_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__a211o_1
X_16601_ _04098_ _04300_ _04304_ _04313_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__a31o_4
X_14087__232 clknet_1_0__leaf__08493_ VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__inv_2
X_17581_ _04996_ _05142_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__and2_1
X_14793_ _08549_ VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16532_ _04075_ _04241_ _04246_ _04042_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10956_ _06982_ VGND VGND VPWR VPWR _07008_ sky130_fd_sc_hd__buf_2
XFILLER_0_156_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16463_ _06109_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10887_ CPU.aluReg\[6\] CPU.aluReg\[4\] _06939_ VGND VGND VPWR VPWR _06955_ sky130_fd_sc_hd__mux2_1
X_15414_ CPU.registerFile\[30\]\[27\] CPU.registerFile\[31\]\[27\] _03291_ VGND VGND
+ VPWR VPWR _03469_ sky130_fd_sc_hd__mux2_1
X_18202_ net1213 net1344 VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[3\] sky130_fd_sc_hd__dfxtp_1
X_12626_ _06617_ net2165 _08004_ VGND VGND VPWR VPWR _08005_ sky130_fd_sc_hd__mux2_1
X_19182_ clknet_leaf_0_clk _02700_ VGND VGND VPWR VPWR per_uart.uart0.rx_ack sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16394_ CPU.registerFile\[5\]\[9\] CPU.registerFile\[4\]\[9\] _04024_ VGND VGND VPWR
+ VPWR _04112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18133_ net1144 _01661_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_15345_ CPU.registerFile\[27\]\[25\] CPU.registerFile\[26\]\[25\] _03172_ VGND VGND
+ VPWR VPWR _03402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12557_ _07956_ VGND VGND VPWR VPWR _07968_ sky130_fd_sc_hd__buf_4
XFILLER_0_81_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18064_ net1075 _01592_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_11508_ _06464_ VGND VGND VPWR VPWR _07368_ sky130_fd_sc_hd__clkbuf_4
X_15276_ _02964_ _03330_ _03334_ _03092_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__o211a_1
X_12488_ _07919_ VGND VGND VPWR VPWR _07931_ sky130_fd_sc_hd__buf_4
Xhold108 CPU.aluReg\[12\] VGND VGND VPWR VPWR net1405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17015_ _04716_ _04717_ _06535_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__mux2_1
Xhold119 mapped_spi_flash.rcv_data\[22\] VGND VGND VPWR VPWR net1416 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11439_ _07321_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__03653_ clknet_0__03653_ VGND VGND VPWR VPWR clknet_1_1__leaf__03653_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__03684_ _03684_ VGND VGND VPWR VPWR clknet_0__03684_ sky130_fd_sc_hd__clkbuf_16
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _06973_ net1573 VGND VGND VPWR VPWR _08261_ sky130_fd_sc_hd__nand2_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18966_ net740 _02486_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_13323__822 clknet_1_0__leaf__08364_ VGND VGND VPWR VPWR net878 sky130_fd_sc_hd__inv_2
XFILLER_0_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917_ clknet_leaf_17_clk _01445_ VGND VGND VPWR VPWR CPU.Iimm\[4\] sky130_fd_sc_hd__dfxtp_2
X_18897_ net671 _02417_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17848_ net928 _01410_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_17779_ net859 _01341_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13778__1143 clknet_1_1__leaf__08463_ VGND VGND VPWR VPWR net1199 sky130_fd_sc_hd__inv_2
XFILLER_0_45_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09202_ _05545_ _05550_ _05553_ CPU.cycles\[31\] VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15842__590 clknet_1_1__leaf__03679_ VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__inv_2
X_09133_ _05352_ _05483_ _05484_ VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09064_ CPU.rs2\[31\] _05247_ _05251_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold620 CPU.registerFile\[2\]\[18\] VGND VGND VPWR VPWR net1917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold631 CPU.registerFile\[30\]\[20\] VGND VGND VPWR VPWR net1928 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold642 CPU.registerFile\[19\]\[7\] VGND VGND VPWR VPWR net1939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold653 CPU.registerFile\[27\]\[11\] VGND VGND VPWR VPWR net1950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 CPU.registerFile\[3\]\[21\] VGND VGND VPWR VPWR net1961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 CPU.registerFile\[17\]\[0\] VGND VGND VPWR VPWR net1972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 CPU.registerFile\[15\]\[6\] VGND VGND VPWR VPWR net1983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 CPU.registerFile\[7\]\[10\] VGND VGND VPWR VPWR net1994 sky130_fd_sc_hd__dlygate4sd3_1
X_09966_ _05263_ _05265_ _05307_ _05308_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__o31a_1
X_08917_ CPU.aluIn1\[3\] _05268_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__and2_1
X_14036__186 clknet_1_0__leaf__08488_ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__inv_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _06126_ _06230_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__nand2_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1320 CPU.aluIn1\[26\] VGND VGND VPWR VPWR net2617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1331 CPU.registerFile\[25\]\[5\] VGND VGND VPWR VPWR net2628 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13595__979 clknet_1_0__leaf__08444_ VGND VGND VPWR VPWR net1035 sky130_fd_sc_hd__inv_2
Xhold1342 CPU.registerFile\[25\]\[8\] VGND VGND VPWR VPWR net2639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1353 CPU.PC\[22\] VGND VGND VPWR VPWR net2650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1364 CPU.aluIn1\[0\] VGND VGND VPWR VPWR net2661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1375 CPU.aluReg\[13\] VGND VGND VPWR VPWR net2672 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _06896_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__clkbuf_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13859__1217 clknet_1_1__leaf__08470_ VGND VGND VPWR VPWR net1273 sky130_fd_sc_hd__inv_2
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11790_ _06655_ net2407 _07512_ VGND VGND VPWR VPWR _07521_ sky130_fd_sc_hd__mux2_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10741_ net2470 _06413_ _06838_ VGND VGND VPWR VPWR _06844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13460_ _08418_ VGND VGND VPWR VPWR _08419_ sky130_fd_sc_hd__buf_6
XFILLER_0_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10672_ net2637 _06440_ _06799_ VGND VGND VPWR VPWR _06806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15624__426 clknet_1_0__leaf__03640_ VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__inv_2
X_12411_ _07890_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__clkbuf_1
X_13391_ _05577_ _05695_ _05579_ _05515_ VGND VGND VPWR VPWR _08374_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_899 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15130_ CPU.registerFile\[2\]\[19\] CPU.registerFile\[3\]\[19\] _02871_ VGND VGND
+ VPWR VPWR _03193_ sky130_fd_sc_hd__mux2_1
X_12342_ _06607_ net2105 _07848_ VGND VGND VPWR VPWR _07854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15061_ CPU.registerFile\[28\]\[18\] CPU.registerFile\[29\]\[18\] _02808_ VGND VGND
+ VPWR VPWR _03125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12273_ net1482 _07799_ _07810_ _07809_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__o211a_1
X_11224_ _07204_ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__clkbuf_1
X_18820_ net609 _02344_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_11155_ net1327 _07147_ _07159_ _07151_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10106_ _05286_ _06431_ VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__xnor2_1
X_18751_ net540 _02275_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[13\] sky130_fd_sc_hd__dfxtp_1
X_11086_ _06981_ _07110_ _07113_ _07115_ net1555 VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__a32o_1
X_17702_ _05207_ _05225_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__and2_1
X_14914_ _08409_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__buf_4
X_10037_ _05855_ _06203_ _06363_ _06204_ _06364_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__o32a_1
X_18682_ net471 _02206_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_17633_ net1965 VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__clkbuf_1
X_14845_ _02750_ _02896_ _02914_ _02839_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__a211o_1
XFILLER_0_86_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14776_ CPU.registerFile\[20\]\[11\] _08839_ _02846_ _08841_ VGND VGND VPWR VPWR
+ _02847_ sky130_fd_sc_hd__o211a_1
X_17564_ per_uart.tx_busy per_uart.uart0.tx_wr VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__and2b_1
X_11988_ _06649_ net2467 _07620_ VGND VGND VPWR VPWR _07626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16515_ CPU.registerFile\[5\]\[12\] CPU.registerFile\[4\]\[12\] _04024_ VGND VGND
+ VPWR VPWR _04230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10939_ _06996_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17495_ _05022_ _06230_ _05073_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16446_ _04161_ _04162_ _03875_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12609_ _06601_ net1832 _07993_ VGND VGND VPWR VPWR _07996_ sky130_fd_sc_hd__mux2_1
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19165_ clknet_leaf_0_clk _02685_ VGND VGND VPWR VPWR per_uart.rx_data\[4\] sky130_fd_sc_hd__dfxtp_1
X_16377_ _08596_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__buf_2
XFILLER_0_144_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15599__403 clknet_1_0__leaf__03638_ VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__inv_2
XFILLER_0_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_16
X_14141__281 clknet_1_1__leaf__08498_ VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__inv_2
XFILLER_0_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18116_ net1127 _01644_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_15328_ _03027_ _03383_ _03385_ _03111_ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__a211o_1
XFILLER_0_81_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19096_ net79 _02616_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18047_ net1058 _01575_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_15259_ _03155_ _03300_ _03318_ _03243_ VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__a211o_2
XFILLER_0_111_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09820_ _05343_ _05474_ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__xor2_1
X_09751_ _05357_ _06090_ _05354_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__a21oi_1
X_18949_ net723 _02469_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_09682_ _06021_ _06023_ _06024_ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__or3_1
XFILLER_0_146_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13293__795 clknet_1_0__leaf__08361_ VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__inv_2
XFILLER_0_71_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09116_ _05322_ CPU.aluIn1\[13\] VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09047_ CPU.aluIn1\[26\] _05397_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold450 CPU.registerFile\[28\]\[22\] VGND VGND VPWR VPWR net1747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 CPU.registerFile\[10\]\[22\] VGND VGND VPWR VPWR net1758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 CPU.registerFile\[13\]\[7\] VGND VGND VPWR VPWR net1769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 CPU.registerFile\[10\]\[8\] VGND VGND VPWR VPWR net1780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 CPU.registerFile\[6\]\[4\] VGND VGND VPWR VPWR net1791 sky130_fd_sc_hd__dlygate4sd3_1
X_13603__986 clknet_1_0__leaf__08445_ VGND VGND VPWR VPWR net1042 sky130_fd_sc_hd__inv_2
X_09949_ _05976_ _05943_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__and2b_1
X_12960_ net1725 _07314_ _08181_ VGND VGND VPWR VPWR _08183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1150 CPU.registerFile\[31\]\[21\] VGND VGND VPWR VPWR net2447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1161 CPU.registerFile\[2\]\[5\] VGND VGND VPWR VPWR net2458 sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ _07585_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__clkbuf_1
Xhold1172 CPU.registerFile\[25\]\[24\] VGND VGND VPWR VPWR net2469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 CPU.registerFile\[2\]\[12\] VGND VGND VPWR VPWR net2480 sky130_fd_sc_hd__dlygate4sd3_1
X_12891_ _08146_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__clkbuf_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 CPU.registerFile\[21\]\[11\] VGND VGND VPWR VPWR net2491 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ CPU.registerFile\[0\]\[7\] _08706_ _08868_ _08588_ VGND VGND VPWR VPWR _08869_
+ sky130_fd_sc_hd__o211a_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ net1760 _07353_ _07548_ VGND VGND VPWR VPWR _07549_ sky130_fd_sc_hd__mux2_1
X_15849__596 clknet_1_1__leaf__03680_ VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__inv_2
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03656_ clknet_0__03656_ VGND VGND VPWR VPWR clknet_1_0__leaf__03656_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ CPU.registerFile\[20\]\[6\] _08527_ _08800_ _08530_ VGND VGND VPWR VPWR _08801_
+ sky130_fd_sc_hd__o211a_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _07489_ VGND VGND VPWR VPWR _07512_ sky130_fd_sc_hd__clkbuf_4
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ CPU.registerFile\[12\]\[7\] _04017_ _04018_ _04019_ VGND VGND VPWR VPWR _04020_
+ sky130_fd_sc_hd__o211a_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17280_ _03735_ _04971_ _04975_ _03732_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__o211a_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ net2156 _06224_ _06827_ VGND VGND VPWR VPWR _06835_ sky130_fd_sc_hd__mux2_1
X_14492_ _08732_ _08733_ _08695_ VGND VGND VPWR VPWR _08734_ sky130_fd_sc_hd__mux2_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14199__333 clknet_1_0__leaf__08504_ VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__inv_2
X_16231_ CPU.registerFile\[27\]\[5\] CPU.registerFile\[26\]\[5\] _03837_ VGND VGND
+ VPWR VPWR _03953_ sky130_fd_sc_hd__mux2_1
X_13443_ _08405_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__clkbuf_1
X_10655_ net2427 _06245_ _06788_ VGND VGND VPWR VPWR _06797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16162_ CPU.registerFile\[19\]\[3\] CPU.registerFile\[18\]\[3\] _03767_ VGND VGND
+ VPWR VPWR _03886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10586_ _06759_ VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15113_ CPU.registerFile\[24\]\[19\] _02928_ _03174_ _03175_ VGND VGND VPWR VPWR
+ _03176_ sky130_fd_sc_hd__o211a_1
X_12325_ _07842_ _07838_ net1304 mapped_spi_ram.rcv_bitcount\[2\] VGND VGND VPWR VPWR
+ _01684_ sky130_fd_sc_hd__a22o_1
X_16093_ CPU.registerFile\[8\]\[2\] _08394_ _06150_ _03817_ VGND VGND VPWR VPWR _03818_
+ sky130_fd_sc_hd__o211a_1
X_15044_ _02831_ _02832_ CPU.registerFile\[1\]\[17\] VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12256_ net1524 _07799_ _07801_ _07796_ VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__o211a_1
X_11207_ _07188_ _07193_ net1433 VGND VGND VPWR VPWR _07194_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12187_ mapped_spi_ram.cmd_addr\[2\] _07749_ _07706_ CPU.mem_wdata\[3\] _07739_ VGND
+ VGND VPWR VPWR _07753_ sky130_fd_sc_hd__a221o_1
X_13777__1142 clknet_1_1__leaf__08463_ VGND VGND VPWR VPWR net1198 sky130_fd_sc_hd__inv_2
X_15594__399 clknet_1_1__leaf__08511_ VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__inv_2
X_18803_ net592 net1626 VGND VGND VPWR VPWR mapped_spi_flash.rbusy sky130_fd_sc_hd__dfxtp_1
X_11138_ _07001_ VGND VGND VPWR VPWR _07151_ sky130_fd_sc_hd__buf_2
X_16995_ CPU.aluIn1\[23\] _04458_ _04698_ _04663_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__o211a_1
X_13578__963 clknet_1_0__leaf__08443_ VGND VGND VPWR VPWR net1019 sky130_fd_sc_hd__inv_2
X_18734_ net523 _02258_ VGND VGND VPWR VPWR mapped_spi_flash.snd_bitcount\[2\] sky130_fd_sc_hd__dfxtp_1
X_11069_ _07048_ _07102_ VGND VGND VPWR VPWR _07103_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_0_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_16
X_18665_ net454 _02189_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_15877_ clknet_1_1__leaf__03654_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__buf_1
XFILLER_0_155_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17616_ per_uart.d_in_uart\[7\] _05157_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__nand2_1
X_14828_ CPU.registerFile\[13\]\[12\] CPU.registerFile\[12\]\[12\] _08693_ VGND VGND
+ VPWR VPWR _02898_ sky130_fd_sc_hd__mux2_1
X_18596_ net417 _02120_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17547_ CPU.PC\[23\] _05016_ _05114_ _05115_ _06858_ VGND VGND VPWR VPWR _02661_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_928 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14759_ _08566_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17478_ _05016_ CPU.PC\[10\] _05057_ _05059_ _05053_ VGND VGND VPWR VPWR _02648_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_128_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16429_ _03704_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19148_ clknet_leaf_5_clk _02668_ VGND VGND VPWR VPWR per_uart.uart0.tx_count16\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19079_ clknet_leaf_27_clk _02599_ VGND VGND VPWR VPWR per_uart.uart0.rxd_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13858__1216 clknet_1_1__leaf__08470_ VGND VGND VPWR VPWR net1272 sky130_fd_sc_hd__inv_2
X_15954__691 clknet_1_1__leaf__03690_ VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__inv_2
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09803_ _06140_ VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__buf_4
XFILLER_0_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09734_ _05366_ _05521_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__nor2_1
X_09665_ _05764_ _05877_ _05909_ _06008_ VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__a211o_4
XFILLER_0_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _05530_ _05922_ VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__nor2_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14148__287 clknet_1_1__leaf__08499_ VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__inv_2
XFILLER_0_77_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13699__1072 clknet_1_1__leaf__08455_ VGND VGND VPWR VPWR net1128 sky130_fd_sc_hd__inv_2
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10440_ _06681_ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10371_ _06596_ VGND VGND VPWR VPWR _06639_ sky130_fd_sc_hd__buf_4
XFILLER_0_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12110_ net1371 _07693_ _07700_ _07175_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__o211a_1
X_13090_ CPU.registerFile\[4\]\[0\] _06554_ _08216_ VGND VGND VPWR VPWR _08251_ sky130_fd_sc_hd__mux2_1
X_15736__527 clknet_1_1__leaf__03651_ VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__inv_2
X_12041_ _07654_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__clkbuf_1
Xhold280 CPU.rs2\[10\] VGND VGND VPWR VPWR net1577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold291 mapped_spi_flash.snd_bitcount\[4\] VGND VGND VPWR VPWR net1588 sky130_fd_sc_hd__dlygate4sd3_1
X_15800_ _08351_ _03668_ _03661_ VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__a21oi_1
X_16780_ _04479_ _04482_ _04488_ _04446_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__o211a_1
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ _08173_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18450_ net271 _01978_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_12874_ _06413_ net2249 _08131_ VGND VGND VPWR VPWR _08137_ sky130_fd_sc_hd__mux2_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11825_ net2392 _07337_ _07537_ VGND VGND VPWR VPWR _07540_ sky130_fd_sc_hd__mux2_1
X_14613_ _08722_ _08846_ _08850_ _08851_ VGND VGND VPWR VPWR _08852_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_917 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18381_ net202 _01909_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03639_ clknet_0__03639_ VGND VGND VPWR VPWR clknet_1_0__leaf__03639_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14544_ _08580_ VGND VGND VPWR VPWR _08785_ sky130_fd_sc_hd__clkbuf_4
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11756_ _07503_ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__clkbuf_1
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10707_ net2143 _06032_ _06816_ VGND VGND VPWR VPWR _06826_ sky130_fd_sc_hd__mux2_1
X_17263_ _03757_ _04954_ _04958_ _06109_ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__o211a_1
X_14475_ CPU.registerFile\[22\]\[4\] CPU.registerFile\[23\]\[4\] _08523_ VGND VGND
+ VPWR VPWR _08717_ sky130_fd_sc_hd__mux2_1
X_11687_ _07466_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19002_ clknet_leaf_12_clk _02522_ VGND VGND VPWR VPWR CPU.aluIn1\[19\] sky130_fd_sc_hd__dfxtp_2
X_16214_ CPU.registerFile\[15\]\[5\] CPU.registerFile\[14\]\[5\] _03705_ VGND VGND
+ VPWR VPWR _03936_ sky130_fd_sc_hd__mux2_1
X_13426_ _08392_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10638_ _06776_ VGND VGND VPWR VPWR _06788_ sky130_fd_sc_hd__buf_4
X_17194_ CPU.registerFile\[28\]\[29\] CPU.registerFile\[29\]\[29\] _03717_ VGND VGND
+ VPWR VPWR _04892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16145_ CPU.registerFile\[0\]\[3\] _03828_ _03725_ _03868_ VGND VGND VPWR VPWR _03869_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10569_ net2054 _06054_ _06750_ VGND VGND VPWR VPWR _06751_ sky130_fd_sc_hd__mux2_1
X_12308_ mapped_spi_ram.rcv_bitcount\[4\] _07781_ mapped_spi_ram.rcv_bitcount\[5\]
+ VGND VGND VPWR VPWR _07831_ sky130_fd_sc_hd__o21ai_1
X_16076_ CPU.registerFile\[24\]\[1\] _08393_ _03747_ _03801_ VGND VGND VPWR VPWR _03802_
+ sky130_fd_sc_hd__o211a_1
X_15027_ _06363_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__buf_4
X_12239_ net1431 _07785_ _07791_ _07755_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__o211a_1
X_16978_ CPU.registerFile\[28\]\[23\] CPU.registerFile\[29\]\[23\] _04526_ VGND VGND
+ VPWR VPWR _04682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput4 spi_miso_ram VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_2
X_18717_ net506 _02241_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[17\] sky130_fd_sc_hd__dfxtp_1
X_13359__854 clknet_1_0__leaf__08368_ VGND VGND VPWR VPWR net910 sky130_fd_sc_hd__inv_2
X_09450_ CPU.Jimm\[14\] VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__clkinv_4
X_18648_ clknet_leaf_11_clk _02172_ VGND VGND VPWR VPWR CPU.rs2\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09381_ _05542_ _05554_ _05732_ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__or3_4
X_18579_ net400 net36 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08488_ clknet_0__08488_ VGND VGND VPWR VPWR clknet_1_1__leaf__08488_
+ sky130_fd_sc_hd__clkbuf_16
X_09717_ _05659_ _05678_ _06057_ _05683_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__a211o_4
XFILLER_0_96_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09648_ _05991_ _05935_ _05989_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _05545_ _05922_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__and2_2
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14081__227 clknet_1_1__leaf__08492_ VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__inv_2
X_11610_ net2094 _07328_ _07416_ VGND VGND VPWR VPWR _07425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _07985_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11541_ net1698 _07328_ _07379_ VGND VGND VPWR VPWR _07388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11472_ net1915 _07343_ _07333_ VGND VGND VPWR VPWR _07344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13211_ _05800_ _06862_ _08324_ VGND VGND VPWR VPWR _08325_ sky130_fd_sc_hd__mux2_1
X_10423_ _06672_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13142_ CPU.cycles\[9\] _08277_ VGND VGND VPWR VPWR _08279_ sky130_fd_sc_hd__and2_1
X_10354_ _06627_ VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ net1333 VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__clkbuf_1
X_17950_ net961 _01478_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_10285_ net2285 _06337_ _06580_ VGND VGND VPWR VPWR _06583_ sky130_fd_sc_hd__mux2_1
X_12024_ _07645_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__clkbuf_1
X_16901_ CPU.registerFile\[28\]\[21\] CPU.registerFile\[29\]\[21\] _04526_ VGND VGND
+ VPWR VPWR _04607_ sky130_fd_sc_hd__mux2_1
X_17881_ clknet_leaf_20_clk _00031_ VGND VGND VPWR VPWR CPU.cycles\[24\] sky130_fd_sc_hd__dfxtp_1
X_16832_ _04367_ _04537_ _04539_ _04410_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__a211o_1
X_16763_ _06148_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__clkbuf_4
X_13975_ clknet_1_0__leaf__08473_ VGND VGND VPWR VPWR _08482_ sky130_fd_sc_hd__buf_1
X_18502_ net323 _02026_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_12926_ _08164_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__clkbuf_1
X_16694_ CPU.registerFile\[20\]\[16\] CPU.registerFile\[21\]\[16\] _04287_ VGND VGND
+ VPWR VPWR _04405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18433_ net254 _01961_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _06224_ net2122 _08120_ VGND VGND VPWR VPWR _08128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13857__1215 clknet_1_0__leaf__08470_ VGND VGND VPWR VPWR net1271 sky130_fd_sc_hd__inv_2
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ net2081 _07320_ _07526_ VGND VGND VPWR VPWR _07531_ sky130_fd_sc_hd__mux2_1
X_18364_ net185 _01892_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_15576_ _08533_ _03622_ _03626_ _08554_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__o211a_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _08090_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14527_ _08764_ _08765_ _08767_ _08552_ VGND VGND VPWR VPWR _08768_ sky130_fd_sc_hd__a211o_1
X_11739_ _07494_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18295_ net116 _01823_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17246_ _06085_ _04925_ _04942_ _08596_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__a211o_2
XFILLER_0_118_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14458_ _08557_ _08696_ _08700_ _08423_ VGND VGND VPWR VPWR _08701_ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0__08511_ _08511_ VGND VGND VPWR VPWR clknet_0__08511_ sky130_fd_sc_hd__clkbuf_16
X_13250__771 clknet_1_1__leaf__08343_ VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__inv_2
X_13409_ _08383_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__clkbuf_1
X_17177_ CPU.registerFile\[9\]\[29\] _03709_ VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14389_ _08574_ _08628_ _08633_ _08592_ VGND VGND VPWR VPWR _08634_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08442_ _08442_ VGND VGND VPWR VPWR clknet_0__08442_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__08342_ clknet_0__08342_ VGND VGND VPWR VPWR clknet_1_1__leaf__08342_
+ sky130_fd_sc_hd__clkbuf_16
X_16128_ _03842_ _03852_ _08406_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__o21a_1
X_08950_ _05284_ _05285_ _05287_ CPU.aluIn1\[4\] VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__a22o_1
X_16059_ CPU.registerFile\[12\]\[1\] _03707_ _03708_ _03784_ VGND VGND VPWR VPWR _03785_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08881_ net2 VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09502_ _05831_ _05846_ _05847_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09433_ mapped_spi_ram.rcv_data\[5\] _05761_ _05762_ net1381 VGND VGND VPWR VPWR
+ _05783_ sky130_fd_sc_hd__a22o_2
XFILLER_0_78_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18575__32 VGND VGND VPWR VPWR _18575__32/HI net32 sky130_fd_sc_hd__conb_1
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09364_ _05677_ _05663_ _05672_ _05715_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__nor4_1
XANTENNA_20 _04680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09295_ CPU.aluIn1\[22\] _05544_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__nor2_1
XANTENNA_31 _06124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_42 _08541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 clknet_1_0__leaf__08340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 CPU.mem_wdata\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13939__99 clknet_1_0__leaf__08478_ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__inv_2
XANTENNA_75 _08520_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10070_ _06206_ _06393_ _06394_ _06395_ _06396_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__a32o_1
Xclkbuf_1_0__f__08500_ clknet_0__08500_ VGND VGND VPWR VPWR clknet_1_0__leaf__08500_
+ sky130_fd_sc_hd__clkbuf_16
X_10972_ _07008_ _07019_ VGND VGND VPWR VPWR _07020_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_0__f__08362_ clknet_0__08362_ VGND VGND VPWR VPWR clknet_1_0__leaf__08362_
+ sky130_fd_sc_hd__clkbuf_16
X_12711_ _08049_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13946__105 clknet_1_1__leaf__08479_ VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__inv_2
XFILLER_0_155_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15430_ _03133_ _03480_ _03484_ _03188_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__o211a_1
X_12642_ _06634_ net1913 _08004_ VGND VGND VPWR VPWR _08013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15361_ _03416_ _03417_ _08562_ VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__mux2_1
X_12573_ _07976_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17100_ _04574_ _04796_ _04800_ _04584_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__o211a_1
X_11524_ _07378_ VGND VGND VPWR VPWR _07379_ sky130_fd_sc_hd__buf_4
X_14312_ _06061_ VGND VGND VPWR VPWR _08558_ sky130_fd_sc_hd__buf_4
XFILLER_0_80_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18080_ net1091 _01608_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_15292_ _03027_ _03348_ _03350_ _03111_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__a211o_1
XFILLER_0_81_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15894__637 clknet_1_0__leaf__03684_ VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__inv_2
XFILLER_0_123_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17031_ net2361 _04458_ _04733_ _04663_ VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__o211a_1
X_11455_ _06053_ VGND VGND VPWR VPWR _07332_ sky130_fd_sc_hd__buf_4
XFILLER_0_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10406_ _06662_ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11386_ _07290_ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__clkbuf_1
X_13125_ CPU.cycles\[0\] CPU.cycles\[1\] CPU.cycles\[2\] VGND VGND VPWR VPWR _08269_
+ sky130_fd_sc_hd__and3_1
X_10337_ _06615_ net1777 _06597_ VGND VGND VPWR VPWR _06616_ sky130_fd_sc_hd__mux2_1
X_18982_ net756 _02502_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13992__147 clknet_1_1__leaf__08483_ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__inv_2
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ net1336 VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__clkbuf_1
X_17933_ net944 _01461_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_10268_ net1690 _06145_ _06569_ VGND VGND VPWR VPWR _06574_ sky130_fd_sc_hd__mux2_1
X_12007_ net2144 _07314_ _07635_ VGND VGND VPWR VPWR _07637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17864_ clknet_leaf_25_clk _00044_ VGND VGND VPWR VPWR CPU.cycles\[7\] sky130_fd_sc_hd__dfxtp_1
X_10199_ CPU.aluIn1\[0\] _05276_ VGND VGND VPWR VPWR _06521_ sky130_fd_sc_hd__nand2_2
X_16815_ _04305_ _04517_ _04522_ _04476_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__o211a_1
X_17795_ net875 _01357_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_16746_ _04447_ _04455_ _04138_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__o21a_1
XFILLER_0_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12909_ _08155_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16677_ CPU.registerFile\[2\]\[16\] CPU.registerFile\[3\]\[16\] _04027_ VGND VGND
+ VPWR VPWR _04388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18416_ net237 _01944_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18347_ net168 _01875_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15559_ _08581_ _03607_ _03609_ _08535_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__04985_ clknet_0__04985_ VGND VGND VPWR VPWR clknet_1_1__leaf__04985_
+ sky130_fd_sc_hd__clkbuf_16
X_09080_ _05268_ CPU.aluIn1\[3\] VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__or2b_1
XFILLER_0_44_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18278_ net1289 _01806_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13839__1199 clknet_1_1__leaf__08468_ VGND VGND VPWR VPWR net1255 sky130_fd_sc_hd__inv_2
XFILLER_0_141_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17229_ CPU.registerFile\[30\]\[30\] CPU.registerFile\[31\]\[30\] _04605_ VGND VGND
+ VPWR VPWR _04926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold802 CPU.registerFile\[9\]\[25\] VGND VGND VPWR VPWR net2099 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold813 CPU.registerFile\[2\]\[28\] VGND VGND VPWR VPWR net2110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold824 CPU.registerFile\[27\]\[3\] VGND VGND VPWR VPWR net2121 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold835 CPU.registerFile\[11\]\[24\] VGND VGND VPWR VPWR net2132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold846 CPU.registerFile\[20\]\[22\] VGND VGND VPWR VPWR net2143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 CPU.registerFile\[9\]\[15\] VGND VGND VPWR VPWR net2154 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09982_ _06204_ _06311_ _06312_ _05855_ VGND VGND VPWR VPWR _06313_ sky130_fd_sc_hd__o22a_1
Xhold868 CPU.registerFile\[27\]\[21\] VGND VGND VPWR VPWR net2165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 CPU.registerFile\[20\]\[21\] VGND VGND VPWR VPWR net2176 sky130_fd_sc_hd__dlygate4sd3_1
X_08933_ CPU.mem_wdata\[5\] CPU.Bimm\[5\] _05245_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__mux2_4
XFILLER_0_110_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15689__484 clknet_1_0__leaf__03647_ VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__inv_2
XFILLER_0_79_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09416_ _05766_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__clkbuf_4
X_13257__777 clknet_1_1__leaf__08344_ VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__inv_2
X_09347_ mapped_spi_ram.rcv_data\[31\] _05685_ _05698_ net1398 VGND VGND VPWR VPWR
+ _05699_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_81_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09278_ CPU.aluIn1\[20\] _05544_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14193__328 clknet_1_0__leaf__08503_ VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__inv_2
X_11240_ _06617_ net1819 _07212_ VGND VGND VPWR VPWR _07213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11171_ net1648 _07134_ VGND VGND VPWR VPWR _07169_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13856__1214 clknet_1_0__leaf__08470_ VGND VGND VPWR VPWR net1270 sky130_fd_sc_hd__inv_2
X_10122_ _05289_ _05748_ _05535_ CPU.aluReg\[4\] VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10053_ _06380_ _05967_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__xnor2_1
X_14930_ _02751_ _02994_ _02996_ _02759_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__a211o_1
X_18236__20 VGND VGND VPWR VPWR _18236__20/HI net20 sky130_fd_sc_hd__conb_1
X_14861_ CPU.registerFile\[24\]\[13\] _02928_ _02929_ _02771_ VGND VGND VPWR VPWR
+ _02930_ sky130_fd_sc_hd__o211a_1
X_16600_ _04305_ _04308_ _04312_ _04072_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__o211a_1
X_14013__165 clknet_1_1__leaf__08486_ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__inv_2
X_17580_ _05141_ _05136_ _05138_ per_uart.uart0.tx_count16\[3\] VGND VGND VPWR VPWR
+ _05142_ sky130_fd_sc_hd__a22o_1
X_14792_ _02733_ _02734_ CPU.registerFile\[9\]\[11\] VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__a21o_1
X_13572__958 clknet_1_1__leaf__08442_ VGND VGND VPWR VPWR net1014 sky130_fd_sc_hd__inv_2
X_16531_ _04037_ _04243_ _04245_ _04208_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__a211o_1
X_10955_ _06999_ VGND VGND VPWR VPWR _07007_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0__f__08345_ clknet_0__08345_ VGND VGND VPWR VPWR clknet_1_0__leaf__08345_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16462_ _03963_ _04174_ _04178_ _04006_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__a211o_1
X_10886_ _06954_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18201_ net1212 _01729_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15413_ _08581_ _03465_ _03467_ _08535_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__a211o_1
XFILLER_0_156_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19181_ clknet_leaf_27_clk net1364 VGND VGND VPWR VPWR per_uart.uart0.uart_rxd2 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_72_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12625_ _07992_ VGND VGND VPWR VPWR _08004_ sky130_fd_sc_hd__buf_4
X_16393_ CPU.registerFile\[6\]\[9\] CPU.registerFile\[7\]\[9\] _04022_ VGND VGND VPWR
+ VPWR _04111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15902__644 clknet_1_0__leaf__03685_ VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__inv_2
XFILLER_0_26_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18132_ net1143 _01660_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_12556_ _07967_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__clkbuf_1
X_15344_ _03399_ _03400_ _03255_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11507_ _07367_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__clkbuf_1
X_18063_ net1074 _01591_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_15601__405 clknet_1_0__leaf__03638_ VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__inv_2
X_12487_ _07930_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__clkbuf_1
X_15275_ _03006_ _03331_ _03333_ _03218_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold109 _06266_ VGND VGND VPWR VPWR net1406 sky130_fd_sc_hd__dlygate4sd3_1
X_17014_ CPU.registerFile\[28\]\[24\] CPU.registerFile\[29\]\[24\] _04526_ VGND VGND
+ VPWR VPWR _04717_ sky130_fd_sc_hd__mux2_1
X_11438_ net1835 _07320_ _07312_ VGND VGND VPWR VPWR _07321_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__03652_ clknet_0__03652_ VGND VGND VPWR VPWR clknet_1_1__leaf__03652_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__03683_ _03683_ VGND VGND VPWR VPWR clknet_0__03683_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11369_ _07281_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__clkbuf_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ _08256_ _06973_ VGND VGND VPWR VPWR _08260_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18965_ net739 _02485_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ net1642 VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__clkbuf_1
X_17916_ clknet_leaf_23_clk _01444_ VGND VGND VPWR VPWR CPU.Iimm\[3\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18896_ net670 _02416_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17847_ net927 _01409_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_17778_ net858 _01340_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16729_ CPU.registerFile\[28\]\[17\] CPU.registerFile\[29\]\[17\] _04122_ VGND VGND
+ VPWR VPWR _04439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09201_ _05552_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__buf_2
XFILLER_0_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09132_ _05348_ CPU.aluIn1\[19\] VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__or2b_1
XFILLER_0_162_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13549__938 clknet_1_1__leaf__08439_ VGND VGND VPWR VPWR net994 sky130_fd_sc_hd__inv_2
XFILLER_0_161_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09063_ _05255_ _05259_ _05411_ _05414_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__o31a_1
XFILLER_0_13_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold610 CPU.registerFile\[3\]\[18\] VGND VGND VPWR VPWR net1907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 CPU.registerFile\[13\]\[21\] VGND VGND VPWR VPWR net1918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold632 CPU.registerFile\[15\]\[25\] VGND VGND VPWR VPWR net1929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold643 CPU.registerFile\[31\]\[11\] VGND VGND VPWR VPWR net1940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 CPU.registerFile\[17\]\[2\] VGND VGND VPWR VPWR net1951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 mapped_spi_flash.rcv_data\[14\] VGND VGND VPWR VPWR net1962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 CPU.registerFile\[4\]\[16\] VGND VGND VPWR VPWR net1973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 CPU.registerFile\[21\]\[27\] VGND VGND VPWR VPWR net1984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 CPU.registerFile\[22\]\[8\] VGND VGND VPWR VPWR net1995 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ _06273_ _06295_ VGND VGND VPWR VPWR _06296_ sky130_fd_sc_hd__and2_1
Xclkbuf_0__08339_ _08339_ VGND VGND VPWR VPWR clknet_0__08339_ sky130_fd_sc_hd__clkbuf_16
X_08916_ CPU.mem_wdata\[3\] CPU.Iimm\[3\] _05244_ VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__mux2_2
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _05457_ _06229_ VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__xnor2_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13298__800 clknet_1_1__leaf__08361_ VGND VGND VPWR VPWR net856 sky130_fd_sc_hd__inv_2
Xhold1310 CPU.aluReg\[31\] VGND VGND VPWR VPWR net2607 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1321 CPU.registerFile\[2\]\[9\] VGND VGND VPWR VPWR net2618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1332 CPU.registerFile\[1\]\[16\] VGND VGND VPWR VPWR net2629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1343 CPU.registerFile\[1\]\[3\] VGND VGND VPWR VPWR net2640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_528 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1354 mapped_spi_flash.snd_bitcount\[2\] VGND VGND VPWR VPWR net2651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1365 CPU.aluReg\[18\] VGND VGND VPWR VPWR net2662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1376 per_uart.uart0.rx_busy VGND VGND VPWR VPWR net2673 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ _06843_ VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10671_ _06805_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12410_ net1824 _07322_ _07884_ VGND VGND VPWR VPWR _07890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13390_ _08373_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14201__335 clknet_1_0__leaf__08504_ VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__inv_2
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12341_ _07853_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15060_ CPU.registerFile\[30\]\[18\] CPU.registerFile\[31\]\[18\] _02887_ VGND VGND
+ VPWR VPWR _03124_ sky130_fd_sc_hd__mux2_1
X_12272_ mapped_spi_ram.rcv_data\[13\] _07800_ VGND VGND VPWR VPWR _07810_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11223_ _06601_ net1989 _07201_ VGND VGND VPWR VPWR _07204_ sky130_fd_sc_hd__mux2_1
X_11154_ _06057_ _07132_ VGND VGND VPWR VPWR _07159_ sky130_fd_sc_hd__nand2_1
X_10105_ _05289_ _06429_ _06430_ VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__o21ai_1
X_18750_ net539 _02274_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11085_ _07009_ net16 _07114_ VGND VGND VPWR VPWR _07115_ sky130_fd_sc_hd__o21bai_1
X_17701_ CPU.mem_wdata\[3\] per_uart.d_in_uart\[3\] _05218_ VGND VGND VPWR VPWR _05225_
+ sky130_fd_sc_hd__mux2_1
X_14913_ _02728_ _02976_ _02980_ _02784_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__o211a_1
X_10036_ _05699_ _05720_ VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__nand2_1
X_18681_ net470 _02205_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_13838__1198 clknet_1_0__leaf__08468_ VGND VGND VPWR VPWR net1254 sky130_fd_sc_hd__inv_2
X_17632_ net1964 per_uart.uart0.rxd_reg\[6\] _05170_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__mux2_1
X_14844_ _02905_ _02913_ _02837_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__o21a_2
X_17563_ net2619 per_uart.tx_busy _05128_ _05120_ _06858_ VGND VGND VPWR VPWR _02664_
+ sky130_fd_sc_hd__o221a_1
X_14775_ CPU.registerFile\[21\]\[11\] _08718_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__or2_1
X_11987_ _07625_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16514_ CPU.registerFile\[6\]\[12\] CPU.registerFile\[7\]\[12\] _04022_ VGND VGND
+ VPWR VPWR _04229_ sky130_fd_sc_hd__mux2_1
X_17494_ CPU.state\[1\] VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__buf_2
X_10938_ _06992_ _06995_ VGND VGND VPWR VPWR _06996_ sky130_fd_sc_hd__and2_1
X_15826__575 clknet_1_1__leaf__03678_ VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__inv_2
X_13353__849 clknet_1_0__leaf__08367_ VGND VGND VPWR VPWR net905 sky130_fd_sc_hd__inv_2
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16445_ CPU.registerFile\[28\]\[10\] CPU.registerFile\[29\]\[10\] _04122_ VGND VGND
+ VPWR VPWR _04162_ sky130_fd_sc_hd__mux2_1
X_10869_ CPU.aluReg\[10\] _06941_ _06922_ VGND VGND VPWR VPWR _06942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12608_ _07995_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__clkbuf_1
X_19164_ clknet_leaf_0_clk _02684_ VGND VGND VPWR VPWR per_uart.rx_data\[3\] sky130_fd_sc_hd__dfxtp_1
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16376_ _04085_ _04094_ _08406_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__o21a_1
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18115_ net1126 _01643_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15327_ CPU.registerFile\[0\]\[24\] _08411_ _03384_ _03195_ VGND VGND VPWR VPWR _03385_
+ sky130_fd_sc_hd__o211a_1
X_12539_ net2360 _07314_ _07957_ VGND VGND VPWR VPWR _07959_ sky130_fd_sc_hd__mux2_1
X_19095_ net78 _02615_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14176__312 clknet_1_0__leaf__08502_ VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__inv_2
XFILLER_0_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18046_ net1057 _01574_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_15258_ _03309_ _03317_ _03241_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__o21a_2
XFILLER_0_151_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15189_ CPU.registerFile\[21\]\[21\] _02960_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_74 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09750_ _05344_ _05347_ _05358_ VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__o21a_1
X_18948_ net722 _02468_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09681_ _05379_ _05521_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__nor2_1
X_18879_ net653 _02399_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_13555__942 clknet_1_1__leaf__08441_ VGND VGND VPWR VPWR net998 sky130_fd_sc_hd__inv_2
XFILLER_0_89_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13855__1213 clknet_1_0__leaf__08470_ VGND VGND VPWR VPWR net1269 sky130_fd_sc_hd__inv_2
XFILLER_0_17_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09115_ _05466_ _05458_ VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__and2b_1
XFILLER_0_127_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09046_ CPU.aluIn1\[26\] _05397_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold440 CPU.registerFile\[5\]\[20\] VGND VGND VPWR VPWR net1737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 CPU.registerFile\[27\]\[9\] VGND VGND VPWR VPWR net1748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 CPU.registerFile\[28\]\[29\] VGND VGND VPWR VPWR net1759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 CPU.registerFile\[15\]\[13\] VGND VGND VPWR VPWR net1770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 CPU.registerFile\[27\]\[19\] VGND VGND VPWR VPWR net1781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 CPU.registerFile\[19\]\[26\] VGND VGND VPWR VPWR net1792 sky130_fd_sc_hd__dlygate4sd3_1
X_15931__670 clknet_1_0__leaf__03688_ VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__inv_2
X_09948_ _05315_ _06269_ _06270_ _06279_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__a211o_1
X_09879_ _06184_ _06213_ _05425_ VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__a21oi_1
Xhold1140 CPU.registerFile\[20\]\[4\] VGND VGND VPWR VPWR net2437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 CPU.registerFile\[23\]\[15\] VGND VGND VPWR VPWR net2448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 CPU.registerFile\[7\]\[26\] VGND VGND VPWR VPWR net2459 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ _06638_ net2445 _07584_ VGND VGND VPWR VPWR _07585_ sky130_fd_sc_hd__mux2_1
Xhold1173 CPU.registerFile\[20\]\[6\] VGND VGND VPWR VPWR net2470 sky130_fd_sc_hd__dlygate4sd3_1
X_12890_ _05734_ net2023 _08145_ VGND VGND VPWR VPWR _08146_ sky130_fd_sc_hd__mux2_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 CPU.registerFile\[29\]\[22\] VGND VGND VPWR VPWR net2481 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1195 CPU.registerFile\[12\]\[18\] VGND VGND VPWR VPWR net2492 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _07525_ VGND VGND VPWR VPWR _07548_ sky130_fd_sc_hd__buf_4
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03655_ clknet_0__03655_ VGND VGND VPWR VPWR clknet_1_0__leaf__03655_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14560_ CPU.registerFile\[21\]\[6\] _08718_ VGND VGND VPWR VPWR _08800_ sky130_fd_sc_hd__or2_1
X_11772_ _07511_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__clkbuf_1
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _06834_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__clkbuf_1
X_14491_ CPU.registerFile\[13\]\[4\] CPU.registerFile\[12\]\[4\] _08693_ VGND VGND
+ VPWR VPWR _08733_ sky130_fd_sc_hd__mux2_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14125__266 clknet_1_1__leaf__08497_ VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__inv_2
XFILLER_0_64_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16230_ _03950_ _03951_ _03875_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10654_ _06796_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__clkbuf_1
X_13442_ CPU.Jimm\[18\] _08404_ _08388_ VGND VGND VPWR VPWR _08405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16161_ _03882_ _03884_ _03763_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__mux2_1
X_10585_ net2337 _06245_ _06750_ VGND VGND VPWR VPWR _06759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15112_ _06035_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12324_ _07779_ _07843_ net1303 VGND VGND VPWR VPWR _07844_ sky130_fd_sc_hd__o21bai_1
X_16092_ CPU.registerFile\[9\]\[2\] _03698_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15043_ CPU.registerFile\[2\]\[17\] CPU.registerFile\[3\]\[17\] _02871_ VGND VGND
+ VPWR VPWR _03108_ sky130_fd_sc_hd__mux2_1
X_12255_ net1516 _07800_ VGND VGND VPWR VPWR _07801_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11206_ mapped_spi_flash.rcv_bitcount\[1\] mapped_spi_flash.rcv_bitcount\[0\] mapped_spi_flash.state\[3\]
+ VGND VGND VPWR VPWR _07193_ sky130_fd_sc_hd__o21a_1
X_12186_ net1355 _07738_ _07752_ _07737_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__o211a_1
X_11137_ net1593 _07149_ VGND VGND VPWR VPWR _07150_ sky130_fd_sc_hd__or2_1
X_18802_ net591 net1654 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfxtp_4
X_15713__506 clknet_1_0__leaf__03649_ VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__inv_2
X_14019__171 clknet_1_0__leaf__08486_ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__inv_2
X_16994_ _04545_ _04680_ _04697_ _04500_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__a211o_2
X_18733_ net522 _02257_ VGND VGND VPWR VPWR mapped_spi_flash.snd_bitcount\[1\] sky130_fd_sc_hd__dfxtp_1
X_11068_ mapped_spi_flash.cmd_addr\[2\] _05704_ _06976_ VGND VGND VPWR VPWR _07102_
+ sky130_fd_sc_hd__mux2_1
X_10019_ _05427_ _06347_ VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__nand2_1
X_18664_ net453 _02188_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_17615_ net1478 _05159_ _05165_ _07108_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__o22a_1
X_14827_ CPU.registerFile\[15\]\[12\] CPU.registerFile\[14\]\[12\] _08771_ VGND VGND
+ VPWR VPWR _02897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18595_ net416 net52 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_15908__650 clknet_1_1__leaf__03685_ VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__inv_2
X_17546_ _05904_ _05022_ _08255_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14758_ CPU.registerFile\[2\]\[10\] CPU.registerFile\[3\]\[10\] _08629_ VGND VGND
+ VPWR VPWR _02830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13709_ clknet_1_1__leaf__08451_ VGND VGND VPWR VPWR _08456_ sky130_fd_sc_hd__buf_1
X_17477_ _05058_ _06299_ _08255_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__a21bo_1
X_15607__411 clknet_1_1__leaf__03638_ VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__inv_2
XFILLER_0_156_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14689_ CPU.registerFile\[21\]\[9\] _08718_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__or2_1
X_16428_ _04099_ _04142_ _04144_ _04105_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__a211o_1
XFILLER_0_143_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19147_ clknet_leaf_5_clk _02667_ VGND VGND VPWR VPWR per_uart.uart0.tx_count16\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16359_ _04076_ _04077_ _03875_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_859 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19078_ net70 _02598_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18029_ net1040 _01557_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09802_ mapped_spi_ram.rcv_data\[9\] _05857_ _05859_ mapped_spi_flash.rcv_data\[9\]
+ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__a22o_4
Xclkbuf_0__03649_ _03649_ VGND VGND VPWR VPWR clknet_0__03649_ sky130_fd_sc_hd__clkbuf_16
X_09733_ _05363_ _05531_ _05534_ CPU.aluReg\[20\] _06073_ VGND VGND VPWR VPWR _06074_
+ sky130_fd_sc_hd__a221o_1
X_14230__361 clknet_1_0__leaf__08507_ VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__inv_2
X_09664_ _05912_ _06007_ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__nor2_1
X_09595_ CPU.PC\[13\] _05938_ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__xor2_2
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13837__1197 clknet_1_1__leaf__08468_ VGND VGND VPWR VPWR net1253 sky130_fd_sc_hd__inv_2
X_10370_ _06291_ VGND VGND VPWR VPWR _06638_ sky130_fd_sc_hd__buf_4
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09029_ _05367_ _05370_ _05374_ _05379_ _05380_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_14_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12040_ CPU.registerFile\[24\]\[14\] _07347_ _07646_ VGND VGND VPWR VPWR _07654_
+ sky130_fd_sc_hd__mux2_1
Xhold270 _01706_ VGND VGND VPWR VPWR net1567 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold281 mapped_spi_flash.rcv_data\[25\] VGND VGND VPWR VPWR net1578 sky130_fd_sc_hd__dlygate4sd3_1
X_13382__875 clknet_1_1__leaf__08370_ VGND VGND VPWR VPWR net931 sky130_fd_sc_hd__inv_2
Xhold292 CPU.rs2\[29\] VGND VGND VPWR VPWR net1589 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15730_ clknet_1_1__leaf__03643_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__buf_1
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12942_ _06413_ net2303 _08167_ VGND VGND VPWR VPWR _08173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _08136_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__clkbuf_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14612_ _08422_ VGND VGND VPWR VPWR _08851_ sky130_fd_sc_hd__clkbuf_4
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _07539_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__clkbuf_1
X_18380_ net201 _01908_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_929 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03638_ clknet_0__03638_ VGND VGND VPWR VPWR clknet_1_0__leaf__03638_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14207__341 clknet_1_1__leaf__08504_ VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__inv_2
XFILLER_0_96_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14543_ _08781_ _08782_ _08783_ VGND VGND VPWR VPWR _08784_ sky130_fd_sc_hd__mux2_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _06620_ net2475 _07501_ VGND VGND VPWR VPWR _07503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17262_ _03765_ _04955_ _04957_ _06141_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__a211o_1
X_10706_ _06825_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14474_ _08415_ _08713_ _08715_ _08420_ VGND VGND VPWR VPWR _08716_ sky130_fd_sc_hd__a211o_1
X_11686_ net2526 _07335_ _07464_ VGND VGND VPWR VPWR _07466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19001_ clknet_leaf_12_clk _02521_ VGND VGND VPWR VPWR CPU.aluIn1\[18\] sky130_fd_sc_hd__dfxtp_4
X_16213_ _08398_ _03932_ _03934_ _08401_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__a211o_1
X_13425_ _05514_ _06205_ _08388_ VGND VGND VPWR VPWR _08392_ sky130_fd_sc_hd__mux2_1
X_10637_ _06787_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__clkbuf_1
X_17193_ CPU.registerFile\[30\]\[29\] CPU.registerFile\[31\]\[29\] _04605_ VGND VGND
+ VPWR VPWR _04891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16144_ _03726_ _03727_ CPU.registerFile\[1\]\[3\] VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__a21o_1
X_13356_ clknet_1_1__leaf__08366_ VGND VGND VPWR VPWR _08368_ sky130_fd_sc_hd__buf_1
X_10568_ _06738_ VGND VGND VPWR VPWR _06750_ sky130_fd_sc_hd__buf_4
XFILLER_0_134_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15938__676 clknet_1_1__leaf__03689_ VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__inv_2
XFILLER_0_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12307_ net1323 VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__clkbuf_1
X_16075_ _03749_ _03751_ CPU.registerFile\[25\]\[1\] VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__a21o_1
X_10499_ _06701_ VGND VGND VPWR VPWR _06713_ sky130_fd_sc_hd__buf_4
X_15026_ _03006_ _03088_ _03090_ _02814_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12238_ mapped_spi_ram.rcv_data\[28\] _07787_ VGND VGND VPWR VPWR _07791_ sky130_fd_sc_hd__or2_1
X_12169_ mapped_spi_ram.cmd_addr\[9\] _05708_ _07724_ VGND VGND VPWR VPWR _07742_
+ sky130_fd_sc_hd__mux2_1
X_13854__1212 clknet_1_0__leaf__08470_ VGND VGND VPWR VPWR net1268 sky130_fd_sc_hd__inv_2
X_16977_ CPU.registerFile\[30\]\[23\] CPU.registerFile\[31\]\[23\] _04605_ VGND VGND
+ VPWR VPWR _04681_ sky130_fd_sc_hd__mux2_1
X_18716_ net505 _02240_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18647_ clknet_leaf_15_clk _02171_ VGND VGND VPWR VPWR CPU.rs2\[19\] sky130_fd_sc_hd__dfxtp_1
X_09380_ _05556_ _05687_ _05731_ VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__o21a_1
X_18578_ net399 net35 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17529_ _05055_ _06067_ _05061_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__or3_1
X_15683__479 clknet_1_1__leaf__03646_ VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__inv_2
X_17325__738 clknet_1_1__leaf__04982_ VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__inv_2
XFILLER_0_157_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08487_ clknet_0__08487_ VGND VGND VPWR VPWR clknet_1_1__leaf__08487_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14154__292 clknet_1_0__leaf__08500_ VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__inv_2
X_09716_ net1619 VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__inv_2
X_09647_ _05988_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__inv_2
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09578_ CPU.instr\[3\] CPU.instr\[4\] VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__nor2_2
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15742__532 clknet_1_1__leaf__03652_ VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__inv_2
XFILLER_0_136_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11540_ _07387_ VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11471_ _06168_ VGND VGND VPWR VPWR _07343_ sky130_fd_sc_hd__buf_4
XFILLER_0_107_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10422_ _06609_ net2413 _06665_ VGND VGND VPWR VPWR _06672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13210_ _05513_ _05816_ _08322_ _08323_ VGND VGND VPWR VPWR _08324_ sky130_fd_sc_hd__or4_1
XFILLER_0_104_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10353_ _06626_ net1930 _06618_ VGND VGND VPWR VPWR _06627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13141_ _08277_ net1544 VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__nor2_1
X_14237__367 clknet_1_1__leaf__08508_ VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__inv_2
X_13072_ CPU.registerFile\[4\]\[9\] net1332 _08239_ VGND VGND VPWR VPWR _08242_ sky130_fd_sc_hd__mux2_1
X_10284_ _06582_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__clkbuf_1
X_12023_ CPU.registerFile\[24\]\[22\] _07330_ _07635_ VGND VGND VPWR VPWR _07645_
+ sky130_fd_sc_hd__mux2_1
X_16900_ CPU.registerFile\[30\]\[21\] CPU.registerFile\[31\]\[21\] _04605_ VGND VGND
+ VPWR VPWR _04606_ sky130_fd_sc_hd__mux2_1
X_17880_ clknet_leaf_19_clk _00030_ VGND VGND VPWR VPWR CPU.cycles\[23\] sky130_fd_sc_hd__dfxtp_1
X_16831_ CPU.registerFile\[16\]\[19\] _04252_ _04494_ _04538_ VGND VGND VPWR VPWR
+ _04539_ sky130_fd_sc_hd__o211a_1
X_16762_ CPU.registerFile\[2\]\[18\] CPU.registerFile\[3\]\[18\] _04431_ VGND VGND
+ VPWR VPWR _04471_ sky130_fd_sc_hd__mux2_1
X_18501_ net322 _02025_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_12925_ _06224_ net2325 _08156_ VGND VGND VPWR VPWR _08164_ sky130_fd_sc_hd__mux2_1
X_16693_ CPU.registerFile\[22\]\[16\] CPU.registerFile\[23\]\[16\] _04362_ VGND VGND
+ VPWR VPWR _04404_ sky130_fd_sc_hd__mux2_1
X_18432_ net253 _01960_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _08127_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18363_ net184 _01891_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_11807_ _07530_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__clkbuf_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _08543_ _03623_ _03625_ _03307_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__a211o_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _06643_ net2317 _08087_ VGND VGND VPWR VPWR _08090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ CPU.registerFile\[24\]\[5\] _08686_ _08766_ _08550_ VGND VGND VPWR VPWR _08767_
+ sky130_fd_sc_hd__o211a_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ _06603_ net2262 _07490_ VGND VGND VPWR VPWR _07494_ sky130_fd_sc_hd__mux2_1
X_18294_ net115 _01822_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17245_ _04933_ _04941_ _06474_ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__o21a_1
X_14457_ _08520_ _08697_ _08699_ _08661_ VGND VGND VPWR VPWR _08700_ sky130_fd_sc_hd__a211o_1
X_11669_ net2359 _07318_ _07453_ VGND VGND VPWR VPWR _07457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__08510_ _08510_ VGND VGND VPWR VPWR clknet_0__08510_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13408_ CPU.instr\[6\] _06389_ _00000_ VGND VGND VPWR VPWR _08383_ sky130_fd_sc_hd__mux2_1
X_17176_ CPU.registerFile\[10\]\[29\] CPU.registerFile\[11\]\[29\] _06173_ VGND VGND
+ VPWR VPWR _04874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14388_ _08581_ _08630_ _08632_ _08590_ VGND VGND VPWR VPWR _08633_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__08441_ _08441_ VGND VGND VPWR VPWR clknet_0__08441_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__08341_ clknet_0__08341_ VGND VGND VPWR VPWR clknet_1_1__leaf__08341_
+ sky130_fd_sc_hd__clkbuf_16
X_16127_ _03758_ _03845_ _03851_ _03775_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15871__616 clknet_1_0__leaf__03682_ VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__inv_2
XFILLER_0_122_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16058_ CPU.registerFile\[13\]\[1\] _03709_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15009_ CPU.registerFile\[19\]\[17\] CPU.registerFile\[18\]\[17\] _02753_ VGND VGND
+ VPWR VPWR _03074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09501_ _05831_ _05846_ _05424_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__o21ai_1
X_13836__1196 clknet_1_1__leaf__08468_ VGND VGND VPWR VPWR net1252 sky130_fd_sc_hd__inv_2
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09432_ CPU.Bimm\[9\] _05758_ _05759_ CPU.cycles\[29\] VGND VGND VPWR VPWR _05782_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09363_ _05235_ _05710_ _05714_ VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09294_ CPU.aluIn1\[22\] _05544_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_10 _03495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18590__47 VGND VGND VPWR VPWR _18590__47/HI net47 sky130_fd_sc_hd__conb_1
XANTENNA_21 _04698_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 _06124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 _08794_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_54 clknet_1_0__leaf__08340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_65 CPU.mem_wdata\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_76 _08549_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10971_ mapped_spi_flash.cmd_addr\[16\] _05671_ _07009_ VGND VGND VPWR VPWR _07019_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__08361_ clknet_0__08361_ VGND VGND VPWR VPWR clknet_1_0__leaf__08361_
+ sky130_fd_sc_hd__clkbuf_16
X_12710_ _06634_ net2520 _08040_ VGND VGND VPWR VPWR _08049_ sky130_fd_sc_hd__mux2_1
X_15666__463 clknet_1_0__leaf__03645_ VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__inv_2
XFILLER_0_84_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17308__722 clknet_1_0__leaf__04981_ VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__inv_2
X_12641_ _08012_ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15360_ CPU.registerFile\[5\]\[25\] CPU.registerFile\[4\]\[25\] _03105_ VGND VGND
+ VPWR VPWR _03417_ sky130_fd_sc_hd__mux2_1
X_12572_ net2627 _07347_ _07968_ VGND VGND VPWR VPWR _07976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14311_ _08532_ VGND VGND VPWR VPWR _08557_ sky130_fd_sc_hd__buf_4
X_13234__756 clknet_1_1__leaf__08342_ VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__inv_2
X_11523_ _07236_ _07310_ VGND VGND VPWR VPWR _07378_ sky130_fd_sc_hd__nor2_4
X_15291_ CPU.registerFile\[0\]\[23\] _08411_ _03349_ _03195_ VGND VGND VPWR VPWR _03350_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17030_ _04545_ _04715_ _04732_ _04500_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__a211o_2
X_14242_ clknet_1_1__leaf__08506_ VGND VGND VPWR VPWR _08509_ sky130_fd_sc_hd__buf_1
XFILLER_0_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11454_ _07331_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10405_ _06661_ net2184 _06596_ VGND VGND VPWR VPWR _06662_ sky130_fd_sc_hd__mux2_1
X_11385_ net2009 _06145_ _07285_ VGND VGND VPWR VPWR _07290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13124_ net1448 net1609 VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__xor2_1
XFILLER_0_150_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10336_ _06031_ VGND VGND VPWR VPWR _06615_ sky130_fd_sc_hd__clkbuf_4
X_18981_ net755 _02501_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14170__307 clknet_1_1__leaf__08501_ VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__inv_2
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ CPU.registerFile\[4\]\[17\] _06144_ _08228_ VGND VGND VPWR VPWR _08233_ sky130_fd_sc_hd__mux2_1
X_17932_ net943 _01460_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_10267_ _06573_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__clkbuf_1
X_12006_ _07636_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__clkbuf_1
X_17863_ clknet_leaf_25_clk _00043_ VGND VGND VPWR VPWR CPU.cycles\[6\] sky130_fd_sc_hd__dfxtp_1
X_10198_ _06519_ _05438_ VGND VGND VPWR VPWR _06520_ sky130_fd_sc_hd__xnor2_1
X_16814_ _04347_ _04518_ _04520_ _04521_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__a211o_1
X_17794_ net874 _01356_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16745_ _04170_ _04450_ _04454_ _04180_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__o211a_1
X_12908_ _06032_ net2485 _08145_ VGND VGND VPWR VPWR _08155_ sky130_fd_sc_hd__mux2_1
X_16676_ _04385_ _04386_ _04153_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18415_ net236 _01943_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12839_ _08118_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18346_ net167 _01874_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15558_ CPU.registerFile\[20\]\[31\] _08523_ _03608_ _08578_ VGND VGND VPWR VPWR
+ _03609_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04984_ clknet_0__04984_ VGND VGND VPWR VPWR clknet_1_1__leaf__04984_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_44_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14509_ _07163_ VGND VGND VPWR VPWR _08751_ sky130_fd_sc_hd__clkbuf_4
X_18277_ net1288 _01805_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15489_ CPU.registerFile\[27\]\[29\] CPU.registerFile\[26\]\[29\] _08576_ VGND VGND
+ VPWR VPWR _03542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17228_ _03755_ _04912_ _04916_ _04924_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold803 CPU.registerFile\[7\]\[1\] VGND VGND VPWR VPWR net2100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 CPU.registerFile\[11\]\[20\] VGND VGND VPWR VPWR net2111 sky130_fd_sc_hd__dlygate4sd3_1
X_17159_ _04856_ _04857_ _06535_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__mux2_1
Xhold825 CPU.registerFile\[29\]\[14\] VGND VGND VPWR VPWR net2122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold836 CPU.registerFile\[19\]\[8\] VGND VGND VPWR VPWR net2133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 CPU.registerFile\[24\]\[30\] VGND VGND VPWR VPWR net2144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 CPU.registerFile\[28\]\[9\] VGND VGND VPWR VPWR net2155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 CPU.registerFile\[7\]\[27\] VGND VGND VPWR VPWR net2166 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ _05693_ _05827_ VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__or2_1
X_08932_ CPU.aluIn1\[5\] VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09415_ _05745_ _05757_ _05760_ _05765_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__a211o_4
XFILLER_0_109_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09346_ _05659_ _05678_ _05683_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_63_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09277_ _05563_ _05566_ _05626_ _05628_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13526__917 clknet_1_0__leaf__08437_ VGND VGND VPWR VPWR net973 sky130_fd_sc_hd__inv_2
X_11170_ net1381 _07160_ _07168_ _07164_ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10121_ _06443_ _06445_ _05800_ VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__a21oi_1
X_10052_ _05968_ _05947_ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__or2b_1
X_14860_ _08808_ _08809_ CPU.registerFile\[25\]\[13\] VGND VGND VPWR VPWR _02929_
+ sky130_fd_sc_hd__a21o_1
X_14791_ CPU.registerFile\[10\]\[11\] CPU.registerFile\[11\]\[11\] _02779_ VGND VGND
+ VPWR VPWR _02862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16530_ CPU.registerFile\[24\]\[12\] _03915_ _04165_ _04244_ VGND VGND VPWR VPWR
+ _04245_ sky130_fd_sc_hd__o211a_1
X_13742_ clknet_1_0__leaf__08451_ VGND VGND VPWR VPWR _08459_ sky130_fd_sc_hd__buf_1
X_10954_ _07006_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__08344_ clknet_0__08344_ VGND VGND VPWR VPWR clknet_1_0__leaf__08344_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16461_ CPU.registerFile\[16\]\[10\] _03848_ _04090_ _04177_ VGND VGND VPWR VPWR
+ _04178_ sky130_fd_sc_hd__o211a_1
X_10885_ net2575 _06953_ _06868_ VGND VGND VPWR VPWR _06954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18200_ net1211 net1315 VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[1\] sky130_fd_sc_hd__dfxtp_1
X_15412_ CPU.registerFile\[20\]\[27\] _08523_ _03466_ _08578_ VGND VGND VPWR VPWR
+ _03467_ sky130_fd_sc_hd__o211a_1
X_19180_ clknet_leaf_27_clk net1 VGND VGND VPWR VPWR per_uart.uart0.uart_rxd1 sky130_fd_sc_hd__dfxtp_1
X_12624_ _08003_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__clkbuf_1
X_16392_ _04015_ _04107_ _04109_ _03979_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13697__1071 clknet_1_1__leaf__08454_ VGND VGND VPWR VPWR net1127 sky130_fd_sc_hd__inv_2
X_18131_ net1142 _01659_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15343_ CPU.registerFile\[28\]\[25\] CPU.registerFile\[29\]\[25\] _03212_ VGND VGND
+ VPWR VPWR _03400_ sky130_fd_sc_hd__mux2_1
X_12555_ net2191 _07330_ _07957_ VGND VGND VPWR VPWR _07967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18062_ net1073 _01590_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_11506_ net1736 _07366_ _07354_ VGND VGND VPWR VPWR _07367_ sky130_fd_sc_hd__mux2_1
X_15274_ CPU.registerFile\[24\]\[23\] _08582_ _03332_ _03175_ VGND VGND VPWR VPWR
+ _03333_ sky130_fd_sc_hd__o211a_1
X_12486_ net2170 _07330_ _07920_ VGND VGND VPWR VPWR _07930_ sky130_fd_sc_hd__mux2_1
X_17013_ CPU.registerFile\[30\]\[24\] CPU.registerFile\[31\]\[24\] _04605_ VGND VGND
+ VPWR VPWR _04716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03651_ clknet_0__03651_ VGND VGND VPWR VPWR clknet_1_1__leaf__03651_
+ sky130_fd_sc_hd__clkbuf_16
X_11437_ net1339 VGND VGND VPWR VPWR _07320_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13835__1195 clknet_1_1__leaf__08468_ VGND VGND VPWR VPWR net1251 sky130_fd_sc_hd__inv_2
XFILLER_0_10_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__03682_ _03682_ VGND VGND VPWR VPWR clknet_0__03682_ sky130_fd_sc_hd__clkbuf_16
X_11368_ net1740 _05853_ _07274_ VGND VGND VPWR VPWR _07281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ _06980_ _08259_ _06856_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _06603_ net2021 _06597_ VGND VGND VPWR VPWR _06604_ sky130_fd_sc_hd__mux2_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18964_ net738 _02484_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _07244_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__clkbuf_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ CPU.registerFile\[4\]\[25\] _05852_ _08217_ VGND VGND VPWR VPWR _08224_ sky130_fd_sc_hd__mux2_1
X_17915_ clknet_leaf_14_clk _01443_ VGND VGND VPWR VPWR CPU.Iimm\[2\] sky130_fd_sc_hd__dfxtp_2
X_18895_ net669 _02415_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17846_ net926 _01408_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_17777_ net857 _01339_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_14989_ _02798_ _03039_ _03044_ _03054_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16728_ CPU.registerFile\[30\]\[17\] CPU.registerFile\[31\]\[17\] _04201_ VGND VGND
+ VPWR VPWR _04438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16659_ _04367_ _04368_ _04370_ _04006_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09200_ _05422_ _05538_ CPU.instr\[6\] _05551_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__and4_1
XFILLER_0_151_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09131_ _05356_ _05481_ _05482_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__a21oi_1
X_18329_ net150 _01857_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09062_ _05413_ VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold600 CPU.registerFile\[13\]\[17\] VGND VGND VPWR VPWR net1897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 CPU.registerFile\[6\]\[22\] VGND VGND VPWR VPWR net1908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold622 CPU.registerFile\[22\]\[13\] VGND VGND VPWR VPWR net1919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 CPU.registerFile\[15\]\[17\] VGND VGND VPWR VPWR net1930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold644 CPU.registerFile\[17\]\[6\] VGND VGND VPWR VPWR net1941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 CPU.registerFile\[30\]\[28\] VGND VGND VPWR VPWR net1952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold666 CPU.registerFile\[18\]\[4\] VGND VGND VPWR VPWR net1963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 CPU.registerFile\[30\]\[31\] VGND VGND VPWR VPWR net1974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 CPU.registerFile\[5\]\[24\] VGND VGND VPWR VPWR net1985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 CPU.registerFile\[21\]\[29\] VGND VGND VPWR VPWR net1996 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ _05310_ _05461_ _06272_ VGND VGND VPWR VPWR _06295_ sky130_fd_sc_hd__nand3_1
X_08915_ _05263_ _05266_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__or2_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ _05316_ _05321_ VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__nor2_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1300 CPU.registerFile\[12\]\[12\] VGND VGND VPWR VPWR net2597 sky130_fd_sc_hd__dlygate4sd3_1
X_13263__782 clknet_1_1__leaf__08345_ VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__inv_2
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1311 CPU.registerFile\[12\]\[15\] VGND VGND VPWR VPWR net2608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 per_uart.uart0.tx_wr VGND VGND VPWR VPWR net2619 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1333 CPU.PC\[13\] VGND VGND VPWR VPWR net2630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1344 CPU.PC\[12\] VGND VGND VPWR VPWR net2641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1355 CPU.registerFile\[2\]\[6\] VGND VGND VPWR VPWR net2652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1366 CPU.registerFile\[2\]\[8\] VGND VGND VPWR VPWR net2663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1377 mapped_spi_ram.state\[1\] VGND VGND VPWR VPWR net2674 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10670_ CPU.registerFile\[1\]\[6\] _06413_ _06799_ VGND VGND VPWR VPWR _06805_ sky130_fd_sc_hd__mux2_1
X_09329_ _05671_ _05667_ _05680_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__and3b_1
XFILLER_0_35_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12340_ _06605_ net1597 _07848_ VGND VGND VPWR VPWR _07853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15778__564 clknet_1_1__leaf__03656_ VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__inv_2
X_12271_ net1489 _07799_ _07808_ _07809_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17341__2 clknet_1_1__leaf__04984_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__inv_2
XFILLER_0_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11222_ _07203_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__clkbuf_1
X_13307__808 clknet_1_1__leaf__08362_ VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__inv_2
XFILLER_0_102_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11153_ net1619 _07147_ _07158_ _07151_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__o211a_1
X_13923__84 clknet_1_0__leaf__08477_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__inv_2
X_10104_ CPU.aluIn1\[4\] _05287_ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__nand2_1
X_11084_ _06981_ _07110_ VGND VGND VPWR VPWR _07114_ sky130_fd_sc_hd__nand2_2
X_14912_ _08857_ _02977_ _02979_ _02903_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__a211o_1
X_10035_ _05722_ _05723_ VGND VGND VPWR VPWR _06363_ sky130_fd_sc_hd__nand2_4
X_17700_ _05224_ VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__clkbuf_1
X_18680_ net469 _02204_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_14843_ _02826_ _02908_ _02912_ _02746_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__o211a_1
X_17631_ net1960 VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__clkbuf_1
X_17562_ _05117_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__inv_2
X_14774_ CPU.registerFile\[22\]\[11\] CPU.registerFile\[23\]\[11\] _08756_ VGND VGND
+ VPWR VPWR _02845_ sky130_fd_sc_hd__mux2_1
X_11986_ _06647_ net2457 _07620_ VGND VGND VPWR VPWR _07625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16513_ _04015_ _04225_ _04227_ _03979_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__a211o_1
XFILLER_0_105_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17493_ _05070_ _05071_ _05020_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__a21oi_1
X_10937_ mapped_spi_flash.cmd_addr\[27\] _06983_ _06985_ mapped_spi_flash.cmd_addr\[26\]
+ VGND VGND VPWR VPWR _06995_ sky130_fd_sc_hd__a22o_1
X_16444_ CPU.registerFile\[30\]\[10\] CPU.registerFile\[31\]\[10\] _03796_ VGND VGND
+ VPWR VPWR _04161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10868_ CPU.aluIn1\[10\] _06940_ _06914_ VGND VGND VPWR VPWR _06941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12607_ _06599_ net1744 _07993_ VGND VGND VPWR VPWR _07995_ sky130_fd_sc_hd__mux2_1
X_19163_ clknet_leaf_0_clk _02683_ VGND VGND VPWR VPWR per_uart.rx_data\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16375_ _03758_ _04088_ _04093_ _03775_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__o211a_1
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13587_ clknet_1_1__leaf__08440_ VGND VGND VPWR VPWR _08444_ sky130_fd_sc_hd__buf_1
XFILLER_0_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10799_ CPU.aluIn1\[26\] _06887_ _06881_ VGND VGND VPWR VPWR _06888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18114_ net1125 _01642_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_15326_ _03235_ _03236_ CPU.registerFile\[1\]\[24\] VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12538_ _07958_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19094_ net77 _02614_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18045_ net1056 _01573_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_15257_ _03230_ _03312_ _03316_ _03151_ VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__o211a_1
X_12469_ _07921_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14208_ clknet_1_0__leaf__08495_ VGND VGND VPWR VPWR _08505_ sky130_fd_sc_hd__buf_1
X_15188_ CPU.registerFile\[22\]\[21\] CPU.registerFile\[23\]\[21\] _02998_ VGND VGND
+ VPWR VPWR _03249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18947_ net721 _02467_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_09680_ _05376_ _05531_ _05534_ CPU.aluReg\[22\] _06022_ VGND VGND VPWR VPWR _06023_
+ sky130_fd_sc_hd__a221o_1
X_18878_ net652 _02398_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_17829_ net909 _01391_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_17423__44 clknet_1_1__leaf__05015_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__inv_2
XFILLER_0_76_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09114_ _05459_ _05312_ _05465_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09045_ CPU.rs2\[26\] _05247_ _05251_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__o21a_1
XFILLER_0_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold430 CPU.registerFile\[10\]\[2\] VGND VGND VPWR VPWR net1727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold441 CPU.registerFile\[28\]\[19\] VGND VGND VPWR VPWR net1738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 CPU.registerFile\[19\]\[12\] VGND VGND VPWR VPWR net1749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 CPU.registerFile\[9\]\[11\] VGND VGND VPWR VPWR net1760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold474 CPU.registerFile\[15\]\[26\] VGND VGND VPWR VPWR net1771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 CPU.registerFile\[11\]\[11\] VGND VGND VPWR VPWR net1782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 CPU.registerFile\[10\]\[12\] VGND VGND VPWR VPWR net1793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09947_ _06126_ _06275_ _06278_ _05818_ VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__o211a_1
X_13696__1070 clknet_1_1__leaf__08454_ VGND VGND VPWR VPWR net1126 sky130_fd_sc_hd__inv_2
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _05333_ _05468_ _06183_ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__or3_1
Xhold1130 CPU.registerFile\[1\]\[13\] VGND VGND VPWR VPWR net2427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 CPU.registerFile\[20\]\[27\] VGND VGND VPWR VPWR net2438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1152 CPU.registerFile\[23\]\[26\] VGND VGND VPWR VPWR net2449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1163 CPU.registerFile\[2\]\[2\] VGND VGND VPWR VPWR net2460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1174 CPU.registerFile\[25\]\[12\] VGND VGND VPWR VPWR net2471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 CPU.registerFile\[8\]\[3\] VGND VGND VPWR VPWR net2482 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1196 CPU.registerFile\[14\]\[6\] VGND VGND VPWR VPWR net2493 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _07547_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__clkbuf_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03654_ clknet_0__03654_ VGND VGND VPWR VPWR clknet_1_0__leaf__03654_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13834__1194 clknet_1_0__leaf__08468_ VGND VGND VPWR VPWR net1250 sky130_fd_sc_hd__inv_2
XFILLER_0_68_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _06636_ net1801 _07501_ VGND VGND VPWR VPWR _07511_ sky130_fd_sc_hd__mux2_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10722_ net1904 _06200_ _06827_ VGND VGND VPWR VPWR _06834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14490_ CPU.registerFile\[15\]\[4\] CPU.registerFile\[14\]\[4\] _08558_ VGND VGND
+ VPWR VPWR _08732_ sky130_fd_sc_hd__mux2_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13441_ _08403_ VGND VGND VPWR VPWR _08404_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10653_ net2565 _06224_ _06788_ VGND VGND VPWR VPWR _06796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16160_ CPU.registerFile\[20\]\[3\] CPU.registerFile\[21\]\[3\] _03883_ VGND VGND
+ VPWR VPWR _03884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10584_ _06758_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15111_ _03049_ _03050_ CPU.registerFile\[25\]\[19\] VGND VGND VPWR VPWR _03174_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12323_ mapped_spi_ram.rcv_bitcount\[1\] mapped_spi_ram.rcv_bitcount\[0\] VGND VGND
+ VPWR VPWR _07843_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16091_ CPU.registerFile\[10\]\[2\] CPU.registerFile\[11\]\[2\] _03694_ VGND VGND
+ VPWR VPWR _03816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15042_ _03104_ _03106_ _03025_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__mux2_1
X_12254_ _07786_ VGND VGND VPWR VPWR _07800_ sky130_fd_sc_hd__clkbuf_2
X_11205_ _07127_ _07190_ _07192_ net1444 VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__a2bb2o_1
X_12185_ net1343 _07749_ _07706_ CPU.mem_wdata\[4\] _07739_ VGND VGND VPWR VPWR _07752_
+ sky130_fd_sc_hd__a221o_1
X_18801_ net590 _02325_ VGND VGND VPWR VPWR CPU.aluReg\[31\] sky130_fd_sc_hd__dfxtp_1
X_11136_ _07134_ VGND VGND VPWR VPWR _07149_ sky130_fd_sc_hd__buf_2
X_16993_ _04688_ _04696_ _04542_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__o21a_1
X_13504__897 clknet_1_0__leaf__08435_ VGND VGND VPWR VPWR net953 sky130_fd_sc_hd__inv_2
X_18732_ net521 _02256_ VGND VGND VPWR VPWR mapped_spi_flash.snd_bitcount\[0\] sky130_fd_sc_hd__dfxtp_1
X_15944_ clknet_1_0__leaf__03686_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__buf_1
X_11067_ net1513 _07054_ _07101_ _07069_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__o211a_1
X_10018_ _05307_ _06346_ VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__or2_1
X_18663_ net452 _02187_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_14826_ _02798_ _02882_ _02886_ _02895_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__a31o_1
X_17614_ per_uart.d_in_uart\[6\] _05134_ _05157_ net1449 VGND VGND VPWR VPWR _05165_
+ sky130_fd_sc_hd__o22a_1
X_18594_ net415 net51 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14757_ _02827_ _02828_ _08783_ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17545_ _05112_ _05113_ _05058_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11969_ _06630_ net2448 _07609_ VGND VGND VPWR VPWR _07616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17476_ _05880_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__clkbuf_4
X_14688_ CPU.registerFile\[22\]\[9\] CPU.registerFile\[23\]\[9\] _08756_ VGND VGND
+ VPWR VPWR _02761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16427_ CPU.registerFile\[8\]\[10\] _04101_ _04102_ _04143_ VGND VGND VPWR VPWR _04144_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16358_ CPU.registerFile\[28\]\[8\] CPU.registerFile\[29\]\[8\] _03739_ VGND VGND
+ VPWR VPWR _04077_ sky130_fd_sc_hd__mux2_1
X_19146_ clknet_leaf_5_clk _02666_ VGND VGND VPWR VPWR per_uart.uart0.tx_count16\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15309_ _03049_ _03050_ CPU.registerFile\[25\]\[24\] VGND VGND VPWR VPWR _03367_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19077_ net69 _02597_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_16289_ _03692_ _03991_ _04009_ _03601_ VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__a211o_1
XFILLER_0_152_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18028_ net1039 _01556_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13661__1039 clknet_1_1__leaf__08450_ VGND VGND VPWR VPWR net1095 sky130_fd_sc_hd__inv_2
XFILLER_0_100_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15915__655 clknet_1_1__leaf__03687_ VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__inv_2
X_09801_ CPU.Jimm\[17\] _05550_ _05790_ CPU.cycles\[17\] _06138_ VGND VGND VPWR VPWR
+ _06139_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__03648_ _03648_ VGND VGND VPWR VPWR clknet_0__03648_ sky130_fd_sc_hd__clkbuf_16
X_13902__65 clknet_1_1__leaf__08475_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__inv_2
X_09732_ _05364_ _05747_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__nor2_1
X_09663_ _05916_ _06006_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09594_ CPU.Jimm\[13\] _05921_ _05923_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__a21o_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13336__834 clknet_1_0__leaf__08365_ VGND VGND VPWR VPWR net890 sky130_fd_sc_hd__inv_2
XFILLER_0_49_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15961__697 clknet_1_0__leaf__03691_ VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__inv_2
XFILLER_0_9_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17302__717 clknet_1_1__leaf__04980_ VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__inv_2
X_15660__458 clknet_1_0__leaf__03644_ VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__inv_2
XFILLER_0_33_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09028_ CPU.aluIn1\[21\] _05368_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold260 _01708_ VGND VGND VPWR VPWR net1557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 CPU.cycles\[6\] VGND VGND VPWR VPWR net1568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _02250_ VGND VGND VPWR VPWR net1579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 per_uart.uart0.enable16_counter\[5\] VGND VGND VPWR VPWR net1590 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12941_ _08172_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__clkbuf_1
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _06386_ net2102 _08131_ VGND VGND VPWR VPWR _08136_ sky130_fd_sc_hd__mux2_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _08764_ _08847_ _08849_ _08552_ VGND VGND VPWR VPWR _08850_ sky130_fd_sc_hd__a211o_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ net2464 _07335_ _07537_ VGND VGND VPWR VPWR _07539_ sky130_fd_sc_hd__mux2_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17402__25 clknet_1_0__leaf__05013_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__inv_2
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _08540_ VGND VGND VPWR VPWR _08783_ sky130_fd_sc_hd__buf_4
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14049__198 clknet_1_0__leaf__08489_ VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__inv_2
XFILLER_0_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _07502_ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__clkbuf_1
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17261_ CPU.registerFile\[0\]\[31\] _04637_ _03741_ _04956_ VGND VGND VPWR VPWR _04957_
+ sky130_fd_sc_hd__o211a_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ net1876 _06010_ _06816_ VGND VGND VPWR VPWR _06825_ sky130_fd_sc_hd__mux2_1
X_14473_ CPU.registerFile\[16\]\[4\] _08412_ _08714_ _06037_ VGND VGND VPWR VPWR _08715_
+ sky130_fd_sc_hd__o211a_1
X_11685_ _07465_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16212_ CPU.registerFile\[8\]\[5\] _08394_ _06150_ _03933_ VGND VGND VPWR VPWR _03934_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19000_ clknet_leaf_14_clk _02520_ VGND VGND VPWR VPWR CPU.aluIn1\[17\] sky130_fd_sc_hd__dfxtp_4
X_13424_ _08391_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__clkbuf_1
X_17192_ _03755_ _04877_ _04881_ _04889_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__a31o_1
X_10636_ CPU.registerFile\[1\]\[22\] _06032_ _06777_ VGND VGND VPWR VPWR _06787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16143_ CPU.registerFile\[2\]\[3\] CPU.registerFile\[3\]\[3\] _03693_ VGND VGND VPWR
+ VPWR _03867_ sky130_fd_sc_hd__mux2_1
X_10567_ _06749_ VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12306_ _07001_ net1322 _07829_ VGND VGND VPWR VPWR _07830_ sky130_fd_sc_hd__and3_1
X_16074_ CPU.registerFile\[27\]\[1\] CPU.registerFile\[26\]\[1\] _03745_ VGND VGND
+ VPWR VPWR _03800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10498_ _06712_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__clkbuf_1
X_15025_ CPU.registerFile\[24\]\[17\] _02928_ _03089_ _02771_ VGND VGND VPWR VPWR
+ _03090_ sky130_fd_sc_hd__o211a_1
X_12237_ net1435 _07785_ _07790_ _07755_ VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__o211a_1
X_15637__438 clknet_1_1__leaf__03641_ VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__inv_2
X_12168_ net1460 _07738_ _07741_ _07737_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__o211a_1
X_11119_ net1390 _07135_ VGND VGND VPWR VPWR _07140_ sky130_fd_sc_hd__or2_1
X_16976_ _04502_ _04667_ _04671_ _04679_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__a31o_2
X_12099_ _07692_ VGND VGND VPWR VPWR _07693_ sky130_fd_sc_hd__clkbuf_4
X_18715_ net504 _02239_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18646_ clknet_leaf_14_clk _02170_ VGND VGND VPWR VPWR CPU.rs2\[18\] sky130_fd_sc_hd__dfxtp_1
X_14809_ CPU.registerFile\[19\]\[12\] CPU.registerFile\[18\]\[12\] _02753_ VGND VGND
+ VPWR VPWR _02879_ sky130_fd_sc_hd__mux2_1
X_18577_ net398 net34 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_15789_ per_uart.uart0.enable16_counter\[2\] _08346_ VGND VGND VPWR VPWR _03662_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_148_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17528_ _05075_ _05025_ _06080_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_59_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17459_ _05022_ _06375_ _08256_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14260__388 clknet_1_1__leaf__08510_ VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__inv_2
XFILLER_0_116_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19129_ clknet_leaf_10_clk _02649_ VGND VGND VPWR VPWR CPU.PC\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__08486_ clknet_0__08486_ VGND VGND VPWR VPWR clknet_1_1__leaf__08486_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13833__1193 clknet_1_0__leaf__08468_ VGND VGND VPWR VPWR net1249 sky130_fd_sc_hd__inv_2
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09715_ _06056_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__clkbuf_1
X_09646_ _05988_ _05989_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__and2_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _05547_ CPU.instr\[4\] VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__or2_2
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11470_ _07342_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10421_ _06671_ VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13140_ CPU.cycles\[7\] _08275_ net1543 VGND VGND VPWR VPWR _08278_ sky130_fd_sc_hd__a21oi_1
X_10352_ _06144_ VGND VGND VPWR VPWR _06626_ sky130_fd_sc_hd__buf_4
XFILLER_0_104_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13071_ net1354 VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__clkbuf_1
X_10283_ net1750 _06316_ _06580_ VGND VGND VPWR VPWR _06582_ sky130_fd_sc_hd__mux2_1
X_12022_ _07644_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__clkbuf_1
X_16830_ _04175_ _04176_ CPU.registerFile\[17\]\[19\] VGND VGND VPWR VPWR _04538_
+ sky130_fd_sc_hd__a21o_1
X_16761_ _04468_ _04469_ _04153_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__mux2_1
X_18500_ net321 _02024_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_12924_ _08163_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__clkbuf_1
X_16692_ _04075_ _04398_ _04402_ _04042_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__o211a_1
X_18431_ net252 _01959_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ _06200_ net2410 _08120_ VGND VGND VPWR VPWR _08127_ sky130_fd_sc_hd__mux2_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13660__1038 clknet_1_1__leaf__08450_ VGND VGND VPWR VPWR net1094 sky130_fd_sc_hd__inv_2
X_11806_ net2153 _07318_ _07526_ VGND VGND VPWR VPWR _07530_ sky130_fd_sc_hd__mux2_1
X_13616__998 clknet_1_1__leaf__08446_ VGND VGND VPWR VPWR net1054 sky130_fd_sc_hd__inv_2
X_15574_ CPU.registerFile\[8\]\[31\] _08545_ _03624_ _08550_ VGND VGND VPWR VPWR _03625_
+ sky130_fd_sc_hd__o211a_1
X_18362_ net183 _01890_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _08089_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__clkbuf_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14525_ _08546_ _08547_ CPU.registerFile\[25\]\[5\] VGND VGND VPWR VPWR _08766_ sky130_fd_sc_hd__a21o_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_924 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _07493_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18293_ net114 _01821_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_14456_ CPU.registerFile\[8\]\[3\] _08526_ _08698_ _08622_ VGND VGND VPWR VPWR _08699_
+ sky130_fd_sc_hd__o211a_1
X_17244_ _03735_ _04936_ _04940_ _03732_ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__o211a_1
X_11668_ _07456_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13407_ _08382_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10619_ _06778_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__clkbuf_1
X_17175_ CPU.aluIn1\[28\] _08513_ _04873_ _04663_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14387_ CPU.registerFile\[0\]\[1\] _08584_ _08631_ _08588_ VGND VGND VPWR VPWR _08632_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11599_ _07419_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08440_ _08440_ VGND VGND VPWR VPWR clknet_0__08440_ sky130_fd_sc_hd__clkbuf_16
X_16126_ _03766_ _03846_ _03850_ _06142_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_1__f__08340_ clknet_0__08340_ VGND VGND VPWR VPWR clknet_1_1__leaf__08340_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_51_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16057_ CPU.registerFile\[15\]\[1\] CPU.registerFile\[14\]\[1\] _03705_ VGND VGND
+ VPWR VPWR _03783_ sky130_fd_sc_hd__mux2_1
X_13269_ net1590 _08349_ VGND VGND VPWR VPWR _08350_ sky130_fd_sc_hd__or2_1
X_13365__860 clknet_1_1__leaf__08368_ VGND VGND VPWR VPWR net916 sky130_fd_sc_hd__inv_2
X_15008_ net1646 _02797_ _03073_ _02993_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__o211a_1
X_17331__743 clknet_1_0__leaf__04983_ VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__inv_2
X_16959_ CPU.aluIn1\[22\] _04458_ _04662_ _04663_ VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09500_ _05388_ _05808_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09431_ _05255_ _05769_ _05770_ CPU.aluReg\[29\] _05780_ VGND VGND VPWR VPWR _05781_
+ sky130_fd_sc_hd__a221o_2
X_18629_ clknet_leaf_24_clk _02153_ VGND VGND VPWR VPWR CPU.mem_wdata\[1\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_59_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09362_ _05558_ _05712_ _05713_ _05235_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09293_ _05560_ _05629_ _05632_ _05630_ _05644_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__a311o_1
XANTENNA_11 _03637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_22 _04733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 _06171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 clknet_1_1__leaf__08340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_66 _06009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_77 _08549_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__08469_ clknet_0__08469_ VGND VGND VPWR VPWR clknet_1_1__leaf__08469_
+ sky130_fd_sc_hd__clkbuf_16
X_15772__559 clknet_1_1__leaf__03655_ VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__inv_2
XFILLER_0_98_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap13 _08330_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
X_10970_ net1515 _07007_ _07018_ _07014_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__o211a_1
X_09629_ _05945_ _05971_ _05972_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__a21o_1
X_18566__23 VGND VGND VPWR VPWR _18566__23/HI net23 sky130_fd_sc_hd__conb_1
XFILLER_0_66_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12640_ _06632_ net1922 _08004_ VGND VGND VPWR VPWR _08012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12571_ _07975_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__clkbuf_1
X_14243__372 clknet_1_0__leaf__08509_ VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__inv_2
XFILLER_0_148_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14310_ _08515_ _08519_ _08534_ _08555_ VGND VGND VPWR VPWR _08556_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11522_ _07377_ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__clkbuf_1
X_15290_ _03235_ _03236_ CPU.registerFile\[1\]\[23\] VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11453_ net2076 _07330_ _07312_ VGND VGND VPWR VPWR _07331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10404_ _06554_ VGND VGND VPWR VPWR _06661_ sky130_fd_sc_hd__clkbuf_4
X_11384_ _07289_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13123_ _08268_ _05538_ _05243_ _08266_ _06858_ VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__o311a_1
XFILLER_0_150_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10335_ _06614_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__clkbuf_1
X_18980_ net754 _02500_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ net1420 VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__clkbuf_1
X_17931_ net942 _01459_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_10266_ net1701 _06124_ _06569_ VGND VGND VPWR VPWR _06573_ sky130_fd_sc_hd__mux2_1
X_12005_ net2563 _07309_ _07635_ VGND VGND VPWR VPWR _07636_ sky130_fd_sc_hd__mux2_1
X_17862_ clknet_leaf_25_clk _00042_ VGND VGND VPWR VPWR CPU.cycles\[5\] sky130_fd_sc_hd__dfxtp_1
X_10197_ _05436_ _05274_ VGND VGND VPWR VPWR _06519_ sky130_fd_sc_hd__nand2_2
X_16813_ _06140_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__clkbuf_4
X_17793_ net873 _01355_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_16744_ _04367_ _04451_ _04453_ _04410_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__a211o_1
X_15749__539 clknet_1_1__leaf__03652_ VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__inv_2
X_12907_ _08154_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__clkbuf_1
X_16675_ CPU.registerFile\[5\]\[16\] CPU.registerFile\[4\]\[16\] _04024_ VGND VGND
+ VPWR VPWR _04386_ sky130_fd_sc_hd__mux2_1
X_13887_ clknet_1_1__leaf__08473_ VGND VGND VPWR VPWR _08474_ sky130_fd_sc_hd__buf_1
Xclkbuf_1_0__f__08489_ clknet_0__08489_ VGND VGND VPWR VPWR clknet_1_0__leaf__08489_
+ sky130_fd_sc_hd__clkbuf_16
X_18414_ net235 _01942_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12838_ _06010_ net2042 _08109_ VGND VGND VPWR VPWR _08118_ sky130_fd_sc_hd__mux2_1
X_13832__1192 clknet_1_0__leaf__08468_ VGND VGND VPWR VPWR net1248 sky130_fd_sc_hd__inv_2
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18345_ net166 _01873_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _08080_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15557_ CPU.registerFile\[21\]\[31\] _02752_ VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__04983_ clknet_0__04983_ VGND VGND VPWR VPWR clknet_1_1__leaf__04983_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14508_ _08425_ _08731_ _08749_ _08597_ VGND VGND VPWR VPWR _08750_ sky130_fd_sc_hd__a211o_1
X_15488_ _03539_ _03540_ _03255_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__mux2_1
X_18276_ net1287 _01804_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17227_ _03757_ _04919_ _04923_ _06109_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14439_ CPU.registerFile\[30\]\[3\] CPU.registerFile\[31\]\[3\] _08645_ VGND VGND
+ VPWR VPWR _08682_ sky130_fd_sc_hd__mux2_1
X_13929__90 clknet_1_1__leaf__08477_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__inv_2
XFILLER_0_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17158_ CPU.registerFile\[28\]\[28\] CPU.registerFile\[29\]\[28\] _04526_ VGND VGND
+ VPWR VPWR _04857_ sky130_fd_sc_hd__mux2_1
Xhold804 CPU.registerFile\[17\]\[23\] VGND VGND VPWR VPWR net2101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 CPU.registerFile\[26\]\[21\] VGND VGND VPWR VPWR net2112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold826 CPU.registerFile\[30\]\[15\] VGND VGND VPWR VPWR net2123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 CPU.registerFile\[21\]\[8\] VGND VGND VPWR VPWR net2134 sky130_fd_sc_hd__dlygate4sd3_1
X_16109_ CPU.registerFile\[30\]\[2\] CPU.registerFile\[31\]\[2\] _03796_ VGND VGND
+ VPWR VPWR _03834_ sky130_fd_sc_hd__mux2_1
Xhold848 CPU.registerFile\[29\]\[11\] VGND VGND VPWR VPWR net2145 sky130_fd_sc_hd__dlygate4sd3_1
X_17089_ _04484_ _04485_ CPU.registerFile\[25\]\[26\] VGND VGND VPWR VPWR _04790_
+ sky130_fd_sc_hd__a21o_1
X_09980_ mapped_spi_ram.rcv_data\[18\] _05761_ _05698_ net1351 VGND VGND VPWR VPWR
+ _06311_ sky130_fd_sc_hd__a22o_1
Xhold859 CPU.registerFile\[20\]\[14\] VGND VGND VPWR VPWR net2156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08931_ _05271_ _05281_ _05282_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09414_ _05556_ _05763_ _05764_ VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09345_ _05692_ _05694_ _05696_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09276_ _05561_ _05564_ _05627_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15854__601 clknet_1_0__leaf__03680_ VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__inv_2
XFILLER_0_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10120_ _05794_ _06444_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__or2_1
X_10051_ _05517_ _06372_ _06376_ _06378_ VGND VGND VPWR VPWR _06379_ sky130_fd_sc_hd__a31o_1
X_13952__111 clknet_1_0__leaf__08479_ VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__inv_2
XFILLER_0_100_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14790_ _02859_ _02860_ _08695_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10953_ _06992_ _07005_ VGND VGND VPWR VPWR _07006_ sky130_fd_sc_hd__and2_1
Xclkbuf_1_0__f__08343_ clknet_0__08343_ VGND VGND VPWR VPWR clknet_1_0__leaf__08343_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16460_ _04175_ _04176_ CPU.registerFile\[17\]\[10\] VGND VGND VPWR VPWR _04177_
+ sky130_fd_sc_hd__a21o_1
X_10884_ CPU.aluIn1\[6\] _06952_ _06880_ VGND VGND VPWR VPWR _06953_ sky130_fd_sc_hd__mux2_1
X_12623_ _06615_ net1763 _07993_ VGND VGND VPWR VPWR _08003_ sky130_fd_sc_hd__mux2_1
X_15411_ CPU.registerFile\[21\]\[27\] _02752_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16391_ CPU.registerFile\[12\]\[9\] _04017_ _04018_ _04108_ VGND VGND VPWR VPWR _04109_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_23_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_16
X_18130_ net1141 _01658_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_15342_ CPU.registerFile\[30\]\[25\] CPU.registerFile\[31\]\[25\] _03291_ VGND VGND
+ VPWR VPWR _03399_ sky130_fd_sc_hd__mux2_1
X_12554_ _07966_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11505_ _06439_ VGND VGND VPWR VPWR _07366_ sky130_fd_sc_hd__clkbuf_4
X_18061_ net1072 _01589_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_15273_ _03049_ _03050_ CPU.registerFile\[25\]\[23\] VGND VGND VPWR VPWR _03332_
+ sky130_fd_sc_hd__a21o_1
X_12485_ _07929_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17012_ _04502_ _04702_ _04706_ _04714_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__a31o_2
XFILLER_0_80_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11436_ _07319_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__03650_ clknet_0__03650_ VGND VGND VPWR VPWR clknet_1_1__leaf__03650_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14094__239 clknet_1_0__leaf__08493_ VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__inv_2
Xclkbuf_0__03681_ _03681_ VGND VGND VPWR VPWR clknet_0__03681_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11367_ _07280_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13106_ _06974_ net1488 mapped_spi_flash.state\[3\] VGND VGND VPWR VPWR _08259_ sky130_fd_sc_hd__o21a_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ _05804_ VGND VGND VPWR VPWR _06603_ sky130_fd_sc_hd__buf_2
X_18963_ net737 _02483_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_14086_ clknet_1_0__leaf__08484_ VGND VGND VPWR VPWR _08493_ sky130_fd_sc_hd__buf_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ net2473 _05839_ _07238_ VGND VGND VPWR VPWR _07244_ sky130_fd_sc_hd__mux2_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ net1443 VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__clkbuf_1
X_17914_ clknet_leaf_14_clk _01442_ VGND VGND VPWR VPWR CPU.Iimm\[1\] sky130_fd_sc_hd__dfxtp_2
X_10249_ net1792 _05839_ _06558_ VGND VGND VPWR VPWR _06564_ sky130_fd_sc_hd__mux2_1
X_18894_ net668 _02414_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17845_ net925 _01407_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_17776_ net856 _01338_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14988_ _02964_ _03047_ _03053_ _08851_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__o211a_1
X_16727_ _04098_ _04418_ _04425_ _04436_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__a31o_2
XFILLER_0_49_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16658_ CPU.registerFile\[16\]\[15\] _04252_ _04090_ _04369_ VGND VGND VPWR VPWR
+ _04370_ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16589_ CPU.registerFile\[13\]\[14\] _03976_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_14_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_16
X_09130_ _05353_ CPU.aluIn1\[18\] VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18328_ net149 _01856_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13330__829 clknet_1_1__leaf__08364_ VGND VGND VPWR VPWR net885 sky130_fd_sc_hd__inv_2
XFILLER_0_161_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09061_ _05253_ _05412_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__or2_2
X_18259_ net1270 _01787_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold601 CPU.registerFile\[5\]\[3\] VGND VGND VPWR VPWR net1898 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold612 CPU.registerFile\[2\]\[30\] VGND VGND VPWR VPWR net1909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold623 CPU.registerFile\[30\]\[14\] VGND VGND VPWR VPWR net1920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 CPU.registerFile\[9\]\[1\] VGND VGND VPWR VPWR net1931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 CPU.registerFile\[3\]\[13\] VGND VGND VPWR VPWR net1942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold656 CPU.registerFile\[22\]\[26\] VGND VGND VPWR VPWR net1953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 per_uart.rx_data\[5\] VGND VGND VPWR VPWR net1964 sky130_fd_sc_hd__dlygate4sd3_1
X_15695__490 clknet_1_1__leaf__03647_ VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__inv_2
Xhold678 CPU.registerFile\[15\]\[4\] VGND VGND VPWR VPWR net1975 sky130_fd_sc_hd__dlygate4sd3_1
X_09963_ _06294_ VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__clkbuf_1
Xhold689 CPU.registerFile\[7\]\[9\] VGND VGND VPWR VPWR net1986 sky130_fd_sc_hd__dlygate4sd3_1
X_08914_ CPU.aluIn1\[8\] _05262_ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__nor2_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _05425_ _06227_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__or2_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1301 CPU.registerFile\[25\]\[1\] VGND VGND VPWR VPWR net2598 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1312 CPU.registerFile\[8\]\[21\] VGND VGND VPWR VPWR net2609 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1323 CPU.registerFile\[12\]\[13\] VGND VGND VPWR VPWR net2620 sky130_fd_sc_hd__dlygate4sd3_1
X_13852__1211 clknet_1_1__leaf__08469_ VGND VGND VPWR VPWR net1267 sky130_fd_sc_hd__inv_2
Xhold1334 per_uart.uart0.rxd_reg\[8\] VGND VGND VPWR VPWR net2631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1345 CPU.PC\[20\] VGND VGND VPWR VPWR net2642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1356 CPU.aluReg\[16\] VGND VGND VPWR VPWR net2653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1367 mapped_spi_flash.rcv_data\[0\] VGND VGND VPWR VPWR net2664 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13532__922 clknet_1_0__leaf__08438_ VGND VGND VPWR VPWR net978 sky130_fd_sc_hd__inv_2
XFILLER_0_48_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09328_ _05677_ _05663_ VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09259_ CPU.aluIn1\[15\] CPU.Bimm\[12\] VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__xor2_1
XFILLER_0_161_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12270_ _07163_ VGND VGND VPWR VPWR _07809_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_160_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13908__71 clknet_1_0__leaf__08475_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__inv_2
X_11221_ _06599_ net2086 _07201_ VGND VGND VPWR VPWR _07203_ sky130_fd_sc_hd__mux2_1
X_11152_ mapped_spi_flash.rcv_data\[13\] _07149_ VGND VGND VPWR VPWR _07158_ sky130_fd_sc_hd__or2_1
X_10103_ _05269_ _05283_ _05291_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__o21ai_1
X_11083_ mapped_spi_flash.state\[1\] _07111_ net16 mapped_spi_flash.state\[2\] VGND
+ VGND VPWR VPWR _07113_ sky130_fd_sc_hd__a31o_1
X_14911_ CPU.registerFile\[8\]\[14\] _08776_ _02978_ _02864_ VGND VGND VPWR VPWR _02979_
+ sky130_fd_sc_hd__o211a_1
X_10034_ _06362_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__clkbuf_1
X_17630_ net1959 per_uart.uart0.rxd_reg\[5\] _05170_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__mux2_1
X_14842_ _08785_ _02909_ _02911_ _08870_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__a211o_1
X_17561_ _05127_ VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__clkbuf_1
X_11985_ _07624_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__clkbuf_1
X_14773_ _02751_ _02841_ _02843_ _02759_ VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__a211o_1
XFILLER_0_58_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16512_ CPU.registerFile\[12\]\[12\] _04017_ _04018_ _04226_ VGND VGND VPWR VPWR
+ _04227_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10936_ _06994_ VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__clkbuf_1
X_17492_ _05055_ _06237_ _05061_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__or3_1
XFILLER_0_156_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16443_ _04098_ _04145_ _04150_ _04159_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__a31o_2
XFILLER_0_67_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10867_ CPU.aluReg\[11\] CPU.aluReg\[9\] _06939_ VGND VGND VPWR VPWR _06940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12606_ _07994_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__clkbuf_1
X_19162_ clknet_leaf_27_clk _02682_ VGND VGND VPWR VPWR per_uart.rx_data\[1\] sky130_fd_sc_hd__dfxtp_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16374_ _03963_ _04089_ _04092_ _04006_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__a211o_1
XFILLER_0_143_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10798_ CPU.aluReg\[27\] CPU.aluReg\[25\] _06872_ VGND VGND VPWR VPWR _06887_ sky130_fd_sc_hd__mux2_1
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13774__1141 clknet_1_0__leaf__08461_ VGND VGND VPWR VPWR net1197 sky130_fd_sc_hd__inv_2
XFILLER_0_143_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18113_ net1124 _01641_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_12537_ net2544 _07309_ _07957_ VGND VGND VPWR VPWR _07958_ sky130_fd_sc_hd__mux2_1
X_15325_ CPU.registerFile\[2\]\[24\] CPU.registerFile\[3\]\[24\] _03275_ VGND VGND
+ VPWR VPWR _03383_ sky130_fd_sc_hd__mux2_1
X_19093_ net76 _02613_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_14102__246 clknet_1_0__leaf__08494_ VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__inv_2
X_18044_ net1055 _01572_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_12468_ net2346 _07309_ _07920_ VGND VGND VPWR VPWR _07921_ sky130_fd_sc_hd__mux2_1
X_15256_ _03027_ _03313_ _03315_ _03111_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13959__117 clknet_1_0__leaf__08480_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__inv_2
X_11419_ _07307_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__clkbuf_1
X_15187_ _03156_ _03245_ _03247_ _03163_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__a211o_1
X_12399_ _07883_ VGND VGND VPWR VPWR _07884_ sky130_fd_sc_hd__buf_4
XFILLER_0_111_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18946_ net720 _02466_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_3_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_146_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18877_ net651 _02397_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_17408__31 clknet_1_1__leaf__05013_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__inv_2
X_17828_ net908 _01390_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17759_ clknet_leaf_6_clk net1501 VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09113_ _05453_ _05464_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09044_ _05395_ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14077__223 clknet_1_1__leaf__08492_ VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__inv_2
XFILLER_0_103_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold420 CPU.registerFile\[5\]\[9\] VGND VGND VPWR VPWR net1717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold431 CPU.registerFile\[19\]\[6\] VGND VGND VPWR VPWR net1728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 CPU.registerFile\[6\]\[20\] VGND VGND VPWR VPWR net1739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 CPU.registerFile\[19\]\[10\] VGND VGND VPWR VPWR net1750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold464 CPU.registerFile\[5\]\[2\] VGND VGND VPWR VPWR net1761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 CPU.registerFile\[5\]\[10\] VGND VGND VPWR VPWR net1772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 CPU.registerFile\[28\]\[1\] VGND VGND VPWR VPWR net1783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold497 CPU.registerFile\[5\]\[18\] VGND VGND VPWR VPWR net1794 sky130_fd_sc_hd__dlygate4sd3_1
X_09946_ _06126_ _06277_ VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1120 CPU.registerFile\[8\]\[2\] VGND VGND VPWR VPWR net2417 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _05334_ _06187_ VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__xnor2_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 CPU.registerFile\[12\]\[0\] VGND VGND VPWR VPWR net2428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1142 CPU.registerFile\[8\]\[18\] VGND VGND VPWR VPWR net2439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 CPU.registerFile\[7\]\[6\] VGND VGND VPWR VPWR net2450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1164 CPU.registerFile\[8\]\[29\] VGND VGND VPWR VPWR net2461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1175 CPU.registerFile\[23\]\[0\] VGND VGND VPWR VPWR net2472 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1186 CPU.registerFile\[26\]\[0\] VGND VGND VPWR VPWR net2483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1197 CPU.registerFile\[22\]\[5\] VGND VGND VPWR VPWR net2494 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03653_ clknet_0__03653_ VGND VGND VPWR VPWR clknet_1_0__leaf__03653_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _07510_ VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__clkbuf_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _06833_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__clkbuf_1
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13440_ _06495_ VGND VGND VPWR VPWR _08403_ sky130_fd_sc_hd__clkbuf_8
X_10652_ _06795_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__clkbuf_1
X_13313__813 clknet_1_0__leaf__08363_ VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__inv_2
XFILLER_0_119_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10583_ net1924 _06224_ _06750_ VGND VGND VPWR VPWR _06758_ sky130_fd_sc_hd__mux2_1
X_12322_ _07780_ VGND VGND VPWR VPWR _07842_ sky130_fd_sc_hd__inv_2
X_15110_ CPU.registerFile\[27\]\[19\] CPU.registerFile\[26\]\[19\] _03172_ VGND VGND
+ VPWR VPWR _03173_ sky130_fd_sc_hd__mux2_1
X_16090_ CPU.aluIn1\[1\] _03566_ _03815_ _03390_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15041_ CPU.registerFile\[5\]\[17\] CPU.registerFile\[4\]\[17\] _03105_ VGND VGND
+ VPWR VPWR _03106_ sky130_fd_sc_hd__mux2_1
X_12253_ _07784_ VGND VGND VPWR VPWR _07799_ sky130_fd_sc_hd__buf_2
X_17350__11 clknet_1_0__leaf__04984_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__inv_2
XFILLER_0_32_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11204_ mapped_spi_flash.state\[3\] _07126_ _07188_ VGND VGND VPWR VPWR _07192_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12184_ net1360 _07738_ _07751_ _07737_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__o211a_1
X_18800_ net589 _02324_ VGND VGND VPWR VPWR CPU.aluReg\[30\] sky130_fd_sc_hd__dfxtp_1
X_11135_ net1593 _07147_ _07148_ _07138_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16992_ _04574_ _04691_ _04695_ _04584_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__o211a_1
X_18731_ net520 _02255_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[31\] sky130_fd_sc_hd__dfxtp_1
X_11066_ _07048_ _07100_ VGND VGND VPWR VPWR _07101_ sky130_fd_sc_hd__or2_1
X_15832__581 clknet_1_1__leaf__03678_ VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__inv_2
X_10017_ _05267_ _05306_ VGND VGND VPWR VPWR _06346_ sky130_fd_sc_hd__and2_1
X_18662_ net451 _02186_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17613_ net1510 _05159_ _05164_ _07108_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__o22a_1
X_14825_ _08722_ _02890_ _02894_ _08851_ VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__o211a_1
X_18593_ net414 net50 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_17544_ _08310_ _05895_ net13 VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__or3_1
X_14756_ CPU.registerFile\[5\]\[10\] CPU.registerFile\[4\]\[10\] _08864_ VGND VGND
+ VPWR VPWR _02828_ sky130_fd_sc_hd__mux2_1
X_11968_ _07615_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10919_ mapped_spi_flash.state\[1\] _06974_ _06975_ _06980_ VGND VGND VPWR VPWR _06981_
+ sky130_fd_sc_hd__a211oi_4
X_17475_ _05054_ _05056_ _05020_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11899_ _06628_ net2138 _07573_ VGND VGND VPWR VPWR _07579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14687_ _02751_ _02754_ _02758_ _02759_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__a211o_1
X_16426_ CPU.registerFile\[9\]\[10\] _04056_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14026__177 clknet_1_0__leaf__08487_ VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__inv_2
X_19145_ clknet_leaf_4_clk _02665_ VGND VGND VPWR VPWR per_uart.uart0.tx_count16\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16357_ CPU.registerFile\[30\]\[8\] CPU.registerFile\[31\]\[8\] _03796_ VGND VGND
+ VPWR VPWR _04076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13851__1210 clknet_1_1__leaf__08469_ VGND VGND VPWR VPWR net1266 sky130_fd_sc_hd__inv_2
XFILLER_0_70_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15308_ CPU.registerFile\[27\]\[24\] CPU.registerFile\[26\]\[24\] _03172_ VGND VGND
+ VPWR VPWR _03366_ sky130_fd_sc_hd__mux2_1
X_19076_ net68 _02596_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_16288_ _03999_ _04008_ _08406_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__o21a_1
XFILLER_0_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18027_ net1038 _01555_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15239_ _02964_ _03294_ _03298_ _03092_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13899__62 clknet_1_1__leaf__08475_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__inv_2
X_09800_ _05910_ _06135_ _06137_ _05881_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__o22ai_2
Xclkbuf_0__03647_ _03647_ VGND VGND VPWR VPWR clknet_0__03647_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15614__417 clknet_1_0__leaf__03639_ VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__inv_2
X_09731_ _06017_ _06068_ _06071_ _05516_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__o211a_1
X_18929_ net703 _02449_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_09662_ _05918_ _06004_ _06005_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__a21oi_1
X_09593_ _05935_ _05936_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09027_ _05378_ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold250 CPU.cycles\[23\] VGND VGND VPWR VPWR net1547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold261 mapped_spi_ram.rcv_data\[19\] VGND VGND VPWR VPWR net1558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 CPU.cycles\[2\] VGND VGND VPWR VPWR net1569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 CPU.rs2\[24\] VGND VGND VPWR VPWR net1580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 mapped_spi_flash.rcv_data\[26\] VGND VGND VPWR VPWR net1591 sky130_fd_sc_hd__dlygate4sd3_1
X_09929_ _05978_ _05941_ VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__or2b_1
X_13773__1140 clknet_1_0__leaf__08461_ VGND VGND VPWR VPWR net1196 sky130_fd_sc_hd__inv_2
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12940_ _06386_ net2400 _08167_ VGND VGND VPWR VPWR _08172_ sky130_fd_sc_hd__mux2_1
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _08135_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__clkbuf_1
X_17399__22 clknet_1_0__leaf__05013_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__inv_2
X_13988__143 clknet_1_0__leaf__08483_ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__inv_2
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ CPU.registerFile\[24\]\[7\] _08686_ _08848_ _08550_ VGND VGND VPWR VPWR _08849_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _07538_ VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__clkbuf_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14541_ CPU.registerFile\[5\]\[5\] CPU.registerFile\[4\]\[5\] _08576_ VGND VGND VPWR
+ VPWR _08782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11753_ _06617_ net2329 _07501_ VGND VGND VPWR VPWR _07502_ sky130_fd_sc_hd__mux2_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _06824_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__clkbuf_1
X_17260_ _03748_ _03750_ CPU.registerFile\[1\]\[31\] VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__a21o_1
XFILLER_0_154_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11684_ net2609 _07332_ _07464_ VGND VGND VPWR VPWR _07465_ sky130_fd_sc_hd__mux2_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14472_ CPU.registerFile\[17\]\[4\] _06456_ VGND VGND VPWR VPWR _08714_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16211_ CPU.registerFile\[9\]\[5\] _03698_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__or2_1
X_10635_ _06786_ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__clkbuf_1
X_13423_ _05856_ _06240_ _08388_ VGND VGND VPWR VPWR _08391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17191_ _03757_ _04884_ _04888_ _06109_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16142_ _03864_ _03865_ _03720_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__mux2_1
X_10566_ net2532 _06032_ _06739_ VGND VGND VPWR VPWR _06749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12305_ _07687_ _05238_ net1321 VGND VGND VPWR VPWR _07829_ sky130_fd_sc_hd__or3_1
X_16073_ _03797_ _03798_ _03742_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__mux2_1
X_10497_ net2117 _06032_ _06702_ VGND VGND VPWR VPWR _06712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12236_ mapped_spi_ram.rcv_data\[29\] _07787_ VGND VGND VPWR VPWR _07790_ sky130_fd_sc_hd__or2_1
X_15024_ _03049_ _03050_ CPU.registerFile\[25\]\[17\] VGND VGND VPWR VPWR _03089_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12167_ _07739_ _07740_ VGND VGND VPWR VPWR _07741_ sky130_fd_sc_hd__or2_1
X_13283__786 clknet_1_0__leaf__08345_ VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__inv_2
X_14214__347 clknet_1_0__leaf__08505_ VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__inv_2
X_11118_ net1390 _07133_ _07139_ _07138_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__o211a_1
X_16975_ _04305_ _04674_ _04678_ _04476_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__o211a_1
X_12098_ _07670_ net1312 _07688_ _07691_ VGND VGND VPWR VPWR _07692_ sky130_fd_sc_hd__o211a_2
X_18714_ net503 _02238_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[14\] sky130_fd_sc_hd__dfxtp_1
X_11049_ mapped_spi_flash.cmd_addr\[6\] _07086_ _07039_ VGND VGND VPWR VPWR _07087_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18645_ clknet_leaf_14_clk _02169_ VGND VGND VPWR VPWR CPU.rs2\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14808_ net1637 _02797_ _02878_ _08751_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__o211a_1
X_18576_ net397 net33 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_15788_ _08346_ _03657_ _03661_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17527_ _05069_ CPU.PC\[19\] _05098_ _05099_ _06858_ VGND VGND VPWR VPWR _02657_
+ sky130_fd_sc_hd__o221a_1
X_14739_ CPU.registerFile\[27\]\[10\] CPU.registerFile\[26\]\[10\] _02768_ VGND VGND
+ VPWR VPWR _02811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17458_ _06381_ _08336_ _05042_ _08334_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__o211a_1
X_16409_ CPU.registerFile\[24\]\[9\] _03915_ _03747_ _04126_ VGND VGND VPWR VPWR _04127_
+ sky130_fd_sc_hd__o211a_1
X_17389_ _04996_ _05011_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19128_ clknet_leaf_10_clk _02648_ VGND VGND VPWR VPWR CPU.PC\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19059_ net801 _02579_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08485_ clknet_0__08485_ VGND VGND VPWR VPWR clknet_1_1__leaf__08485_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_112_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15839__587 clknet_1_1__leaf__03679_ VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__inv_2
XFILLER_0_112_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14189__324 clknet_1_1__leaf__08503_ VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__inv_2
X_09714_ net2385 _06054_ _06055_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09645_ CPU.PC\[16\] _05987_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__or2_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ CPU.PC\[21\] _05919_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__or2_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13568__954 clknet_1_0__leaf__08442_ VGND VGND VPWR VPWR net1010 sky130_fd_sc_hd__inv_2
XFILLER_0_18_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10420_ _06607_ net2398 _06665_ VGND VGND VPWR VPWR _06671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10351_ _06625_ VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13070_ CPU.registerFile\[4\]\[10\] net1353 _08239_ VGND VGND VPWR VPWR _08241_ sky130_fd_sc_hd__mux2_1
X_10282_ _06581_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12021_ CPU.registerFile\[24\]\[23\] _07328_ _07635_ VGND VGND VPWR VPWR _07644_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16760_ CPU.registerFile\[5\]\[18\] CPU.registerFile\[4\]\[18\] _04428_ VGND VGND
+ VPWR VPWR _04469_ sky130_fd_sc_hd__mux2_1
X_13729__1100 clknet_1_1__leaf__08457_ VGND VGND VPWR VPWR net1156 sky130_fd_sc_hd__inv_2
X_13893__57 clknet_1_1__leaf__08474_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__inv_2
X_12923_ _06200_ net2253 _08156_ VGND VGND VPWR VPWR _08163_ sky130_fd_sc_hd__mux2_1
X_16691_ _04037_ _04399_ _04401_ _04208_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__a211o_2
X_18430_ net251 _01958_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _08126_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__clkbuf_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ net182 _01889_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_11805_ _07529_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__clkbuf_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _08546_ _08547_ CPU.registerFile\[9\]\[31\] VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _06641_ net2142 _08087_ VGND VGND VPWR VPWR _08089_ sky130_fd_sc_hd__mux2_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ CPU.registerFile\[27\]\[5\] CPU.registerFile\[26\]\[5\] _06063_ VGND VGND
+ VPWR VPWR _08765_ sky130_fd_sc_hd__mux2_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ _06601_ net1996 _07490_ VGND VGND VPWR VPWR _07493_ sky130_fd_sc_hd__mux2_1
X_18292_ net113 _01820_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15643__443 clknet_1_0__leaf__03642_ VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__inv_2
X_17243_ _08397_ _04937_ _04939_ _08400_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__a211o_1
XFILLER_0_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14455_ _08567_ _08569_ CPU.registerFile\[9\]\[3\] VGND VGND VPWR VPWR _08698_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11667_ net2461 _07316_ _07453_ VGND VGND VPWR VPWR _07456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13406_ _05422_ _06416_ _00000_ VGND VGND VPWR VPWR _08382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10618_ net2519 _05734_ _06777_ VGND VGND VPWR VPWR _06778_ sky130_fd_sc_hd__mux2_1
X_17174_ _04545_ _04855_ _04872_ _08596_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__a211o_2
X_11598_ net1890 _07316_ _07416_ VGND VGND VPWR VPWR _07419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14386_ _08585_ _08586_ CPU.registerFile\[1\]\[1\] VGND VGND VPWR VPWR _08631_ sky130_fd_sc_hd__a21o_1
X_16125_ CPU.registerFile\[16\]\[2\] _03848_ _03769_ _03849_ VGND VGND VPWR VPWR _03850_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10549_ _06740_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08370_ _08370_ VGND VGND VPWR VPWR clknet_0__08370_ sky130_fd_sc_hd__clkbuf_16
X_16056_ _08398_ _03779_ _03781_ _08401_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__a211o_1
XFILLER_0_110_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13268_ net1582 _08348_ VGND VGND VPWR VPWR _08349_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14138__278 clknet_1_1__leaf__08498_ VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__inv_2
X_15007_ _02750_ _03055_ _03072_ _02839_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__a211o_1
X_12219_ mapped_spi_ram.snd_bitcount\[0\] _07749_ _07764_ VGND VGND VPWR VPWR _07777_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13199_ _06548_ _06549_ _05440_ VGND VGND VPWR VPWR _08313_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_47_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16958_ _06855_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__clkbuf_4
X_16889_ _04419_ _04592_ _04594_ _04383_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__a211o_1
X_09430_ _05256_ _05771_ _05774_ _05779_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__a2bb2o_1
X_18628_ clknet_leaf_24_clk _02152_ VGND VGND VPWR VPWR CPU.mem_wdata\[0\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15726__518 clknet_1_1__leaf__03650_ VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__inv_2
X_09361_ CPU.PC\[2\] _05643_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__or2_1
X_18559_ net380 _02083_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09292_ CPU.aluIn1\[21\] _05544_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17393__17 clknet_1_1__leaf__04985_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__inv_2
XFILLER_0_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_12 _03833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_947 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_23 _04768_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_34 _06336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_45 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 clknet_1_1__leaf__08462_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 _06053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_78 _08569_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__08468_ clknet_0__08468_ VGND VGND VPWR VPWR clknet_1_1__leaf__08468_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__08499_ _08499_ VGND VGND VPWR VPWR clknet_0__08499_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09628_ CPU.PC\[9\] CPU.Bimm\[9\] _05914_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__and3_1
X_09559_ _05379_ _05902_ _05376_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_65_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12570_ net2608 _07345_ _07968_ VGND VGND VPWR VPWR _07975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18581__38 VGND VGND VPWR VPWR _18581__38/HI net38 sky130_fd_sc_hd__conb_1
X_11521_ net1691 _07376_ _07311_ VGND VGND VPWR VPWR _07377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11452_ _06031_ VGND VGND VPWR VPWR _07330_ sky130_fd_sc_hd__clkbuf_4
X_10403_ _06660_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11383_ net1710 _06124_ _07285_ VGND VGND VPWR VPWR _07289_ sky130_fd_sc_hd__mux2_1
X_13349__845 clknet_1_1__leaf__08367_ VGND VGND VPWR VPWR net901 sky130_fd_sc_hd__inv_2
XFILLER_0_132_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10334_ _06613_ net1936 _06597_ VGND VGND VPWR VPWR _06614_ sky130_fd_sc_hd__mux2_1
X_13122_ _05422_ VGND VGND VPWR VPWR _08268_ sky130_fd_sc_hd__inv_2
X_13053_ CPU.registerFile\[4\]\[18\] _06123_ _08228_ VGND VGND VPWR VPWR _08232_ sky130_fd_sc_hd__mux2_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17930_ net941 _01458_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_10265_ _06572_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__clkbuf_1
X_12004_ _07634_ VGND VGND VPWR VPWR _07635_ sky130_fd_sc_hd__clkbuf_4
X_17861_ clknet_leaf_1_clk _00041_ VGND VGND VPWR VPWR CPU.cycles\[4\] sky130_fd_sc_hd__dfxtp_1
X_10196_ CPU.PC\[1\] _06368_ _06382_ _06517_ VGND VGND VPWR VPWR _06518_ sky130_fd_sc_hd__a22o_1
X_16812_ CPU.registerFile\[0\]\[19\] _04233_ _04472_ _04519_ VGND VGND VPWR VPWR _04520_
+ sky130_fd_sc_hd__o211a_1
X_17792_ net872 _01354_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16743_ CPU.registerFile\[16\]\[17\] _04252_ _04090_ _04452_ VGND VGND VPWR VPWR
+ _04453_ sky130_fd_sc_hd__o211a_1
X_12906_ _06010_ net2416 _08145_ VGND VGND VPWR VPWR _08154_ sky130_fd_sc_hd__mux2_1
X_16674_ CPU.registerFile\[6\]\[16\] CPU.registerFile\[7\]\[16\] _04022_ VGND VGND
+ VPWR VPWR _04385_ sky130_fd_sc_hd__mux2_1
X_13886_ clknet_1_0__leaf__08339_ VGND VGND VPWR VPWR _08473_ sky130_fd_sc_hd__buf_1
X_18413_ net234 _01941_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[13\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__08488_ clknet_0__08488_ VGND VGND VPWR VPWR clknet_1_0__leaf__08488_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12837_ _08117_ VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__clkbuf_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18344_ net165 _01872_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15556_ CPU.registerFile\[22\]\[31\] CPU.registerFile\[23\]\[31\] _08584_ VGND VGND
+ VPWR VPWR _03607_ sky130_fd_sc_hd__mux2_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _06624_ net2254 _08076_ VGND VGND VPWR VPWR _08080_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__04982_ clknet_0__04982_ VGND VGND VPWR VPWR clknet_1_1__leaf__04982_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14507_ _08739_ _08748_ _08594_ VGND VGND VPWR VPWR _08749_ sky130_fd_sc_hd__o21a_1
X_11719_ net2503 _07368_ _07475_ VGND VGND VPWR VPWR _07483_ sky130_fd_sc_hd__mux2_1
X_18275_ net1286 _01803_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_15487_ CPU.registerFile\[28\]\[29\] CPU.registerFile\[29\]\[29\] _03212_ VGND VGND
+ VPWR VPWR _03540_ sky130_fd_sc_hd__mux2_1
X_12699_ _08043_ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17226_ _03765_ _04920_ _04922_ _06141_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__a211o_1
XFILLER_0_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14438_ _08521_ _08678_ _08680_ _08533_ VGND VGND VPWR VPWR _08681_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17157_ CPU.registerFile\[30\]\[28\] CPU.registerFile\[31\]\[28\] _04605_ VGND VGND
+ VPWR VPWR _04856_ sky130_fd_sc_hd__mux2_1
X_14369_ _08543_ _08611_ _08613_ _08552_ VGND VGND VPWR VPWR _08614_ sky130_fd_sc_hd__a211o_1
Xhold805 CPU.registerFile\[29\]\[7\] VGND VGND VPWR VPWR net2102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold816 CPU.registerFile\[3\]\[26\] VGND VGND VPWR VPWR net2113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16108_ _08404_ _03819_ _03823_ _03832_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__a31o_2
Xhold827 CPU.registerFile\[30\]\[7\] VGND VGND VPWR VPWR net2124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 CPU.registerFile\[3\]\[10\] VGND VGND VPWR VPWR net2135 sky130_fd_sc_hd__dlygate4sd3_1
X_17088_ CPU.registerFile\[27\]\[26\] CPU.registerFile\[26\]\[26\] _04646_ VGND VGND
+ VPWR VPWR _04789_ sky130_fd_sc_hd__mux2_1
Xhold849 CPU.registerFile\[18\]\[26\] VGND VGND VPWR VPWR net2146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16039_ _03765_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__clkbuf_8
X_08930_ CPU.aluIn1\[2\] _05270_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14071__218 clknet_1_1__leaf__08491_ VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__inv_2
XFILLER_0_0_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09413_ _05731_ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__buf_4
XFILLER_0_47_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09344_ _05577_ _05695_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_733 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09275_ CPU.aluIn1\[17\] CPU.aluIn1\[16\] _05544_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10050_ _05294_ _05532_ _05534_ CPU.aluReg\[7\] _06377_ VGND VGND VPWR VPWR _06378_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10952_ mapped_spi_flash.cmd_addr\[22\] _06983_ _06984_ mapped_spi_flash.cmd_addr\[21\]
+ VGND VGND VPWR VPWR _07005_ sky130_fd_sc_hd__a22o_1
Xclkbuf_1_0__f__08342_ clknet_0__08342_ VGND VGND VPWR VPWR clknet_1_0__leaf__08342_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15709__502 clknet_1_0__leaf__03649_ VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__inv_2
XFILLER_0_39_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10883_ CPU.aluReg\[7\] CPU.aluReg\[5\] _06939_ VGND VGND VPWR VPWR _06952_ sky130_fd_sc_hd__mux2_1
X_15410_ CPU.registerFile\[22\]\[27\] CPU.registerFile\[23\]\[27\] _08584_ VGND VGND
+ VPWR VPWR _03465_ sky130_fd_sc_hd__mux2_1
X_12622_ _08002_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__clkbuf_1
X_16390_ CPU.registerFile\[13\]\[9\] _03976_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15341_ _03078_ _03395_ _03397_ _03043_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__a211o_1
XFILLER_0_148_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12553_ net2522 _07328_ _07957_ VGND VGND VPWR VPWR _07966_ sky130_fd_sc_hd__mux2_1
X_18060_ net1071 _01588_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11504_ _07365_ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__clkbuf_1
X_15272_ CPU.registerFile\[27\]\[23\] CPU.registerFile\[26\]\[23\] _03172_ VGND VGND
+ VPWR VPWR _03331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12484_ net2087 _07328_ _07920_ VGND VGND VPWR VPWR _07929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17011_ _03757_ _04709_ _04713_ _04476_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11435_ net2061 _07318_ _07312_ VGND VGND VPWR VPWR _07319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__03680_ _03680_ VGND VGND VPWR VPWR clknet_0__03680_ sky130_fd_sc_hd__clkbuf_16
X_11366_ net1842 _05839_ _07274_ VGND VGND VPWR VPWR _07280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10317_ _06602_ VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__clkbuf_1
X_13105_ _07687_ _07779_ _07782_ _06858_ VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__o31ai_1
X_15755__544 clknet_1_0__leaf__03653_ VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__inv_2
X_18962_ net736 _02482_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11297_ _07243_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__clkbuf_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ CPU.registerFile\[4\]\[26\] _05838_ _08217_ VGND VGND VPWR VPWR _08223_ sky130_fd_sc_hd__mux2_1
X_10248_ _06563_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__clkbuf_1
X_17913_ clknet_leaf_17_clk _01441_ VGND VGND VPWR VPWR CPU.Iimm\[0\] sky130_fd_sc_hd__dfxtp_2
X_18893_ net667 _02413_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_17844_ net924 _01406_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_10179_ _06500_ _06501_ _05794_ VGND VGND VPWR VPWR _06502_ sky130_fd_sc_hd__o21ai_1
X_17775_ net855 _01337_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_14987_ _03006_ _03048_ _03052_ _02814_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__a211o_2
XFILLER_0_88_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16726_ _04305_ _04430_ _04435_ _04072_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16657_ _04175_ _04176_ CPU.registerFile\[17\]\[15\] VGND VGND VPWR VPWR _04369_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15608_ clknet_1_1__leaf__08506_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__buf_1
X_16588_ CPU.registerFile\[15\]\[14\] CPU.registerFile\[14\]\[14\] _04146_ VGND VGND
+ VPWR VPWR _04301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18327_ net148 _01855_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15539_ _08533_ _03586_ _03590_ _08554_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09060_ CPU.aluIn1\[30\] _05252_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__nor2_1
X_18258_ net1269 _01786_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17209_ _04898_ _04906_ _06474_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__o21a_1
X_18189_ net1200 net1432 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold602 CPU.registerFile\[30\]\[12\] VGND VGND VPWR VPWR net1899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 CPU.registerFile\[10\]\[6\] VGND VGND VPWR VPWR net1910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold624 CPU.registerFile\[13\]\[18\] VGND VGND VPWR VPWR net1921 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold635 CPU.registerFile\[10\]\[18\] VGND VGND VPWR VPWR net1932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 CPU.registerFile\[19\]\[11\] VGND VGND VPWR VPWR net1943 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 CPU.registerFile\[17\]\[26\] VGND VGND VPWR VPWR net1954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold668 _05176_ VGND VGND VPWR VPWR net1965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 CPU.registerFile\[20\]\[17\] VGND VGND VPWR VPWR net1976 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ net2363 _06292_ _06293_ VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08913_ CPU.aluIn1\[9\] _05264_ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__and2_2
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _06183_ _06226_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1302 CPU.aluShamt\[2\] VGND VGND VPWR VPWR net2599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1313 CPU.registerFile\[25\]\[28\] VGND VGND VPWR VPWR net2610 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1324 CPU.registerFile\[25\]\[0\] VGND VGND VPWR VPWR net2621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1335 _05178_ VGND VGND VPWR VPWR net2632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 CPU.aluReg\[30\] VGND VGND VPWR VPWR net2643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1357 CPU.aluIn1\[6\] VGND VGND VPWR VPWR net2654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1368 CPU.aluReg\[11\] VGND VGND VPWR VPWR net2665 sky130_fd_sc_hd__dlygate4sd3_1
X_15884__628 clknet_1_0__leaf__03683_ VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__inv_2
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13982__138 clknet_1_1__leaf__08482_ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__inv_2
XFILLER_0_153_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09327_ net1409 VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09258_ _05609_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15704__498 clknet_1_1__leaf__03648_ VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__inv_2
X_09189_ _05540_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__buf_4
XFILLER_0_105_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11220_ _07202_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11151_ net2612 _07147_ _07157_ _07151_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__o211a_1
X_14054__202 clknet_1_0__leaf__08490_ VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__inv_2
X_10102_ _05286_ _05431_ _05445_ _06427_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__a31o_1
X_11082_ mapped_spi_flash.snd_bitcount\[4\] mapped_spi_flash.snd_bitcount\[1\] mapped_spi_flash.snd_bitcount\[0\]
+ _06978_ VGND VGND VPWR VPWR _07112_ sky130_fd_sc_hd__nor4_1
X_14910_ _02733_ _02734_ CPU.registerFile\[9\]\[14\] VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__a21o_1
Xclkbuf_1_0__f__04985_ clknet_0__04985_ VGND VGND VPWR VPWR clknet_1_0__leaf__04985_
+ sky130_fd_sc_hd__clkbuf_16
X_10033_ net2425 _06361_ _06293_ VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__mux2_1
X_14841_ CPU.registerFile\[0\]\[12\] _08706_ _02910_ _02791_ VGND VGND VPWR VPWR _02911_
+ sky130_fd_sc_hd__o211a_1
X_17560_ net5 net1762 _06855_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__mux2_1
X_14772_ CPU.registerFile\[16\]\[11\] _02755_ _02842_ _02757_ VGND VGND VPWR VPWR
+ _02843_ sky130_fd_sc_hd__o211a_1
X_11984_ _06645_ net2243 _07620_ VGND VGND VPWR VPWR _07624_ sky130_fd_sc_hd__mux2_1
X_16511_ CPU.registerFile\[13\]\[12\] _03976_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17491_ _08379_ _05017_ _06235_ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__o21bai_1
X_10935_ _06992_ _06993_ VGND VGND VPWR VPWR _06994_ sky130_fd_sc_hd__and2_1
X_16442_ _03901_ _04154_ _04158_ _04072_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10866_ _06871_ VGND VGND VPWR VPWR _06939_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12605_ _06593_ net2036 _07993_ VGND VGND VPWR VPWR _07994_ sky130_fd_sc_hd__mux2_1
X_19161_ clknet_leaf_27_clk _02681_ VGND VGND VPWR VPWR per_uart.rx_data\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16373_ CPU.registerFile\[16\]\[8\] _03848_ _04090_ _04091_ VGND VGND VPWR VPWR _04092_
+ sky130_fd_sc_hd__o211a_1
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10797_ _06886_ VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18112_ net1123 _01640_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[22\] sky130_fd_sc_hd__dfxtp_1
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15324_ _03380_ _03381_ _03025_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__mux2_1
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12536_ _07956_ VGND VGND VPWR VPWR _07957_ sky130_fd_sc_hd__buf_4
X_19092_ net75 _02612_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_18043_ net1054 _01571_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_15255_ CPU.registerFile\[0\]\[22\] _02948_ _03314_ _03195_ VGND VGND VPWR VPWR _03315_
+ sky130_fd_sc_hd__o211a_1
X_12467_ _07919_ VGND VGND VPWR VPWR _07920_ sky130_fd_sc_hd__buf_4
XFILLER_0_151_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11418_ net1783 _06530_ _07273_ VGND VGND VPWR VPWR _07307_ sky130_fd_sc_hd__mux2_1
X_15679__475 clknet_1_0__leaf__03646_ VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__inv_2
X_15186_ CPU.registerFile\[16\]\[21\] _03159_ _03246_ _03161_ VGND VGND VPWR VPWR
+ _03247_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12398_ _07236_ _07451_ VGND VGND VPWR VPWR _07883_ sky130_fd_sc_hd__nor2_4
X_13789__1153 clknet_1_0__leaf__08464_ VGND VGND VPWR VPWR net1209 sky130_fd_sc_hd__inv_2
XFILLER_0_39_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11349_ _07270_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13247__768 clknet_1_1__leaf__08343_ VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__inv_2
X_18945_ net719 _02465_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_13019_ _08213_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__clkbuf_1
X_18876_ net650 _02396_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_17827_ net907 _01389_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_17758_ clknet_leaf_1_clk _00003_ VGND VGND VPWR VPWR CPU.state\[3\] sky130_fd_sc_hd__dfxtp_1
X_14183__319 clknet_1_1__leaf__08502_ VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__inv_2
XFILLER_0_77_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16709_ _03702_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__clkbuf_4
X_17689_ _05207_ _05216_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09112_ _05310_ _05462_ _05463_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09043_ _05393_ _05394_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__04979_ _04979_ VGND VGND VPWR VPWR clknet_0__04979_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_103_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14003__156 clknet_1_1__leaf__08485_ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__inv_2
XFILLER_0_25_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold410 CPU.PC\[3\] VGND VGND VPWR VPWR net1707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold421 CPU.registerFile\[10\]\[11\] VGND VGND VPWR VPWR net1718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13562__949 clknet_1_0__leaf__08441_ VGND VGND VPWR VPWR net1005 sky130_fd_sc_hd__inv_2
Xhold432 CPU.registerFile\[18\]\[25\] VGND VGND VPWR VPWR net1729 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 CPU.registerFile\[28\]\[25\] VGND VGND VPWR VPWR net1740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 CPU.registerFile\[5\]\[30\] VGND VGND VPWR VPWR net1751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold465 per_uart.uart_ctrl\[2\] VGND VGND VPWR VPWR net1762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 CPU.registerFile\[6\]\[25\] VGND VGND VPWR VPWR net1773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 CPU.registerFile\[20\]\[25\] VGND VGND VPWR VPWR net1784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold498 CPU.registerFile\[28\]\[13\] VGND VGND VPWR VPWR net1795 sky130_fd_sc_hd__dlygate4sd3_1
X_09945_ _05453_ _06276_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _05331_ _05533_ _05536_ CPU.aluReg\[14\] _06210_ VGND VGND VPWR VPWR _06211_
+ sky130_fd_sc_hd__a221o_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1110 CPU.registerFile\[21\]\[3\] VGND VGND VPWR VPWR net2407 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 CPU.registerFile\[17\]\[21\] VGND VGND VPWR VPWR net2418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1132 CPU.registerFile\[3\]\[4\] VGND VGND VPWR VPWR net2429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1143 CPU.registerFile\[23\]\[20\] VGND VGND VPWR VPWR net2440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 CPU.rs2\[31\] VGND VGND VPWR VPWR net2451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1165 CPU.registerFile\[29\]\[4\] VGND VGND VPWR VPWR net2462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 CPU.registerFile\[2\]\[26\] VGND VGND VPWR VPWR net2473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 CPU.registerFile\[14\]\[30\] VGND VGND VPWR VPWR net2484 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03652_ clknet_0__03652_ VGND VGND VPWR VPWR clknet_1_0__leaf__03652_
+ sky130_fd_sc_hd__clkbuf_16
Xhold1198 CPU.registerFile\[29\]\[17\] VGND VGND VPWR VPWR net2495 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ net2340 _06169_ _06827_ VGND VGND VPWR VPWR _06833_ sky130_fd_sc_hd__mux2_1
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10651_ net2559 _06200_ _06788_ VGND VGND VPWR VPWR _06795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10582_ _06757_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12321_ net1310 net1303 _07838_ _07841_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15040_ _06062_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__buf_4
X_12252_ net1516 _07785_ _07798_ _07796_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11203_ _07128_ _07190_ _07191_ net1446 VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__a2bb2o_1
X_12183_ net1355 _07749_ _07706_ CPU.mem_wdata\[5\] _07739_ VGND VGND VPWR VPWR _07751_
+ sky130_fd_sc_hd__a221o_1
X_11134_ net1602 _07135_ VGND VGND VPWR VPWR _07148_ sky130_fd_sc_hd__or2_1
X_16991_ _04367_ _04692_ _04694_ _04410_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__a211o_1
X_18730_ net519 _02254_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[30\] sky130_fd_sc_hd__dfxtp_1
X_11065_ mapped_spi_flash.cmd_addr\[3\] _05708_ _06976_ VGND VGND VPWR VPWR _07100_
+ sky130_fd_sc_hd__mux2_1
X_10016_ _06271_ _06344_ VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__and2_1
X_15867__612 clknet_1_0__leaf__03682_ VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__inv_2
X_13539__929 clknet_1_1__leaf__08438_ VGND VGND VPWR VPWR net985 sky130_fd_sc_hd__inv_2
X_18661_ net450 _02185_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_14824_ _08764_ _02891_ _02893_ _02814_ VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__a211o_2
X_17612_ per_uart.d_in_uart\[5\] _05134_ _05157_ net1478 VGND VGND VPWR VPWR _05164_
+ sky130_fd_sc_hd__o22a_1
X_18592_ net413 net49 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17543_ _05075_ _05025_ _06007_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__o21bai_1
X_14755_ CPU.registerFile\[6\]\[10\] CPU.registerFile\[7\]\[10\] _08740_ VGND VGND
+ VPWR VPWR _02827_ sky130_fd_sc_hd__mux2_1
X_11967_ _06628_ net2152 _07609_ VGND VGND VPWR VPWR _07615_ sky130_fd_sc_hd__mux2_1
X_13965__122 clknet_1_0__leaf__08481_ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__inv_2
X_10918_ _06976_ _06979_ VGND VGND VPWR VPWR _06980_ sky130_fd_sc_hd__nor2_2
X_17474_ _05055_ _06308_ _08331_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__or3_1
XFILLER_0_157_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14686_ _08419_ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__clkbuf_4
X_11898_ _07578_ VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__clkbuf_1
X_16425_ CPU.registerFile\[10\]\[10\] CPU.registerFile\[11\]\[10\] _03931_ VGND VGND
+ VPWR VPWR _04142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10849_ _06926_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19144_ clknet_leaf_4_clk _02664_ VGND VGND VPWR VPWR per_uart.tx_busy sky130_fd_sc_hd__dfxtp_2
X_16356_ _03713_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_109_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15307_ _03363_ _03364_ _03255_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__mux2_1
X_12519_ _07947_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19075_ net67 _02595_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_16287_ _03758_ _04002_ _04007_ _03775_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__o211a_1
X_18026_ net1037 _01554_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_15238_ _03006_ _03295_ _03297_ _03218_ VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__a211o_1
XFILLER_0_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15169_ CPU.registerFile\[6\]\[20\] CPU.registerFile\[7\]\[20\] _02982_ VGND VGND
+ VPWR VPWR _03231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0__03646_ _03646_ VGND VGND VPWR VPWR clknet_0__03646_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09730_ _06017_ _06070_ VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__nand2_1
X_18928_ net702 _02448_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_09661_ CPU.PC\[22\] _05917_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__and2_1
X_18859_ net633 _02379_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09592_ CPU.PC\[15\] _05934_ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13830__1191 clknet_1_0__leaf__08467_ VGND VGND VPWR VPWR net1247 sky130_fd_sc_hd__inv_2
XFILLER_0_18_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09026_ _05376_ _05377_ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold240 _01705_ VGND VGND VPWR VPWR net1537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 _08298_ VGND VGND VPWR VPWR net1548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 CPU.cycles\[9\] VGND VGND VPWR VPWR net1559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _08270_ VGND VGND VPWR VPWR net1570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 CPU.rs2\[27\] VGND VGND VPWR VPWR net1581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 mapped_spi_flash.rcv_data\[2\] VGND VGND VPWR VPWR net1592 sky130_fd_sc_hd__dlygate4sd3_1
X_09928_ _06257_ _06259_ _06260_ _05744_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__o31a_1
X_09859_ _05937_ _05986_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__xnor2_1
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14166__303 clknet_1_0__leaf__08501_ VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__inv_2
X_12870_ _06361_ net2397 _08131_ VGND VGND VPWR VPWR _08135_ sky130_fd_sc_hd__mux2_1
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ net2313 _07332_ _07537_ VGND VGND VPWR VPWR _07538_ sky130_fd_sc_hd__mux2_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ CPU.registerFile\[6\]\[5\] CPU.registerFile\[7\]\[5\] _08740_ VGND VGND VPWR
+ VPWR _08781_ sky130_fd_sc_hd__mux2_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13788__1152 clknet_1_0__leaf__08464_ VGND VGND VPWR VPWR net1208 sky130_fd_sc_hd__inv_2
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _07489_ VGND VGND VPWR VPWR _07501_ sky130_fd_sc_hd__buf_4
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ net1845 _05873_ _06816_ VGND VGND VPWR VPWR _06824_ sky130_fd_sc_hd__mux2_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14471_ CPU.registerFile\[19\]\[4\] CPU.registerFile\[18\]\[4\] _06064_ VGND VGND
+ VPWR VPWR _08713_ sky130_fd_sc_hd__mux2_1
X_11683_ _07452_ VGND VGND VPWR VPWR _07464_ sky130_fd_sc_hd__buf_4
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16210_ CPU.registerFile\[10\]\[5\] CPU.registerFile\[11\]\[5\] _03931_ VGND VGND
+ VPWR VPWR _03932_ sky130_fd_sc_hd__mux2_1
X_13422_ _08390_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10634_ net2648 _06010_ _06777_ VGND VGND VPWR VPWR _06786_ sky130_fd_sc_hd__mux2_1
X_17190_ _03765_ _04885_ _04887_ _06141_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16141_ CPU.registerFile\[5\]\[3\] CPU.registerFile\[4\]\[3\] _03704_ VGND VGND VPWR
+ VPWR _03865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10565_ _06748_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12304_ _05238_ net1321 _07687_ VGND VGND VPWR VPWR _07828_ sky130_fd_sc_hd__o21ai_1
X_16072_ CPU.registerFile\[28\]\[1\] CPU.registerFile\[29\]\[1\] _03739_ VGND VGND
+ VPWR VPWR _03798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10496_ _06711_ VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__clkbuf_1
X_15023_ CPU.registerFile\[27\]\[17\] CPU.registerFile\[26\]\[17\] _02768_ VGND VGND
+ VPWR VPWR _03088_ sky130_fd_sc_hd__mux2_1
X_12235_ net1437 _07785_ _07789_ _07755_ VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12166_ mapped_spi_ram.cmd_addr\[10\] _07097_ _07724_ VGND VGND VPWR VPWR _07740_
+ sky130_fd_sc_hd__mux2_1
X_11117_ net1366 _07135_ VGND VGND VPWR VPWR _07139_ sky130_fd_sc_hd__or2_1
X_16974_ _04347_ _04675_ _04677_ _04521_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__a211o_1
X_12097_ net1312 net14 VGND VGND VPWR VPWR _07691_ sky130_fd_sc_hd__nand2_1
X_18713_ net502 _02237_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[13\] sky130_fd_sc_hd__dfxtp_1
X_11048_ _07023_ _07084_ _07085_ _06853_ VGND VGND VPWR VPWR _07086_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18644_ clknet_leaf_15_clk _02168_ VGND VGND VPWR VPWR CPU.rs2\[16\] sky130_fd_sc_hd__dfxtp_1
X_14032__182 clknet_1_0__leaf__08488_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__inv_2
X_18587__44 VGND VGND VPWR VPWR _18587__44/HI net44 sky130_fd_sc_hd__conb_1
XFILLER_0_87_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14807_ _02750_ _02858_ _02877_ _02839_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__a211o_1
X_13869__1226 clknet_1_1__leaf__08471_ VGND VGND VPWR VPWR net1282 sky130_fd_sc_hd__inv_2
X_15787_ _03660_ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__buf_2
X_18575_ net396 net32 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_13591__975 clknet_1_1__leaf__08444_ VGND VGND VPWR VPWR net1031 sky130_fd_sc_hd__inv_2
X_12999_ _08180_ VGND VGND VPWR VPWR _08203_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17526_ _08335_ _06092_ _05073_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__o21ai_1
X_14738_ _02807_ _02809_ _08609_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17457_ _08310_ _06370_ _08330_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__or3_1
X_14669_ _08585_ _08586_ CPU.registerFile\[1\]\[8\] VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__a21o_1
XFILLER_0_157_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16408_ _04080_ _04081_ CPU.registerFile\[25\]\[9\] VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__a21o_1
X_15921__661 clknet_1_0__leaf__03687_ VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__inv_2
XFILLER_0_129_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17388_ per_uart.uart0.uart_rxd2 _04992_ _04993_ per_uart.uart0.rxd_reg\[9\] VGND
+ VGND VPWR VPWR _05011_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16339_ CPU.registerFile\[8\]\[8\] _08394_ _06150_ _04057_ VGND VGND VPWR VPWR _04058_
+ sky130_fd_sc_hd__o211a_1
X_19127_ clknet_leaf_10_clk _02647_ VGND VGND VPWR VPWR CPU.PC\[9\] sky130_fd_sc_hd__dfxtp_2
X_15620__422 clknet_1_1__leaf__03640_ VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__inv_2
XFILLER_0_42_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19058_ net800 _02578_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__08484_ clknet_0__08484_ VGND VGND VPWR VPWR clknet_1_1__leaf__08484_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13485__880 clknet_1_0__leaf__08370_ VGND VGND VPWR VPWR net936 sky130_fd_sc_hd__inv_2
XFILLER_0_11_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18009_ net1020 _01537_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13342__840 clknet_1_1__leaf__08365_ VGND VGND VPWR VPWR net896 sky130_fd_sc_hd__inv_2
X_14115__257 clknet_1_1__leaf__08496_ VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__inv_2
X_09713_ net15 VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__buf_4
X_09644_ CPU.PC\[16\] _05987_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09575_ CPU.Iimm\[1\] _05545_ _05914_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__mux2_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14161__299 clknet_1_1__leaf__08500_ VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__inv_2
XFILLER_0_150_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10350_ _06624_ net1818 _06618_ VGND VGND VPWR VPWR _06625_ sky130_fd_sc_hd__mux2_1
X_09009_ _05350_ _05360_ _05349_ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__o21ba_1
X_10281_ net1943 _06292_ _06580_ VGND VGND VPWR VPWR _06581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12020_ _07643_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__clkbuf_1
X_12922_ _08162_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__clkbuf_1
X_16690_ CPU.registerFile\[24\]\[16\] _04319_ _04165_ _04400_ VGND VGND VPWR VPWR
+ _04401_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15641_ clknet_1_0__leaf__08506_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__buf_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12853_ _06169_ net2324 _08120_ VGND VGND VPWR VPWR _08126_ sky130_fd_sc_hd__mux2_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ net2302 _07316_ _07526_ VGND VGND VPWR VPWR _07529_ sky130_fd_sc_hd__mux2_1
X_18360_ net181 _01888_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ CPU.registerFile\[10\]\[31\] CPU.registerFile\[11\]\[31\] _08522_ VGND VGND
+ VPWR VPWR _03623_ sky130_fd_sc_hd__mux2_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _08088_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _06418_ VGND VGND VPWR VPWR _08764_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_139_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _07492_ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__clkbuf_1
X_18291_ net112 _01819_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17242_ CPU.registerFile\[16\]\[30\] _04656_ _06149_ _04938_ VGND VGND VPWR VPWR
+ _04939_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14454_ CPU.registerFile\[10\]\[3\] CPU.registerFile\[11\]\[3\] _08564_ VGND VGND
+ VPWR VPWR _08697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11666_ _07455_ VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_924 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13405_ _08381_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__clkbuf_1
X_10617_ _06776_ VGND VGND VPWR VPWR _06777_ sky130_fd_sc_hd__buf_4
X_17173_ _04863_ _04871_ _04542_ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__o21a_1
XFILLER_0_153_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14385_ CPU.registerFile\[2\]\[1\] CPU.registerFile\[3\]\[1\] _08629_ VGND VGND VPWR
+ VPWR _08630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11597_ _07418_ VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__clkbuf_1
X_16124_ _03770_ _03771_ CPU.registerFile\[17\]\[2\] VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__a21o_1
X_10548_ net2163 _05734_ _06739_ VGND VGND VPWR VPWR _06740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16055_ CPU.registerFile\[8\]\[1\] _08394_ _06150_ _03780_ VGND VGND VPWR VPWR _03781_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13267_ per_uart.uart0.enable16_counter\[3\] _08347_ VGND VGND VPWR VPWR _08348_
+ sky130_fd_sc_hd__or2_1
X_10479_ net2088 _05734_ _06702_ VGND VGND VPWR VPWR _06703_ sky130_fd_sc_hd__mux2_1
X_15006_ _03063_ _03071_ _02837_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__o21a_2
X_12218_ mapped_spi_ram.snd_bitcount\[0\] _07704_ _07764_ VGND VGND VPWR VPWR _07776_
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_121_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13198_ _06043_ _06112_ _06185_ _06186_ VGND VGND VPWR VPWR _08312_ sky130_fd_sc_hd__or4_1
X_13708__1081 clknet_1_0__leaf__08455_ VGND VGND VPWR VPWR net1137 sky130_fd_sc_hd__inv_2
X_12149_ _07715_ _07727_ VGND VGND VPWR VPWR _07728_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16957_ _04545_ _04642_ _04661_ _04500_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__a211o_1
XFILLER_0_47_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16888_ CPU.registerFile\[12\]\[21\] _04421_ _04422_ _04593_ VGND VGND VPWR VPWR
+ _04594_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18627_ net448 _02151_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__05015_ _05015_ VGND VGND VPWR VPWR clknet_0__05015_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09360_ _05711_ _05581_ VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__xnor2_1
X_18558_ net379 _02082_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15845__592 clknet_1_0__leaf__03680_ VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__inv_2
X_17509_ _05055_ _06156_ _05061_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__or3_1
X_13372__866 clknet_1_1__leaf__08369_ VGND VGND VPWR VPWR net922 sky130_fd_sc_hd__inv_2
XFILLER_0_157_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09291_ _05636_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__buf_2
X_18489_ net310 _02013_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[21\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_13 _04033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_24 _04785_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 _07360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_46 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_57 clknet_1_1__leaf__08462_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 _06058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 clknet_1_1__leaf__08448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__08467_ clknet_0__08467_ VGND VGND VPWR VPWR clknet_1_1__leaf__08467_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_112_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_859 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08498_ _08498_ VGND VGND VPWR VPWR clknet_0__08498_ sky130_fd_sc_hd__clkbuf_16
X_15590__395 clknet_1_1__leaf__08511_ VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__inv_2
Xmax_cap15 _05741_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
X_09627_ _05946_ _05969_ _05970_ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__a21o_1
X_15928__667 clknet_1_0__leaf__03688_ VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__inv_2
X_09558_ _05367_ _05370_ _05380_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09489_ _05399_ _05533_ _05536_ net1441 _05835_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__a221o_2
X_11520_ _06554_ VGND VGND VPWR VPWR _07376_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11451_ _07329_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10402_ _06659_ net1980 _06596_ VGND VGND VPWR VPWR _06660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11382_ _07288_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13121_ _07108_ _08267_ VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10333_ _06009_ VGND VGND VPWR VPWR _06613_ sky130_fd_sc_hd__clkbuf_4
X_13868__1225 clknet_1_1__leaf__08471_ VGND VGND VPWR VPWR net1281 sky130_fd_sc_hd__inv_2
X_13052_ net1329 VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__clkbuf_1
X_10264_ net1877 _06106_ _06569_ VGND VGND VPWR VPWR _06572_ sky130_fd_sc_hd__mux2_1
X_12003_ _06813_ _07633_ VGND VGND VPWR VPWR _07634_ sky130_fd_sc_hd__nor2b_4
X_17315__729 clknet_1_1__leaf__04981_ VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__inv_2
X_17860_ clknet_leaf_25_clk _00040_ VGND VGND VPWR VPWR CPU.cycles\[3\] sky130_fd_sc_hd__dfxtp_1
X_10195_ _06488_ _06516_ VGND VGND VPWR VPWR _06517_ sky130_fd_sc_hd__and2_1
X_16811_ _04389_ _04390_ CPU.registerFile\[1\]\[19\] VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__a21o_1
X_17791_ net871 _01353_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_16742_ _04175_ _04176_ CPU.registerFile\[17\]\[17\] VGND VGND VPWR VPWR _04452_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12905_ _08153_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__clkbuf_1
X_16673_ _04015_ _04379_ _04382_ _04383_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_0__f__08487_ clknet_0__08487_ VGND VGND VPWR VPWR clknet_1_0__leaf__08487_
+ sky130_fd_sc_hd__clkbuf_16
X_18412_ net233 _01940_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_12836_ _05873_ net2206 _08109_ VGND VGND VPWR VPWR _08117_ sky130_fd_sc_hd__mux2_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18343_ net164 _01871_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_15555_ _08521_ _03603_ _03605_ _08590_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__a211o_1
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _08079_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__04981_ clknet_0__04981_ VGND VGND VPWR VPWR clknet_1_1__leaf__04981_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _08574_ _08743_ _08747_ _08592_ VGND VGND VPWR VPWR _08748_ sky130_fd_sc_hd__o211a_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11718_ _07482_ VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__clkbuf_1
X_18274_ net1285 _01802_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14144__283 clknet_1_0__leaf__08499_ VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__inv_2
X_15486_ CPU.registerFile\[30\]\[29\] CPU.registerFile\[31\]\[29\] _03291_ VGND VGND
+ VPWR VPWR _03539_ sky130_fd_sc_hd__mux2_1
X_12698_ _06622_ net2638 _08040_ VGND VGND VPWR VPWR _08043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17225_ CPU.registerFile\[0\]\[30\] _04637_ _03741_ _04921_ VGND VGND VPWR VPWR _04922_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14437_ CPU.registerFile\[20\]\[3\] _08527_ _08679_ _08530_ VGND VGND VPWR VPWR _08680_
+ sky130_fd_sc_hd__o211a_1
X_11649_ _07445_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17156_ _04502_ _04842_ _04846_ _04854_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__a31o_1
XFILLER_0_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14368_ CPU.registerFile\[24\]\[1\] _08545_ _08612_ _08550_ VGND VGND VPWR VPWR _08613_
+ sky130_fd_sc_hd__o211a_1
Xhold806 CPU.registerFile\[27\]\[8\] VGND VGND VPWR VPWR net2103 sky130_fd_sc_hd__dlygate4sd3_1
X_16107_ _03716_ _03826_ _03831_ _03732_ VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__o211a_1
Xhold817 CPU.registerFile\[31\]\[29\] VGND VGND VPWR VPWR net2114 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold828 CPU.registerFile\[22\]\[9\] VGND VGND VPWR VPWR net2125 sky130_fd_sc_hd__dlygate4sd3_1
X_17087_ _04786_ _04787_ _06535_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__mux2_1
Xhold839 CPU.registerFile\[31\]\[26\] VGND VGND VPWR VPWR net2136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14299_ _08410_ VGND VGND VPWR VPWR _08545_ sky130_fd_sc_hd__buf_4
X_16038_ _08396_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_15732__523 clknet_1_0__leaf__03651_ VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__inv_2
X_13597__981 clknet_1_0__leaf__08444_ VGND VGND VPWR VPWR net1037 sky130_fd_sc_hd__inv_2
X_17989_ net1000 _01517_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09412_ mapped_spi_ram.rcv_data\[6\] _05761_ _05762_ net1346 VGND VGND VPWR VPWR
+ _05763_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14227__358 clknet_1_0__leaf__08507_ VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__inv_2
X_09343_ CPU.aluIn1\[0\] _05576_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__or2_1
XFILLER_0_158_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09274_ _05617_ _05623_ _05624_ _05625_ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13935__95 clknet_1_1__leaf__08478_ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__inv_2
XFILLER_0_140_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08989_ CPU.aluIn1\[16\] _05339_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10951_ _07004_ VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__08341_ clknet_0__08341_ VGND VGND VPWR VPWR clknet_1_0__leaf__08341_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15861__607 clknet_1_1__leaf__03681_ VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__inv_2
X_19197__55 VGND VGND VPWR VPWR _19197__55/HI net55 sky130_fd_sc_hd__conb_1
X_10882_ _06951_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__clkbuf_1
X_12621_ _06613_ net1786 _07993_ VGND VGND VPWR VPWR _08002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_857 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15340_ CPU.registerFile\[20\]\[25\] _03080_ _03396_ _03082_ VGND VGND VPWR VPWR
+ _03397_ sky130_fd_sc_hd__o211a_1
X_13707__1080 clknet_1_0__leaf__08455_ VGND VGND VPWR VPWR net1136 sky130_fd_sc_hd__inv_2
X_12552_ _07965_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11503_ net1753 _07364_ _07354_ VGND VGND VPWR VPWR _07365_ sky130_fd_sc_hd__mux2_1
X_15271_ _03328_ _03329_ _03255_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__mux2_1
X_12483_ _07928_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__clkbuf_1
X_17010_ _04347_ _04710_ _04712_ _04521_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__a211o_1
XFILLER_0_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11434_ _05804_ VGND VGND VPWR VPWR _07318_ sky130_fd_sc_hd__buf_4
XFILLER_0_105_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14153_ clknet_1_1__leaf__08495_ VGND VGND VPWR VPWR _08500_ sky130_fd_sc_hd__buf_1
XFILLER_0_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11365_ _07279_ VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13104_ _07762_ _08258_ _05237_ VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__a21oi_1
X_10316_ _06601_ net1719 _06597_ VGND VGND VPWR VPWR _06602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18961_ net735 _02481_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_11296_ net2338 _05825_ _07238_ VGND VGND VPWR VPWR _07243_ sky130_fd_sc_hd__mux2_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ net1340 VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__clkbuf_1
X_17912_ clknet_leaf_17_clk _01440_ VGND VGND VPWR VPWR CPU.Jimm\[19\] sky130_fd_sc_hd__dfxtp_1
X_10247_ net1796 _05825_ _06558_ VGND VGND VPWR VPWR _06563_ sky130_fd_sc_hd__mux2_1
X_18892_ net666 _02412_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_17843_ net923 _01405_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_10178_ _05440_ _05435_ _05439_ VGND VGND VPWR VPWR _06501_ sky130_fd_sc_hd__and3_1
X_17774_ net854 _01336_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_14986_ CPU.registerFile\[24\]\[16\] _02928_ _03051_ _02771_ VGND VGND VPWR VPWR
+ _03052_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16725_ _04347_ _04432_ _04434_ _04117_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__a211o_1
XFILLER_0_135_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16656_ CPU.registerFile\[19\]\[15\] CPU.registerFile\[18\]\[15\] _04327_ VGND VGND
+ VPWR VPWR _04368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12819_ _05276_ _06861_ _06869_ _08107_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16587_ _04099_ _04297_ _04299_ _04105_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18326_ net147 _01854_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15538_ _08543_ _03587_ _03589_ _03307_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__a211o_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15469_ _03521_ _03522_ _08562_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__mux2_1
X_18257_ net1268 _01785_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17208_ _04574_ _04901_ _04905_ _04584_ VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18188_ net1199 net1430 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[27\] sky130_fd_sc_hd__dfxtp_1
Xhold603 CPU.registerFile\[6\]\[31\] VGND VGND VPWR VPWR net1900 sky130_fd_sc_hd__dlygate4sd3_1
X_15957__693 clknet_1_1__leaf__03691_ VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__inv_2
XFILLER_0_13_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold614 CPU.registerFile\[3\]\[7\] VGND VGND VPWR VPWR net1911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17139_ net2584 _04458_ _04838_ _04663_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__o211a_1
Xhold625 CPU.registerFile\[27\]\[14\] VGND VGND VPWR VPWR net1922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 CPU.registerFile\[2\]\[1\] VGND VGND VPWR VPWR net1933 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 CPU.registerFile\[15\]\[16\] VGND VGND VPWR VPWR net1944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 CPU.registerFile\[20\]\[8\] VGND VGND VPWR VPWR net1955 sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ net15 VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__buf_4
Xhold669 CPU.registerFile\[21\]\[16\] VGND VGND VPWR VPWR net1966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15656__454 clknet_1_1__leaf__03644_ VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__inv_2
X_08912_ CPU.rs2\[9\] CPU.Bimm\[9\] _05244_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _05457_ _06181_ _06182_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__and3b_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1303 CPU.registerFile\[12\]\[4\] VGND VGND VPWR VPWR net2600 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1314 CPU.registerFile\[1\]\[18\] VGND VGND VPWR VPWR net2611 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1325 per_uart.uart0.rx_count16\[0\] VGND VGND VPWR VPWR net2622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1336 CPU.aluReg\[4\] VGND VGND VPWR VPWR net2633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1347 CPU.registerFile\[25\]\[7\] VGND VGND VPWR VPWR net2644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1358 CPU.registerFile\[25\]\[10\] VGND VGND VPWR VPWR net2655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1369 CPU.cycles\[4\] VGND VGND VPWR VPWR net2666 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13867__1224 clknet_1_1__leaf__08471_ VGND VGND VPWR VPWR net1280 sky130_fd_sc_hd__inv_2
XFILLER_0_76_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09326_ _05663_ _05672_ _05677_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_118_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09257_ CPU.aluIn1\[13\] CPU.Bimm\[12\] VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__xor2_2
XFILLER_0_161_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09188_ _05538_ _05539_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__and2_2
XFILLER_0_121_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11150_ mapped_spi_flash.rcv_data\[14\] _07149_ VGND VGND VPWR VPWR _07157_ sky130_fd_sc_hd__or2_1
X_10101_ _05794_ _05446_ VGND VGND VPWR VPWR _06427_ sky130_fd_sc_hd__nand2_1
X_11081_ mapped_spi_flash.snd_bitcount\[5\] VGND VGND VPWR VPWR _07111_ sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__04984_ clknet_0__04984_ VGND VGND VPWR VPWR clknet_1_0__leaf__04984_
+ sky130_fd_sc_hd__clkbuf_16
X_10032_ _06360_ VGND VGND VPWR VPWR _06361_ sky130_fd_sc_hd__buf_4
X_14840_ _02831_ _02832_ CPU.registerFile\[1\]\[12\] VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__a21o_1
X_14771_ CPU.registerFile\[17\]\[11\] _08795_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__or2_1
X_11983_ _07623_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__clkbuf_1
X_16510_ CPU.registerFile\[15\]\[12\] CPU.registerFile\[14\]\[12\] _04146_ VGND VGND
+ VPWR VPWR _04225_ sky130_fd_sc_hd__mux2_1
X_10934_ mapped_spi_flash.cmd_addr\[28\] _06983_ _06985_ mapped_spi_flash.cmd_addr\[27\]
+ VGND VGND VPWR VPWR _06993_ sky130_fd_sc_hd__a22o_1
X_17490_ _08255_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13653_ clknet_1_0__leaf__08440_ VGND VGND VPWR VPWR _08450_ sky130_fd_sc_hd__buf_1
X_16441_ _03943_ _04155_ _04157_ _04117_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__a211o_1
X_10865_ _06938_ VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12604_ _07992_ VGND VGND VPWR VPWR _07993_ sky130_fd_sc_hd__buf_4
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19160_ clknet_leaf_4_clk net1450 VGND VGND VPWR VPWR per_uart.uart0.txd_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16372_ _03770_ _03771_ CPU.registerFile\[17\]\[8\] VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__a21o_1
X_10796_ CPU.aluReg\[27\] _06885_ _06869_ VGND VGND VPWR VPWR _06886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15323_ CPU.registerFile\[5\]\[24\] CPU.registerFile\[4\]\[24\] _03105_ VGND VGND
+ VPWR VPWR _03381_ sky130_fd_sc_hd__mux2_1
X_18111_ net1122 _01639_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12535_ _07955_ _06813_ VGND VGND VPWR VPWR _07956_ sky130_fd_sc_hd__nor2_4
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19091_ net74 _02611_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18042_ net1053 _01570_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_15254_ _03235_ _03236_ CPU.registerFile\[1\]\[22\] VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12466_ _07414_ _07451_ VGND VGND VPWR VPWR _07919_ sky130_fd_sc_hd__nor2_4
XFILLER_0_2_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11417_ _07306_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__clkbuf_1
X_15185_ CPU.registerFile\[17\]\[21\] _03036_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__or2_1
X_12397_ _07882_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14256__384 clknet_1_1__leaf__08510_ VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__inv_2
X_11348_ net2460 _06508_ _07260_ VGND VGND VPWR VPWR _07270_ sky130_fd_sc_hd__mux2_1
X_13914__76 clknet_1_0__leaf__08476_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__inv_2
X_18944_ net718 _02464_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_11279_ _06657_ net2554 _07223_ VGND VGND VPWR VPWR _07233_ sky130_fd_sc_hd__mux2_1
X_13018_ net2614 _07372_ _08203_ VGND VGND VPWR VPWR _08213_ sky130_fd_sc_hd__mux2_1
X_18875_ net649 _02395_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_17826_ net906 _01388_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17757_ clknet_leaf_1_clk _00002_ VGND VGND VPWR VPWR CPU.state\[2\] sky130_fd_sc_hd__dfxtp_1
X_14969_ CPU.registerFile\[19\]\[16\] CPU.registerFile\[18\]\[16\] _02753_ VGND VGND
+ VPWR VPWR _03035_ sky130_fd_sc_hd__mux2_1
X_13516__908 clknet_1_1__leaf__08436_ VGND VGND VPWR VPWR net964 sky130_fd_sc_hd__inv_2
X_16708_ _04099_ _04415_ _04417_ _04105_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17688_ CPU.mem_wdata\[3\] per_uart.uart0.tx_wr _05211_ VGND VGND VPWR VPWR _05216_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16639_ _04347_ _04348_ _04350_ _04117_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__a211o_1
XFILLER_0_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09111_ _05260_ CPU.aluIn1\[10\] VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__or2b_1
XFILLER_0_162_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18309_ net130 _01837_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09042_ CPU.aluIn1\[27\] _05392_ VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13673__1049 clknet_1_0__leaf__08452_ VGND VGND VPWR VPWR net1105 sky130_fd_sc_hd__inv_2
XFILLER_0_13_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold400 CPU.registerFile\[19\]\[31\] VGND VGND VPWR VPWR net1697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 CPU.registerFile\[6\]\[29\] VGND VGND VPWR VPWR net1708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 CPU.registerFile\[15\]\[29\] VGND VGND VPWR VPWR net1719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15890__633 clknet_1_1__leaf__03684_ VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__inv_2
Xhold433 CPU.registerFile\[28\]\[5\] VGND VGND VPWR VPWR net1730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 CPU.registerFile\[11\]\[18\] VGND VGND VPWR VPWR net1741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 CPU.registerFile\[2\]\[25\] VGND VGND VPWR VPWR net1752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 CPU.registerFile\[27\]\[22\] VGND VGND VPWR VPWR net1763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 CPU.registerFile\[31\]\[10\] VGND VGND VPWR VPWR net1774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 CPU.registerFile\[28\]\[10\] VGND VGND VPWR VPWR net1785 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ _05261_ _05311_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__nor2_1
Xhold499 CPU.registerFile\[19\]\[27\] VGND VGND VPWR VPWR net1796 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _05332_ _05749_ VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__nor2_1
Xhold1100 CPU.registerFile\[29\]\[8\] VGND VGND VPWR VPWR net2397 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 CPU.registerFile\[21\]\[23\] VGND VGND VPWR VPWR net2408 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 CPU.registerFile\[12\]\[19\] VGND VGND VPWR VPWR net2419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 CPU.registerFile\[23\]\[12\] VGND VGND VPWR VPWR net2430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 CPU.registerFile\[14\]\[0\] VGND VGND VPWR VPWR net2441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 CPU.registerFile\[20\]\[9\] VGND VGND VPWR VPWR net2452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1166 CPU.registerFile\[20\]\[5\] VGND VGND VPWR VPWR net2463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1177 CPU.registerFile\[17\]\[10\] VGND VGND VPWR VPWR net2474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1188 CPU.registerFile\[31\]\[22\] VGND VGND VPWR VPWR net2485 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03651_ clknet_0__03651_ VGND VGND VPWR VPWR clknet_1_0__leaf__03651_
+ sky130_fd_sc_hd__clkbuf_16
Xhold1199 CPU.registerFile\[1\]\[17\] VGND VGND VPWR VPWR net2496 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414__36 clknet_1_1__leaf__05014_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__inv_2
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10650_ _06794_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__clkbuf_1
X_17717__48 clknet_1_0__leaf__05015_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__inv_2
XFILLER_0_75_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09309_ _05566_ _05660_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10581_ net2044 _06200_ _06750_ VGND VGND VPWR VPWR _06757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12320_ _07781_ _07840_ VGND VGND VPWR VPWR _07841_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12251_ mapped_spi_ram.rcv_data\[22\] _07787_ VGND VGND VPWR VPWR _07798_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11202_ mapped_spi_flash.state\[3\] _07127_ _07188_ VGND VGND VPWR VPWR _07191_ sky130_fd_sc_hd__a21o_1
X_12182_ net1349 _07738_ _07750_ _07737_ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__o211a_1
X_11133_ _07132_ VGND VGND VPWR VPWR _07147_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16990_ CPU.registerFile\[16\]\[23\] _04656_ _04494_ _04693_ VGND VGND VPWR VPWR
+ _04694_ sky130_fd_sc_hd__o211a_1
X_11064_ net1521 _07054_ _07099_ _07069_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__o211a_1
X_10015_ _05267_ _05428_ _05448_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__nand3b_1
X_18660_ net449 _02184_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17611_ net1476 _05159_ _05163_ _07108_ VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__o22a_1
X_14823_ CPU.registerFile\[24\]\[12\] _08686_ _02892_ _02771_ VGND VGND VPWR VPWR
+ _02893_ sky130_fd_sc_hd__o211a_1
X_18591_ net412 net48 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17542_ _05069_ net2650 _05110_ _05111_ _06858_ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__o221a_1
X_14754_ _08532_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__clkbuf_4
X_11966_ _07614_ VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10917_ net1555 net1588 _06977_ _06978_ VGND VGND VPWR VPWR _06979_ sky130_fd_sc_hd__or4_1
X_17473_ _08310_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__clkbuf_2
X_14685_ CPU.registerFile\[16\]\[9\] _02755_ _02756_ _02757_ VGND VGND VPWR VPWR _02758_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11897_ _06626_ net2316 _07573_ VGND VGND VPWR VPWR _07578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16424_ _06085_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__clkbuf_4
X_10848_ net2670 _06925_ _06922_ VGND VGND VPWR VPWR _06926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19143_ clknet_leaf_0_clk _02663_ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_143_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16355_ _08404_ _04059_ _04063_ _04073_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__a31o_4
X_13253__773 clknet_1_0__leaf__08344_ VGND VGND VPWR VPWR net829 sky130_fd_sc_hd__inv_2
X_10779_ _06871_ VGND VGND VPWR VPWR _06872_ sky130_fd_sc_hd__buf_4
XFILLER_0_27_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12518_ net2435 _07362_ _07942_ VGND VGND VPWR VPWR _07947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15306_ CPU.registerFile\[28\]\[24\] CPU.registerFile\[29\]\[24\] _03212_ VGND VGND
+ VPWR VPWR _03364_ sky130_fd_sc_hd__mux2_1
X_19074_ net66 _02594_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16286_ _03963_ _04003_ _04005_ _04006_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13498_ clknet_1_0__leaf__08366_ VGND VGND VPWR VPWR _08435_ sky130_fd_sc_hd__buf_1
X_18025_ net1036 _01553_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_12449_ _07910_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__clkbuf_1
X_15237_ CPU.registerFile\[24\]\[22\] _02928_ _03296_ _03175_ VGND VGND VPWR VPWR
+ _03297_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15168_ _08532_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__buf_2
X_13866__1223 clknet_1_1__leaf__08471_ VGND VGND VPWR VPWR net1279 sky130_fd_sc_hd__inv_2
Xclkbuf_0__03645_ _03645_ VGND VGND VPWR VPWR clknet_0__03645_ sky130_fd_sc_hd__clkbuf_16
X_15099_ CPU.registerFile\[16\]\[19\] _03159_ _03160_ _03161_ VGND VGND VPWR VPWR
+ _03162_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18927_ net701 _02447_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_09660_ _05920_ _06002_ _06003_ VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__a21o_1
X_18858_ net632 _02378_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_17809_ net889 _01371_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_09591_ CPU.PC\[15\] _05934_ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__and2_1
X_18789_ net578 _02313_ VGND VGND VPWR VPWR CPU.aluReg\[19\] sky130_fd_sc_hd__dfxtp_1
X_15768__555 clknet_1_0__leaf__03655_ VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__inv_2
XFILLER_0_82_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09025_ CPU.aluIn1\[22\] _05375_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold230 _02368_ VGND VGND VPWR VPWR net1527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold241 CPU.cycles\[17\] VGND VGND VPWR VPWR net1538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold252 CPU.cycles\[29\] VGND VGND VPWR VPWR net1549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 CPU.cycles\[20\] VGND VGND VPWR VPWR net1560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 CPU.cycles\[15\] VGND VGND VPWR VPWR net1571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 per_uart.uart0.enable16_counter\[4\] VGND VGND VPWR VPWR net1582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 mapped_spi_flash.rcv_data\[20\] VGND VGND VPWR VPWR net1593 sky130_fd_sc_hd__dlygate4sd3_1
X_09927_ _05319_ _05523_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__nor2_1
X_09858_ _06191_ _06193_ _05541_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__o21a_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _05340_ _05344_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__nor2_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _07525_ VGND VGND VPWR VPWR _07537_ sky130_fd_sc_hd__buf_4
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _07500_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__clkbuf_1
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _06823_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__clkbuf_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ CPU.mem_wdata\[3\] _08514_ _08712_ _07822_ VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11682_ _07463_ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__clkbuf_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _05526_ _06247_ _08388_ VGND VGND VPWR VPWR _08390_ sky130_fd_sc_hd__mux2_1
X_10633_ _06785_ VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16140_ CPU.registerFile\[6\]\[3\] CPU.registerFile\[7\]\[3\] _03717_ VGND VGND VPWR
+ VPWR _03864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10564_ net2003 _06010_ _06739_ VGND VGND VPWR VPWR _06748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12303_ mapped_spi_ram.div_counter\[1\] net1320 VGND VGND VPWR VPWR _07827_ sky130_fd_sc_hd__xnor2_1
X_16071_ CPU.registerFile\[30\]\[1\] CPU.registerFile\[31\]\[1\] _03796_ VGND VGND
+ VPWR VPWR _03797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13545__934 clknet_1_0__leaf__08439_ VGND VGND VPWR VPWR net990 sky130_fd_sc_hd__inv_2
X_10495_ net2101 _06010_ _06702_ VGND VGND VPWR VPWR _06711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15022_ _03085_ _03086_ _02851_ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12234_ net1427 _07787_ VGND VGND VPWR VPWR _07789_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12165_ _07695_ VGND VGND VPWR VPWR _07739_ sky130_fd_sc_hd__buf_2
XFILLER_0_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11116_ net1366 _07133_ _07137_ _07138_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__o211a_1
X_12096_ mapped_spi_ram.snd_bitcount\[3\] mapped_spi_ram.snd_bitcount\[2\] mapped_spi_ram.snd_bitcount\[1\]
+ _07689_ VGND VGND VPWR VPWR _07690_ sky130_fd_sc_hd__nor4_1
X_16973_ CPU.registerFile\[0\]\[23\] _04637_ _04472_ _04676_ VGND VGND VPWR VPWR _04677_
+ sky130_fd_sc_hd__o211a_1
X_18712_ net501 _02236_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[12\] sky130_fd_sc_hd__dfxtp_1
X_11047_ CPU.PC\[7\] _05643_ VGND VGND VPWR VPWR _07085_ sky130_fd_sc_hd__or2_1
X_18643_ clknet_leaf_14_clk _02167_ VGND VGND VPWR VPWR CPU.rs2\[15\] sky130_fd_sc_hd__dfxtp_1
X_15855_ clknet_1_1__leaf__03654_ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__buf_1
X_14806_ _02867_ _02876_ _02837_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__o21a_2
X_13672__1048 clknet_1_0__leaf__08452_ VGND VGND VPWR VPWR net1104 sky130_fd_sc_hd__inv_2
X_18574_ net395 net31 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_15786_ _06854_ _03659_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__nand2_1
X_12998_ _08202_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17525_ _05096_ _05097_ _05058_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14737_ CPU.registerFile\[28\]\[10\] CPU.registerFile\[29\]\[10\] _02808_ VGND VGND
+ VPWR VPWR _02809_ sky130_fd_sc_hd__mux2_1
X_11949_ _07605_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__clkbuf_1
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17456_ _05016_ net2603 _05040_ _05041_ _07002_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__o221a_1
XFILLER_0_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14668_ CPU.registerFile\[2\]\[8\] CPU.registerFile\[3\]\[8\] _08629_ VGND VGND VPWR
+ VPWR _02742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16407_ CPU.registerFile\[27\]\[9\] CPU.registerFile\[26\]\[9\] _03837_ VGND VGND
+ VPWR VPWR _04125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17387_ _05010_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__clkbuf_1
X_14599_ CPU.registerFile\[22\]\[7\] CPU.registerFile\[23\]\[7\] _08756_ VGND VGND
+ VPWR VPWR _08838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19126_ clknet_leaf_2_clk _02646_ VGND VGND VPWR VPWR CPU.PC\[8\] sky130_fd_sc_hd__dfxtp_1
X_16338_ CPU.registerFile\[9\]\[8\] _04056_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19057_ net799 _02577_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_16269_ _03901_ _03983_ _03989_ _03732_ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_1__f__08483_ clknet_0__08483_ VGND VGND VPWR VPWR clknet_1_1__leaf__08483_
+ sky130_fd_sc_hd__clkbuf_16
X_18008_ net1019 _01536_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09712_ _06053_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__buf_4
X_09643_ CPU.Jimm\[16\] _05921_ _05923_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__a21o_1
X_09574_ CPU.PC\[22\] _05917_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__or2_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15595__400 clknet_1_1__leaf__08511_ VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__inv_2
XFILLER_0_103_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09008_ CPU.aluIn1\[18\] _05353_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10280_ _06557_ VGND VGND VPWR VPWR _06580_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12921_ _06169_ net2513 _08156_ VGND VGND VPWR VPWR _08162_ sky130_fd_sc_hd__mux2_1
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _08125_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__clkbuf_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _07528_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _03620_ _03621_ _08541_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__mux2_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _06638_ net2078 _08087_ VGND VGND VPWR VPWR _08088_ sky130_fd_sc_hd__mux2_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11734_ _06599_ net2011 _07490_ VGND VGND VPWR VPWR _07492_ sky130_fd_sc_hd__mux2_1
X_14522_ _08761_ _08762_ _08609_ VGND VGND VPWR VPWR _08763_ sky130_fd_sc_hd__mux2_1
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13865__1222 clknet_1_1__leaf__08471_ VGND VGND VPWR VPWR net1278 sky130_fd_sc_hd__inv_2
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18290_ net111 _01818_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _03749_ _03751_ CPU.registerFile\[17\]\[30\] VGND VGND VPWR VPWR _04938_
+ sky130_fd_sc_hd__a21o_1
X_14453_ _08692_ _08694_ _08695_ VGND VGND VPWR VPWR _08696_ sky130_fd_sc_hd__mux2_1
X_11665_ net2183 _07314_ _07453_ VGND VGND VPWR VPWR _07455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10616_ _06774_ _06775_ VGND VGND VPWR VPWR _06776_ sky130_fd_sc_hd__nor2_2
X_13404_ _05538_ _06461_ _00000_ VGND VGND VPWR VPWR _08381_ sky130_fd_sc_hd__mux2_1
X_14384_ _08525_ VGND VGND VPWR VPWR _08629_ sky130_fd_sc_hd__buf_4
X_17172_ _04574_ _04866_ _04870_ _04584_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__o211a_1
X_11596_ net2528 _07314_ _07416_ VGND VGND VPWR VPWR _07418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16123_ _03847_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__clkbuf_4
X_10547_ _06738_ VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__buf_4
XFILLER_0_107_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13266_ per_uart.uart0.enable16_counter\[2\] _08346_ VGND VGND VPWR VPWR _08347_
+ sky130_fd_sc_hd__or2_1
X_16054_ CPU.registerFile\[9\]\[1\] _03698_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__or2_1
X_10478_ _06701_ VGND VGND VPWR VPWR _06702_ sky130_fd_sc_hd__buf_4
XFILLER_0_121_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15005_ _02826_ _03066_ _03070_ _02746_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__o211a_1
X_12217_ mapped_spi_ram.snd_bitcount\[2\] _07764_ _07775_ _07694_ VGND VGND VPWR VPWR
+ _01723_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13197_ _08310_ VGND VGND VPWR VPWR _08311_ sky130_fd_sc_hd__buf_2
X_13326__825 clknet_1_0__leaf__08364_ VGND VGND VPWR VPWR net881 sky130_fd_sc_hd__inv_2
XFILLER_0_20_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15951__688 clknet_1_1__leaf__03690_ VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__inv_2
X_12148_ mapped_spi_ram.cmd_addr\[15\] _07066_ _07724_ VGND VGND VPWR VPWR _07727_
+ sky130_fd_sc_hd__mux2_1
X_12079_ _07670_ _07671_ _07677_ mapped_spi_ram.rbusy VGND VGND VPWR VPWR _07678_
+ sky130_fd_sc_hd__a22o_1
X_16956_ _04651_ _04660_ _04542_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__o21a_1
X_16887_ CPU.registerFile\[13\]\[21\] _04380_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__or2_1
X_18626_ net447 _02150_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__05014_ _05014_ VGND VGND VPWR VPWR clknet_0__05014_ sky130_fd_sc_hd__clkbuf_16
X_18557_ net378 _02081_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_17508_ _05075_ _05025_ _06153_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__o21bai_1
X_09290_ _05638_ _05641_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18488_ net309 _02012_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_14 _04074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17439_ _08334_ _06477_ _08255_ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__o21a_1
XANTENNA_25 _04803_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_36 _07452_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_47 clknet_1_0__leaf__03656_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 clknet_1_1__leaf__08451_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_69 _06105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14121__262 clknet_1_1__leaf__08497_ VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__inv_2
XFILLER_0_42_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19109_ net92 _02629_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14195__330 clknet_1_0__leaf__08503_ VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__inv_2
XFILLER_0_3_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08466_ clknet_0__08466_ VGND VGND VPWR VPWR clknet_1_1__leaf__08466_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__08497_ _08497_ VGND VGND VPWR VPWR clknet_0__08497_ sky130_fd_sc_hd__clkbuf_16
X_14039__189 clknet_1_1__leaf__08488_ VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__inv_2
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap16 _07112_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
X_13574__960 clknet_1_1__leaf__08442_ VGND VGND VPWR VPWR net1016 sky130_fd_sc_hd__inv_2
X_09626_ CPU.PC\[8\] CPU.Bimm\[8\] _05914_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09557_ _05374_ _05900_ VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__xnor2_1
X_15627__429 clknet_1_0__leaf__03640_ VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__inv_2
X_09488_ _05398_ _05829_ _05834_ _05516_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_66_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17344__5 clknet_1_0__leaf__04984_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__inv_2
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11450_ net1686 _07328_ _07312_ VGND VGND VPWR VPWR _07329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10401_ _06529_ VGND VGND VPWR VPWR _06659_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_116_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11381_ net1738 _06106_ _07285_ VGND VGND VPWR VPWR _07288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13120_ _08255_ _06176_ _08266_ CPU.state\[2\] VGND VGND VPWR VPWR _08267_ sky130_fd_sc_hd__o2bb2a_1
X_10332_ _06612_ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13671__1047 clknet_1_0__leaf__08452_ VGND VGND VPWR VPWR net1103 sky130_fd_sc_hd__inv_2
X_13051_ CPU.registerFile\[4\]\[19\] net1328 _08228_ VGND VGND VPWR VPWR _08231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10263_ _06571_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__clkbuf_1
X_12002_ _05738_ _05737_ _05739_ VGND VGND VPWR VPWR _07633_ sky130_fd_sc_hd__and3b_4
X_10194_ CPU.PC\[1\] _05952_ VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__or2_1
X_16810_ CPU.registerFile\[2\]\[19\] CPU.registerFile\[3\]\[19\] _04431_ VGND VGND
+ VPWR VPWR _04518_ sky130_fd_sc_hd__mux2_1
X_14250__379 clknet_1_1__leaf__08509_ VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__inv_2
X_17790_ net870 _01352_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16741_ CPU.registerFile\[19\]\[17\] CPU.registerFile\[18\]\[17\] _04327_ VGND VGND
+ VPWR VPWR _04451_ sky130_fd_sc_hd__mux2_1
X_13953_ clknet_1_0__leaf__08473_ VGND VGND VPWR VPWR _08480_ sky130_fd_sc_hd__buf_1
X_12904_ _05873_ net1658 _08145_ VGND VGND VPWR VPWR _08153_ sky130_fd_sc_hd__mux2_1
X_16672_ _03713_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__buf_4
X_18411_ net232 _01939_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[11\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__08486_ clknet_0__08486_ VGND VGND VPWR VPWR clknet_1_0__leaf__08486_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _08116_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__clkbuf_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ net163 _01870_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ CPU.registerFile\[16\]\[31\] _08527_ _03604_ _08530_ VGND VGND VPWR VPWR
+ _03605_ sky130_fd_sc_hd__o211a_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__04980_ clknet_0__04980_ VGND VGND VPWR VPWR clknet_1_1__leaf__04980_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _06622_ net2281 _08076_ VGND VGND VPWR VPWR _08079_ sky130_fd_sc_hd__mux2_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18572__29 VGND VGND VPWR VPWR _18572__29/HI net29 sky130_fd_sc_hd__conb_1
X_14505_ _08581_ _08744_ _08746_ _08590_ VGND VGND VPWR VPWR _08747_ sky130_fd_sc_hd__a211o_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ net2560 _07366_ _07475_ VGND VGND VPWR VPWR _07482_ sky130_fd_sc_hd__mux2_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ net1284 _01801_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_12697_ _08042_ VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__clkbuf_1
X_15485_ _08581_ _03535_ _03537_ _08535_ VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__a211o_1
X_17224_ _03748_ _03750_ CPU.registerFile\[1\]\[30\] VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__a21o_1
X_11648_ net2534 _07366_ _07438_ VGND VGND VPWR VPWR _07445_ sky130_fd_sc_hd__mux2_1
X_14436_ CPU.registerFile\[21\]\[3\] _08528_ VGND VGND VPWR VPWR _08679_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17155_ _03757_ _04849_ _04853_ _06109_ VGND VGND VPWR VPWR _04854_ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11579_ net2240 _07366_ _07401_ VGND VGND VPWR VPWR _07408_ sky130_fd_sc_hd__mux2_1
X_14367_ _08546_ _08547_ CPU.registerFile\[25\]\[1\] VGND VGND VPWR VPWR _08612_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold807 CPU.registerFile\[29\]\[0\] VGND VGND VPWR VPWR net2104 sky130_fd_sc_hd__dlygate4sd3_1
X_16106_ _03722_ _03827_ _03830_ _03730_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__a211o_1
Xhold818 CPU.registerFile\[27\]\[0\] VGND VGND VPWR VPWR net2115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold829 CPU.registerFile\[14\]\[12\] VGND VGND VPWR VPWR net2126 sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ CPU.registerFile\[27\]\[0\] CPU.registerFile\[26\]\[0\] _06063_ VGND VGND
+ VPWR VPWR _08544_ sky130_fd_sc_hd__mux2_1
X_17086_ CPU.registerFile\[28\]\[26\] CPU.registerFile\[29\]\[26\] _04526_ VGND VGND
+ VPWR VPWR _04787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16037_ _03760_ _03762_ _03763_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17988_ net999 _01516_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_16939_ CPU.registerFile\[28\]\[22\] CPU.registerFile\[29\]\[22\] _04526_ VGND VGND
+ VPWR VPWR _04644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09411_ _05698_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__clkbuf_4
X_18609_ net430 _02133_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13296__798 clknet_1_1__leaf__08361_ VGND VGND VPWR VPWR net854 sky130_fd_sc_hd__inv_2
XFILLER_0_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_16
X_09342_ _05684_ _05686_ _05693_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09273_ CPU.aluIn1\[16\] _05543_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__08449_ clknet_0__08449_ VGND VGND VPWR VPWR clknet_1_1__leaf__08449_
+ sky130_fd_sc_hd__clkbuf_16
X_13606__989 clknet_1_0__leaf__08445_ VGND VGND VPWR VPWR net1045 sky130_fd_sc_hd__inv_2
X_15934__672 clknet_1_1__leaf__03689_ VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__inv_2
XFILLER_0_139_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08988_ CPU.aluIn1\[16\] _05339_ VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10950_ _06992_ _07003_ VGND VGND VPWR VPWR _07004_ sky130_fd_sc_hd__and2_1
Xclkbuf_1_0__f__08340_ clknet_0__08340_ VGND VGND VPWR VPWR clknet_1_0__leaf__08340_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09609_ CPU.Iimm\[2\] CPU.instr\[3\] VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__nand2_1
X_10881_ CPU.aluReg\[7\] _06950_ _06922_ VGND VGND VPWR VPWR _06951_ sky130_fd_sc_hd__mux2_1
X_12620_ _08001_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__clkbuf_1
X_13355__851 clknet_1_0__leaf__08367_ VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__inv_2
XFILLER_0_38_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12551_ net1871 _07326_ _07957_ VGND VGND VPWR VPWR _07965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11502_ _06412_ VGND VGND VPWR VPWR _07364_ sky130_fd_sc_hd__clkbuf_4
X_12482_ net2132 _07326_ _07920_ VGND VGND VPWR VPWR _07928_ sky130_fd_sc_hd__mux2_1
X_15270_ CPU.registerFile\[28\]\[23\] CPU.registerFile\[29\]\[23\] _03212_ VGND VGND
+ VPWR VPWR _03329_ sky130_fd_sc_hd__mux2_1
X_17321__734 clknet_1_0__leaf__04982_ VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__inv_2
XFILLER_0_123_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11433_ _07317_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11364_ net1797 _05825_ _07274_ VGND VGND VPWR VPWR _07279_ sky130_fd_sc_hd__mux2_1
X_13103_ _07687_ _07782_ net1298 VGND VGND VPWR VPWR _08258_ sky130_fd_sc_hd__o21ai_1
X_10315_ _05785_ VGND VGND VPWR VPWR _06601_ sky130_fd_sc_hd__clkbuf_4
X_18960_ net734 _02480_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_11295_ _07242_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ CPU.registerFile\[4\]\[27\] net1339 _08217_ VGND VGND VPWR VPWR _08222_ sky130_fd_sc_hd__mux2_1
X_17911_ clknet_leaf_23_clk _01439_ VGND VGND VPWR VPWR CPU.Jimm\[18\] sky130_fd_sc_hd__dfxtp_1
X_10246_ _06562_ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__clkbuf_1
X_18891_ net665 _02411_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_17842_ net922 _01404_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_10177_ _05435_ _05439_ _05440_ VGND VGND VPWR VPWR _06500_ sky130_fd_sc_hd__a21oi_1
X_17773_ net853 _01335_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_14985_ _03049_ _03050_ CPU.registerFile\[25\]\[16\] VGND VGND VPWR VPWR _03051_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16724_ CPU.registerFile\[0\]\[17\] _04233_ _04068_ _04433_ VGND VGND VPWR VPWR _04434_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16655_ _03765_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__08469_ clknet_0__08469_ VGND VGND VPWR VPWR clknet_1_0__leaf__08469_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12818_ net1634 VGND VGND VPWR VPWR _08107_ sky130_fd_sc_hd__inv_2
X_16586_ CPU.registerFile\[8\]\[14\] _04101_ _04102_ _04298_ VGND VGND VPWR VPWR _04299_
+ sky130_fd_sc_hd__o211a_1
X_13798_ clknet_1_0__leaf__08462_ VGND VGND VPWR VPWR _08465_ sky130_fd_sc_hd__buf_1
XFILLER_0_158_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13786__1151 clknet_1_0__leaf__08463_ VGND VGND VPWR VPWR net1207 sky130_fd_sc_hd__inv_2
X_18325_ net146 _01853_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_15537_ CPU.registerFile\[8\]\[30\] _08545_ _03588_ _03268_ VGND VGND VPWR VPWR _03589_
+ sky130_fd_sc_hd__o211a_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _06605_ net2148 _08065_ VGND VGND VPWR VPWR _08070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18256_ net1267 _01784_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_15468_ CPU.registerFile\[5\]\[28\] CPU.registerFile\[4\]\[28\] _08558_ VGND VGND
+ VPWR VPWR _03522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17207_ _08397_ _04902_ _04904_ _08400_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__a211o_1
XFILLER_0_142_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14419_ _08557_ _08657_ _08662_ _08423_ VGND VGND VPWR VPWR _08663_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18187_ net1198 net1374 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[26\] sky130_fd_sc_hd__dfxtp_1
X_15399_ _03235_ _03236_ CPU.registerFile\[1\]\[26\] VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold604 CPU.registerFile\[6\]\[10\] VGND VGND VPWR VPWR net1901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17138_ _04545_ _04820_ _04837_ _04500_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__a211o_2
XFILLER_0_142_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold615 CPU.registerFile\[3\]\[17\] VGND VGND VPWR VPWR net1912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 CPU.registerFile\[18\]\[10\] VGND VGND VPWR VPWR net1923 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold637 CPU.registerFile\[22\]\[21\] VGND VGND VPWR VPWR net1934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold648 CPU.registerFile\[27\]\[7\] VGND VGND VPWR VPWR net1945 sky130_fd_sc_hd__dlygate4sd3_1
X_17069_ CPU.registerFile\[9\]\[26\] _04460_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__or2_1
Xhold659 CPU.registerFile\[27\]\[18\] VGND VGND VPWR VPWR net1956 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ _06291_ VGND VGND VPWR VPWR _06292_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_6_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08911_ CPU.aluIn1\[8\] _05262_ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__and2_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09891_ _06225_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__clkbuf_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14233__363 clknet_1_0__leaf__08508_ VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__inv_2
XFILLER_0_110_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1304 CPU.registerFile\[12\]\[17\] VGND VGND VPWR VPWR net2601 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1315 mapped_spi_flash.rcv_data\[13\] VGND VGND VPWR VPWR net2612 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1326 CPU.registerFile\[25\]\[18\] VGND VGND VPWR VPWR net2623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1337 mapped_spi_flash.rcv_bitcount\[1\] VGND VGND VPWR VPWR net2634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1348 CPU.aluIn1\[16\] VGND VGND VPWR VPWR net2645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1359 CPU.aluReg\[20\] VGND VGND VPWR VPWR net2656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18233__17 VGND VGND VPWR VPWR _18233__17/HI net17 sky130_fd_sc_hd__conb_1
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13670__1046 clknet_1_0__leaf__08452_ VGND VGND VPWR VPWR net1102 sky130_fd_sc_hd__inv_2
XFILLER_0_95_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09325_ CPU.PC\[19\] _05636_ _05675_ _05676_ net2 VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__o221a_2
XFILLER_0_48_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09256_ _05606_ _05607_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_647 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09187_ CPU.instr\[6\] _05243_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__nor2_1
XFILLER_0_161_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10100_ CPU.cycles\[5\] _05553_ _06368_ _06422_ _06425_ VGND VGND VPWR VPWR _06426_
+ sky130_fd_sc_hd__a221o_1
X_11080_ mapped_spi_flash.state\[2\] mapped_spi_flash.state\[1\] mapped_spi_flash.state\[0\]
+ _05703_ VGND VGND VPWR VPWR _07110_ sky130_fd_sc_hd__o31a_1
Xclkbuf_1_0__f__04983_ clknet_0__04983_ VGND VGND VPWR VPWR clknet_1_0__leaf__04983_
+ sky130_fd_sc_hd__clkbuf_16
X_10031_ _06343_ _06353_ _06359_ VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__or3b_4
XFILLER_0_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14770_ CPU.registerFile\[19\]\[11\] CPU.registerFile\[18\]\[11\] _02753_ VGND VGND
+ VPWR VPWR _02841_ sky130_fd_sc_hd__mux2_1
X_11982_ _06643_ net2089 _07620_ VGND VGND VPWR VPWR _07623_ sky130_fd_sc_hd__mux2_1
X_10933_ _06854_ VGND VGND VPWR VPWR _06992_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16440_ CPU.registerFile\[0\]\[10\] _03828_ _04068_ _04156_ VGND VGND VPWR VPWR _04157_
+ sky130_fd_sc_hd__o211a_1
X_10864_ net2665 _06937_ _06922_ VGND VGND VPWR VPWR _06938_ sky130_fd_sc_hd__mux2_1
X_12603_ _06595_ _07633_ VGND VGND VPWR VPWR _07992_ sky130_fd_sc_hd__nand2_4
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16371_ _06534_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__clkbuf_4
X_10795_ CPU.aluIn1\[27\] _06884_ _06881_ VGND VGND VPWR VPWR _06885_ sky130_fd_sc_hd__mux2_1
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15761__550 clknet_1_1__leaf__03653_ VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__inv_2
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18110_ net1121 _01638_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15322_ CPU.registerFile\[6\]\[24\] CPU.registerFile\[7\]\[24\] _08536_ VGND VGND
+ VPWR VPWR _03380_ sky130_fd_sc_hd__mux2_1
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12534_ _06594_ VGND VGND VPWR VPWR _07955_ sky130_fd_sc_hd__inv_2
X_19090_ net73 _02610_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[2\] sky130_fd_sc_hd__dfxtp_1
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18041_ net1052 _01569_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_15253_ CPU.registerFile\[2\]\[22\] CPU.registerFile\[3\]\[22\] _03275_ VGND VGND
+ VPWR VPWR _03313_ sky130_fd_sc_hd__mux2_1
X_12465_ _07918_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11416_ net2182 _06508_ _07296_ VGND VGND VPWR VPWR _07306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12396_ _06661_ net1990 _07847_ VGND VGND VPWR VPWR _07882_ sky130_fd_sc_hd__mux2_1
X_15184_ CPU.registerFile\[19\]\[21\] CPU.registerFile\[18\]\[21\] _03157_ VGND VGND
+ VPWR VPWR _03245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11347_ _07269_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11278_ _07232_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__clkbuf_1
X_18943_ net717 _02463_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_13017_ _08212_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__clkbuf_1
X_10229_ _06521_ _05520_ _05528_ VGND VGND VPWR VPWR _06550_ sky130_fd_sc_hd__a21oi_1
X_18874_ net648 _02394_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_17825_ net905 _01387_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold1 net1358 VGND VGND VPWR VPWR net1298 sky130_fd_sc_hd__buf_2
XFILLER_0_89_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17756_ clknet_leaf_25_clk _00000_ VGND VGND VPWR VPWR CPU.state\[1\] sky130_fd_sc_hd__dfxtp_2
X_14968_ net1647 _02797_ _03034_ _02993_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__o211a_1
X_16707_ CPU.registerFile\[8\]\[17\] _04101_ _04102_ _04416_ VGND VGND VPWR VPWR _04417_
+ sky130_fd_sc_hd__o211a_1
X_17687_ _05215_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__clkbuf_1
X_14899_ _02965_ _02966_ _02851_ VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16638_ CPU.registerFile\[0\]\[15\] _04233_ _04068_ _04349_ VGND VGND VPWR VPWR _04350_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16569_ CPU.registerFile\[24\]\[13\] _03915_ _04165_ _04282_ VGND VGND VPWR VPWR
+ _04283_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09110_ _05451_ _05460_ _05461_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__o21a_1
X_18308_ net129 _01836_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09041_ CPU.aluIn1\[27\] _05392_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__and2_1
X_18239_ net1250 _01767_ VGND VGND VPWR VPWR mapped_spi_ram.rbusy sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13230__752 clknet_1_1__leaf__08342_ VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__inv_2
XFILLER_0_142_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold401 CPU.registerFile\[6\]\[23\] VGND VGND VPWR VPWR net1698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold412 CPU.registerFile\[5\]\[14\] VGND VGND VPWR VPWR net1709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 CPU.registerFile\[6\]\[8\] VGND VGND VPWR VPWR net1720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 CPU.registerFile\[22\]\[0\] VGND VGND VPWR VPWR net1731 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 CPU.registerFile\[10\]\[20\] VGND VGND VPWR VPWR net1742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold456 CPU.registerFile\[5\]\[6\] VGND VGND VPWR VPWR net1753 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 CPU.registerFile\[10\]\[10\] VGND VGND VPWR VPWR net1764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold478 CPU.registerFile\[30\]\[23\] VGND VGND VPWR VPWR net1775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 CPU.registerFile\[27\]\[23\] VGND VGND VPWR VPWR net1786 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ _05453_ _06274_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__xor2_1
XFILLER_0_96_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _05514_ _05550_ _05553_ CPU.cycles\[14\] VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__a22o_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 CPU.registerFile\[14\]\[26\] VGND VGND VPWR VPWR net2398 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1112 CPU.registerFile\[14\]\[3\] VGND VGND VPWR VPWR net2409 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1123 CPU.aluIn1\[30\] VGND VGND VPWR VPWR net2420 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1134 CPU.registerFile\[25\]\[23\] VGND VGND VPWR VPWR net2431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 CPU.registerFile\[14\]\[2\] VGND VGND VPWR VPWR net2442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1156 CPU.registerFile\[8\]\[12\] VGND VGND VPWR VPWR net2453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 CPU.registerFile\[9\]\[20\] VGND VGND VPWR VPWR net2464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1178 CPU.registerFile\[21\]\[20\] VGND VGND VPWR VPWR net2475 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03650_ clknet_0__03650_ VGND VGND VPWR VPWR clknet_1_0__leaf__03650_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 CPU.registerFile\[17\]\[13\] VGND VGND VPWR VPWR net2486 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09308_ _05626_ _05627_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10580_ _06756_ VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09239_ CPU.aluIn1\[5\] CPU.Bimm\[5\] VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12250_ net1551 _07785_ _07797_ _07796_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11201_ _07130_ _07188_ VGND VGND VPWR VPWR _07190_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12181_ mapped_spi_ram.cmd_addr\[5\] _07749_ _07706_ CPU.mem_wdata\[6\] _07739_ VGND
+ VGND VPWR VPWR _07750_ sky130_fd_sc_hd__a221o_1
X_11132_ net1602 _07133_ _07146_ _07138_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__o211a_1
Xhold990 CPU.registerFile\[8\]\[11\] VGND VGND VPWR VPWR net2287 sky130_fd_sc_hd__dlygate4sd3_1
X_11063_ _07048_ _07098_ VGND VGND VPWR VPWR _07099_ sky130_fd_sc_hd__or2_1
X_13785__1150 clknet_1_0__leaf__08463_ VGND VGND VPWR VPWR net1206 sky130_fd_sc_hd__inv_2
X_10014_ _06202_ _06342_ _06177_ VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__o21a_1
X_17610_ per_uart.d_in_uart\[4\] _05134_ _05157_ per_uart.uart0.txd_reg\[5\] VGND
+ VGND VPWR VPWR _05163_ sky130_fd_sc_hd__o22a_1
X_14822_ _08808_ _08809_ CPU.registerFile\[25\]\[12\] VGND VGND VPWR VPWR _02892_
+ sky130_fd_sc_hd__a21o_1
X_18590_ net411 net47 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17541_ _08335_ _06019_ _05073_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__o21ai_1
X_14753_ _02728_ _02820_ _02824_ _02784_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11965_ _06626_ net2201 _07609_ VGND VGND VPWR VPWR _07614_ sky130_fd_sc_hd__mux2_1
X_10916_ mapped_spi_flash.snd_bitcount\[3\] mapped_spi_flash.snd_bitcount\[2\] VGND
+ VGND VPWR VPWR _06978_ sky130_fd_sc_hd__or2_1
X_17472_ _08379_ _05017_ _06306_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__o21bai_1
X_14684_ _06036_ VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__clkbuf_4
X_11896_ _07577_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__clkbuf_1
X_15685__481 clknet_1_1__leaf__03646_ VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__inv_2
X_17327__740 clknet_1_1__leaf__04982_ VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__inv_2
X_16423_ CPU.aluIn1\[9\] _04054_ _04140_ _03855_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__o211a_1
X_10847_ CPU.aluIn1\[15\] _06924_ _06914_ VGND VGND VPWR VPWR _06925_ sky130_fd_sc_hd__mux2_1
X_19142_ clknet_leaf_7_clk _02662_ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dfxtp_2
X_16354_ _03901_ _04066_ _04071_ _04072_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10778_ _05514_ _06175_ VGND VGND VPWR VPWR _06871_ sky130_fd_sc_hd__nor2_2
X_15305_ CPU.registerFile\[30\]\[24\] CPU.registerFile\[31\]\[24\] _03291_ VGND VGND
+ VPWR VPWR _03363_ sky130_fd_sc_hd__mux2_1
X_12517_ _07946_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__clkbuf_1
X_19073_ net65 _02593_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_16285_ _06141_ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18024_ net1035 _01552_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_15236_ _03049_ _03050_ CPU.registerFile\[25\]\[22\] VGND VGND VPWR VPWR _03296_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12448_ net1780 _07360_ _07906_ VGND VGND VPWR VPWR _07910_ sky130_fd_sc_hd__mux2_1
X_15167_ _03133_ _03224_ _03228_ _03188_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12379_ _07873_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13522__913 clknet_1_1__leaf__08437_ VGND VGND VPWR VPWR net969 sky130_fd_sc_hd__inv_2
Xclkbuf_0__03644_ _03644_ VGND VGND VPWR VPWR clknet_0__03644_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15098_ _06036_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__clkbuf_4
X_18926_ net700 _02446_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18857_ net631 _02377_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_09590_ CPU.Jimm\[15\] _05921_ _05923_ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__a21o_1
X_17808_ net888 _01370_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_18788_ net577 _02312_ VGND VGND VPWR VPWR CPU.aluReg\[18\] sky130_fd_sc_hd__dfxtp_1
X_17739_ net824 _01305_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09024_ CPU.aluIn1\[22\] _05375_ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13750__1119 clknet_1_1__leaf__08459_ VGND VGND VPWR VPWR net1175 sky130_fd_sc_hd__inv_2
Xhold220 _01711_ VGND VGND VPWR VPWR net1517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 CPU.cycles\[11\] VGND VGND VPWR VPWR net1528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 _08290_ VGND VGND VPWR VPWR net1539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _08306_ VGND VGND VPWR VPWR net1550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _08294_ VGND VGND VPWR VPWR net1561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 mapped_spi_ram.rcv_data\[17\] VGND VGND VPWR VPWR net1572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 CPU.cycles\[12\] VGND VGND VPWR VPWR net1583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 CPU.rs2\[25\] VGND VGND VPWR VPWR net1594 sky130_fd_sc_hd__dlygate4sd3_1
X_09926_ _05316_ _05533_ _05535_ net1405 _06258_ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__a221o_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _05326_ _05533_ _05536_ net1414 _06192_ VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__a221o_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _05425_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__clkbuf_4
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13949__108 clknet_1_0__leaf__08479_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__inv_2
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11750_ _06615_ net2226 _07490_ VGND VGND VPWR VPWR _07500_ sky130_fd_sc_hd__mux2_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ net1784 _05853_ _06816_ VGND VGND VPWR VPWR _06823_ sky130_fd_sc_hd__mux2_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11681_ net2402 _07330_ _07453_ VGND VGND VPWR VPWR _07463_ sky130_fd_sc_hd__mux2_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13420_ _08389_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__clkbuf_1
X_10632_ net2596 _05873_ _06777_ VGND VGND VPWR VPWR _06785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10563_ _06747_ VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12302_ net4 _07784_ _07826_ _07822_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__o211a_1
X_16070_ _03736_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__buf_4
XFILLER_0_134_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10494_ _06710_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15021_ CPU.registerFile\[28\]\[17\] CPU.registerFile\[29\]\[17\] _02808_ VGND VGND
+ VPWR VPWR _03086_ sky130_fd_sc_hd__mux2_1
X_12233_ net1427 _07785_ _07788_ _07755_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12164_ _07692_ VGND VGND VPWR VPWR _07738_ sky130_fd_sc_hd__buf_2
X_11115_ _07001_ VGND VGND VPWR VPWR _07138_ sky130_fd_sc_hd__clkbuf_4
X_12095_ mapped_spi_ram.snd_bitcount\[5\] mapped_spi_ram.snd_bitcount\[4\] mapped_spi_ram.snd_bitcount\[0\]
+ VGND VGND VPWR VPWR _07689_ sky130_fd_sc_hd__or3b_1
X_16972_ _04389_ _04390_ CPU.registerFile\[1\]\[23\] VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__a21o_1
X_18711_ net500 _02235_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[11\] sky130_fd_sc_hd__dfxtp_1
X_11046_ _07083_ _05593_ VGND VGND VPWR VPWR _07084_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18642_ clknet_leaf_14_clk _02166_ VGND VGND VPWR VPWR CPU.rs2\[14\] sky130_fd_sc_hd__dfxtp_1
X_14805_ _02826_ _02870_ _02875_ _02746_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__o211a_1
X_18573_ net394 net30 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_14067__214 clknet_1_0__leaf__08491_ VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__inv_2
X_15785_ _03658_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__clkbuf_4
X_12997_ net2306 _07351_ _08192_ VGND VGND VPWR VPWR _08202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17524_ _05055_ _06088_ _05061_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__or3_1
XFILLER_0_86_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14736_ _08409_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__buf_4
X_11948_ _06609_ net2556 _07598_ VGND VGND VPWR VPWR _07605_ sky130_fd_sc_hd__mux2_1
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17455_ _05022_ _06406_ _08256_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__o21ai_1
X_14667_ _02739_ _02740_ _08783_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__mux2_1
X_11879_ _07568_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16406_ _04121_ _04123_ _03875_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__mux2_1
X_17386_ _04996_ _05009_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14598_ _08520_ VGND VGND VPWR VPWR _08837_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19125_ clknet_leaf_10_clk _02645_ VGND VGND VPWR VPWR CPU.PC\[7\] sky130_fd_sc_hd__dfxtp_1
X_16337_ _03697_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__buf_2
XFILLER_0_109_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19056_ net798 _02576_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_16268_ _03943_ _03984_ _03988_ _03730_ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_1__f__08482_ clknet_0__08482_ VGND VGND VPWR VPWR clknet_1_1__leaf__08482_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_124_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18007_ net1018 _01535_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_15219_ _03230_ _03274_ _03279_ _03151_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__o211a_1
X_16199_ _03920_ _03921_ _03763_ VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13303__804 clknet_1_0__leaf__08362_ VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__inv_2
X_09711_ _05764_ _06038_ _06049_ _06052_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__a211o_4
X_18909_ net683 _02429_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_09642_ _05939_ _05979_ _05983_ _05985_ _05982_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__a32o_1
X_18578__35 VGND VGND VPWR VPWR _18578__35/HI net35 sky130_fd_sc_hd__conb_1
X_09573_ CPU.Iimm\[2\] _05545_ _05914_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__mux2_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13492__886 clknet_1_0__leaf__08434_ VGND VGND VPWR VPWR net942 sky130_fd_sc_hd__inv_2
XFILLER_0_136_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09007_ _05344_ _05347_ _05352_ _05357_ _05358_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_130_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09909_ _06202_ _06242_ _06177_ VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__o21a_1
X_14016__168 clknet_1_0__leaf__08486_ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__inv_2
X_12920_ _08161_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__clkbuf_1
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12851_ _06145_ net2495 _08120_ VGND VGND VPWR VPWR _08125_ sky130_fd_sc_hd__mux2_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ net2082 _07314_ _07526_ VGND VGND VPWR VPWR _07528_ sky130_fd_sc_hd__mux2_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ CPU.registerFile\[13\]\[31\] CPU.registerFile\[12\]\[31\] _08794_ VGND VGND
+ VPWR VPWR _03621_ sky130_fd_sc_hd__mux2_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _08064_ VGND VGND VPWR VPWR _08087_ sky130_fd_sc_hd__buf_4
XFILLER_0_68_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ CPU.registerFile\[28\]\[5\] CPU.registerFile\[29\]\[5\] _08538_ VGND VGND
+ VPWR VPWR _08762_ sky130_fd_sc_hd__mux2_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _07491_ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__clkbuf_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15905__647 clknet_1_1__leaf__03685_ VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__inv_2
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17240_ CPU.registerFile\[19\]\[30\] CPU.registerFile\[18\]\[30\] _03745_ VGND VGND
+ VPWR VPWR _04937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14452_ _08540_ VGND VGND VPWR VPWR _08695_ sky130_fd_sc_hd__buf_4
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _07454_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__clkbuf_1
X_15604__408 clknet_1_1__leaf__03638_ VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__inv_2
XFILLER_0_37_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13403_ _08380_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10615_ _05739_ _05737_ _05738_ VGND VGND VPWR VPWR _06775_ sky130_fd_sc_hd__or3_2
X_17171_ _08397_ _04867_ _04869_ _08400_ VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__a211o_1
XFILLER_0_119_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14383_ _08626_ _08627_ _08578_ VGND VGND VPWR VPWR _08628_ sky130_fd_sc_hd__mux2_1
X_11595_ _07417_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16122_ _06171_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10546_ _06737_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__buf_2
X_16053_ CPU.registerFile\[10\]\[1\] CPU.registerFile\[11\]\[1\] _03694_ VGND VGND
+ VPWR VPWR _03779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13265_ net1514 net1500 VGND VGND VPWR VPWR _08346_ sky130_fd_sc_hd__or2_1
X_10477_ _06700_ VGND VGND VPWR VPWR _06701_ sky130_fd_sc_hd__clkbuf_4
X_15004_ _03027_ _03067_ _03069_ _08870_ VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__a211o_1
X_12216_ _07770_ _07774_ _07764_ VGND VGND VPWR VPWR _07775_ sky130_fd_sc_hd__a21oi_1
X_17290__706 clknet_1_1__leaf__04979_ VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__inv_2
X_13196_ _05547_ VGND VGND VPWR VPWR _08310_ sky130_fd_sc_hd__buf_2
X_12147_ net1485 _07714_ _07726_ _07713_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12078_ _07675_ net1302 VGND VGND VPWR VPWR _07677_ sky130_fd_sc_hd__or2_1
X_16955_ _04574_ _04654_ _04659_ _04584_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__o211a_1
X_11029_ net1518 _07054_ _07068_ _07069_ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__o211a_1
X_16886_ CPU.registerFile\[15\]\[21\] CPU.registerFile\[14\]\[21\] _04550_ VGND VGND
+ VPWR VPWR _04592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18625_ net446 _02149_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__05013_ _05013_ VGND VGND VPWR VPWR clknet_0__05013_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13628__1009 clknet_1_1__leaf__08447_ VGND VGND VPWR VPWR net1065 sky130_fd_sc_hd__inv_2
X_18556_ net377 _02080_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14719_ CPU.registerFile\[0\]\[9\] _08706_ _02790_ _02791_ VGND VGND VPWR VPWR _02792_
+ sky130_fd_sc_hd__o211a_1
X_17507_ _05069_ CPU.PC\[15\] _05082_ _05083_ _05053_ VGND VGND VPWR VPWR _02653_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_157_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18487_ net308 _02011_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17438_ _06468_ _05024_ _05026_ _05880_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__a211o_1
XFILLER_0_129_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_15 _04120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _04803_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 _07452_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_48 clknet_1_0__leaf__03656_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17369_ _04998_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_59 clknet_1_0__leaf__08440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19108_ net91 _02628_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_918 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19039_ net781 _02559_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13978__134 clknet_1_0__leaf__08482_ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__08465_ clknet_0__08465_ VGND VGND VPWR VPWR clknet_1_1__leaf__08465_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08496_ _08496_ VGND VGND VPWR VPWR clknet_0__08496_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13500__893 clknet_1_0__leaf__08435_ VGND VGND VPWR VPWR net949 sky130_fd_sc_hd__inv_2
X_09625_ _05947_ _05967_ _05968_ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__a21o_1
X_09556_ _05379_ _05899_ _05493_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09487_ _05793_ _05830_ _05832_ _05833_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14204__338 clknet_1_1__leaf__08504_ VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__inv_2
XFILLER_0_108_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10400_ _06658_ VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11380_ _07287_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10331_ _06611_ net1949 _06597_ VGND VGND VPWR VPWR _06612_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13050_ _08230_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10262_ net1850 _06083_ _06569_ VGND VGND VPWR VPWR _06571_ sky130_fd_sc_hd__mux2_1
X_12001_ _07632_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__clkbuf_1
X_10193_ _06391_ _06511_ _06514_ VGND VGND VPWR VPWR _06515_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16740_ _04448_ _04449_ _04365_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_918 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12903_ _08152_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__clkbuf_1
X_16671_ CPU.registerFile\[12\]\[16\] _04017_ _04018_ _04381_ VGND VGND VPWR VPWR
+ _04382_ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_0__f__08485_ clknet_0__08485_ VGND VGND VPWR VPWR clknet_1_0__leaf__08485_
+ sky130_fd_sc_hd__clkbuf_16
X_18410_ net231 _01938_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12834_ _05853_ net2289 _08109_ VGND VGND VPWR VPWR _08116_ sky130_fd_sc_hd__mux2_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15829__578 clknet_1_0__leaf__03678_ VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__inv_2
XFILLER_0_97_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18341_ net162 _01869_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ CPU.registerFile\[17\]\[31\] _08528_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__or2_1
X_12765_ _08078_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__clkbuf_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14504_ CPU.registerFile\[0\]\[4\] _08706_ _08745_ _08588_ VGND VGND VPWR VPWR _08746_
+ sky130_fd_sc_hd__o211a_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _07481_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__clkbuf_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18272_ net1283 _01800_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15484_ CPU.registerFile\[20\]\[29\] _08523_ _03536_ _08578_ VGND VGND VPWR VPWR
+ _03537_ sky130_fd_sc_hd__o211a_1
X_12696_ _06620_ net2543 _08040_ VGND VGND VPWR VPWR _08042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17223_ CPU.registerFile\[2\]\[30\] CPU.registerFile\[3\]\[30\] _03759_ VGND VGND
+ VPWR VPWR _04920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14435_ CPU.registerFile\[22\]\[3\] CPU.registerFile\[23\]\[3\] _08523_ VGND VGND
+ VPWR VPWR _08678_ sky130_fd_sc_hd__mux2_1
X_11647_ _07444_ VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__clkbuf_1
X_14179__315 clknet_1_0__leaf__08502_ VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__inv_2
XFILLER_0_142_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17154_ _03765_ _04850_ _04852_ _04521_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__a211o_1
X_14366_ CPU.registerFile\[27\]\[1\] CPU.registerFile\[26\]\[1\] _06063_ VGND VGND
+ VPWR VPWR _08611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11578_ _07407_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__clkbuf_1
X_16105_ CPU.registerFile\[0\]\[2\] _03828_ _03725_ _03829_ VGND VGND VPWR VPWR _03830_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold808 CPU.registerFile\[13\]\[26\] VGND VGND VPWR VPWR net2105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17085_ CPU.registerFile\[30\]\[26\] CPU.registerFile\[31\]\[26\] _04605_ VGND VGND
+ VPWR VPWR _04786_ sky130_fd_sc_hd__mux2_1
Xhold819 CPU.registerFile\[23\]\[14\] VGND VGND VPWR VPWR net2116 sky130_fd_sc_hd__dlygate4sd3_1
X_10529_ net2387 _06386_ _06724_ VGND VGND VPWR VPWR _06729_ sky130_fd_sc_hd__mux2_1
X_14297_ _06418_ VGND VGND VPWR VPWR _08543_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16036_ _03741_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__buf_4
XFILLER_0_122_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13179_ _08299_ _08300_ VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__nor2_1
X_17987_ net998 _01515_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_13558__945 clknet_1_1__leaf__08441_ VGND VGND VPWR VPWR net1001 sky130_fd_sc_hd__inv_2
X_16938_ CPU.registerFile\[30\]\[22\] CPU.registerFile\[31\]\[22\] _04605_ VGND VGND
+ VPWR VPWR _04643_ sky130_fd_sc_hd__mux2_1
X_16869_ CPU.registerFile\[20\]\[20\] CPU.registerFile\[21\]\[20\] _04287_ VGND VGND
+ VPWR VPWR _04576_ sky130_fd_sc_hd__mux2_1
X_09410_ _05685_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__buf_2
X_18608_ net429 _02132_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09341_ _05577_ _05579_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__xnor2_4
X_18539_ net360 _02063_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09272_ CPU.aluIn1\[17\] _05543_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14045__194 clknet_1_1__leaf__08489_ VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__inv_2
XFILLER_0_7_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13309__810 clknet_1_1__leaf__08362_ VGND VGND VPWR VPWR net866 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__08448_ clknet_0__08448_ VGND VGND VPWR VPWR clknet_1_1__leaf__08448_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__08479_ _08479_ VGND VGND VPWR VPWR clknet_0__08479_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08987_ CPU.rs2\[16\] _05246_ _05250_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__o21a_1
X_15633__434 clknet_1_0__leaf__03641_ VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__inv_2
XFILLER_0_98_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09608_ CPU.Iimm\[1\] CPU.instr\[3\] _05922_ CPU.Bimm\[1\] VGND VGND VPWR VPWR _05952_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10880_ CPU.aluIn1\[7\] _06949_ _06880_ VGND VGND VPWR VPWR _06950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09539_ CPU.PC\[5\] _05882_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__and2_1
X_14128__269 clknet_1_0__leaf__08497_ VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__inv_2
X_12550_ _07964_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11501_ _07363_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12481_ _07927_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14220_ clknet_1_1__leaf__08506_ VGND VGND VPWR VPWR _08507_ sky130_fd_sc_hd__buf_1
XFILLER_0_62_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11432_ net1700 _07316_ _07312_ VGND VGND VPWR VPWR _07317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11363_ _07278_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13102_ net1623 _08257_ _06856_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__o21a_1
X_13627__1008 clknet_1_1__leaf__08447_ VGND VGND VPWR VPWR net1064 sky130_fd_sc_hd__inv_2
X_10314_ _06600_ VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_934 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11294_ net2110 _05805_ _07238_ VGND VGND VPWR VPWR _07242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15716__509 clknet_1_1__leaf__03649_ VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__inv_2
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ net1403 VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__clkbuf_1
X_17910_ clknet_leaf_23_clk _01438_ VGND VGND VPWR VPWR CPU.Jimm\[17\] sky130_fd_sc_hd__dfxtp_1
X_10245_ net1807 _05805_ _06558_ VGND VGND VPWR VPWR _06562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18890_ net664 _02410_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17841_ net921 _01403_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_10176_ _05424_ _06498_ VGND VGND VPWR VPWR _06499_ sky130_fd_sc_hd__nand2_1
X_17772_ net852 _01334_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_14984_ _06059_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__clkbuf_4
X_16723_ _04389_ _04390_ CPU.registerFile\[1\]\[17\] VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__a21o_1
X_16654_ _04363_ _04364_ _04365_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__08468_ clknet_0__08468_ VGND VGND VPWR VPWR clknet_1_0__leaf__08468_
+ sky130_fd_sc_hd__clkbuf_16
X_12817_ _05434_ _06861_ _08106_ _08104_ _06869_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__o221a_1
X_16585_ CPU.registerFile\[9\]\[14\] _04056_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__or2_1
X_15536_ _08546_ _08547_ CPU.registerFile\[9\]\[30\] VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__a21o_1
X_18324_ net145 _01852_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12748_ _08069_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__clkbuf_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18255_ net1266 _01783_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_15467_ CPU.registerFile\[6\]\[28\] CPU.registerFile\[7\]\[28\] _08536_ VGND VGND
+ VPWR VPWR _03521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12679_ _06603_ net2610 _08029_ VGND VGND VPWR VPWR _08033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17206_ CPU.registerFile\[16\]\[29\] _04656_ _06149_ _04903_ VGND VGND VPWR VPWR
+ _04904_ sky130_fd_sc_hd__o211a_1
X_14418_ _08520_ _08658_ _08660_ _08661_ VGND VGND VPWR VPWR _08662_ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18186_ net1197 _01714_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[25\] sky130_fd_sc_hd__dfxtp_1
X_15398_ CPU.registerFile\[2\]\[26\] CPU.registerFile\[3\]\[26\] _03275_ VGND VGND
+ VPWR VPWR _03454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17137_ _04828_ _04836_ _04542_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__o21a_1
X_14349_ _08573_ _08593_ _08594_ VGND VGND VPWR VPWR _08595_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold605 CPU.registerFile\[13\]\[16\] VGND VGND VPWR VPWR net1902 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold616 CPU.registerFile\[27\]\[13\] VGND VGND VPWR VPWR net1913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold627 CPU.registerFile\[18\]\[14\] VGND VGND VPWR VPWR net1924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 CPU.registerFile\[10\]\[19\] VGND VGND VPWR VPWR net1935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 CPU.registerFile\[19\]\[13\] VGND VGND VPWR VPWR net1946 sky130_fd_sc_hd__dlygate4sd3_1
X_17068_ CPU.registerFile\[10\]\[26\] CPU.registerFile\[11\]\[26\] _06173_ VGND VGND
+ VPWR VPWR _04769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16019_ CPU.registerFile\[27\]\[0\] CPU.registerFile\[26\]\[0\] _03745_ VGND VGND
+ VPWR VPWR _03746_ sky130_fd_sc_hd__mux2_1
X_08910_ CPU.rs2\[8\] CPU.Bimm\[8\] _05245_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__mux2_2
XFILLER_0_110_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ net2173 _06224_ _06055_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__mux2_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1305 CPU.registerFile\[26\]\[1\] VGND VGND VPWR VPWR net2602 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1316 mapped_spi_flash.rcv_data\[10\] VGND VGND VPWR VPWR net2613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1327 per_uart.uart0.rx_busy VGND VGND VPWR VPWR net2624 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1338 CPU.registerFile\[9\]\[3\] VGND VGND VPWR VPWR net2635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1349 CPU.registerFile\[25\]\[3\] VGND VGND VPWR VPWR net2646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09324_ _05674_ _05564_ _05673_ _05557_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13612__994 clknet_1_0__leaf__08446_ VGND VGND VPWR VPWR net1050 sky130_fd_sc_hd__inv_2
XFILLER_0_91_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09255_ CPU.aluIn1\[12\] CPU.Bimm\[12\] VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09186_ CPU.instr\[4\] VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__buf_2
XFILLER_0_43_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13385__878 clknet_1_0__leaf__08370_ VGND VGND VPWR VPWR net934 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__04982_ clknet_0__04982_ VGND VGND VPWR VPWR clknet_1_0__leaf__04982_
+ sky130_fd_sc_hd__clkbuf_16
X_10030_ _05911_ _06355_ _06357_ _06197_ _06358_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__o221a_1
X_11981_ _07622_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__clkbuf_1
X_13720_ clknet_1_1__leaf__08451_ VGND VGND VPWR VPWR _08457_ sky130_fd_sc_hd__buf_1
X_10932_ _06991_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10863_ CPU.aluIn1\[11\] _06936_ _06914_ VGND VGND VPWR VPWR _06937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12602_ _07991_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__clkbuf_1
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16370_ CPU.registerFile\[19\]\[8\] CPU.registerFile\[18\]\[8\] _03923_ VGND VGND
+ VPWR VPWR _04089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14061__209 clknet_1_1__leaf__08490_ VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__inv_2
XFILLER_0_27_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10794_ CPU.aluReg\[28\] CPU.aluReg\[26\] _06872_ VGND VGND VPWR VPWR _06884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15321_ _03133_ _03374_ _03378_ _03188_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12533_ _07954_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__clkbuf_1
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18040_ net1051 _01568_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15252_ _03310_ _03311_ _03025_ VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__mux2_1
X_12464_ net1683 _07376_ _07883_ VGND VGND VPWR VPWR _07918_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11415_ _07305_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__clkbuf_1
X_15183_ net1638 _03201_ _03244_ _02993_ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__o211a_1
X_12395_ _07881_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11346_ net2505 _06486_ _07260_ VGND VGND VPWR VPWR _07269_ sky130_fd_sc_hd__mux2_1
X_18942_ net716 _02462_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_11277_ _06655_ net1885 _07223_ VGND VGND VPWR VPWR _07232_ sky130_fd_sc_hd__mux2_1
X_13016_ net2339 _07370_ _08203_ VGND VGND VPWR VPWR _08212_ sky130_fd_sc_hd__mux2_1
X_10228_ CPU.aluIn1\[0\] _05276_ VGND VGND VPWR VPWR _06549_ sky130_fd_sc_hd__nor2_1
X_18873_ net647 _02393_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17824_ net904 _01386_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold2 _07845_ VGND VGND VPWR VPWR net1299 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10159_ _05818_ _06480_ _06482_ VGND VGND VPWR VPWR _06483_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17755_ clknet_leaf_1_clk _00001_ VGND VGND VPWR VPWR CPU.state\[0\] sky130_fd_sc_hd__dfxtp_1
X_14967_ _02750_ _03012_ _03033_ _02839_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__a211o_1
X_16706_ CPU.registerFile\[9\]\[17\] _04056_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17686_ _05207_ _05214_ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__and2_1
X_14898_ CPU.registerFile\[28\]\[14\] CPU.registerFile\[29\]\[14\] _02808_ VGND VGND
+ VPWR VPWR _02966_ sky130_fd_sc_hd__mux2_1
X_16637_ _03985_ _03986_ CPU.registerFile\[1\]\[15\] VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16568_ _04080_ _04081_ CPU.registerFile\[25\]\[13\] VGND VGND VPWR VPWR _04282_
+ sky130_fd_sc_hd__a21o_1
X_13863__1221 clknet_1_1__leaf__08470_ VGND VGND VPWR VPWR net1277 sky130_fd_sc_hd__inv_2
X_18307_ net128 _01835_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_15519_ CPU.registerFile\[22\]\[30\] CPU.registerFile\[23\]\[30\] _08584_ VGND VGND
+ VPWR VPWR _03571_ sky130_fd_sc_hd__mux2_1
X_15662__460 clknet_1_0__leaf__03644_ VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__inv_2
X_16499_ _04175_ _04176_ CPU.registerFile\[17\]\[11\] VGND VGND VPWR VPWR _04215_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09040_ CPU.rs2\[27\] _05247_ _05251_ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__o21a_1
X_18238_ net1249 _01766_ VGND VGND VPWR VPWR CPU.mem_wbusy sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18169_ net1180 net1455 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold402 CPU.registerFile\[10\]\[4\] VGND VGND VPWR VPWR net1699 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold413 CPU.registerFile\[28\]\[18\] VGND VGND VPWR VPWR net1710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold424 CPU.registerFile\[5\]\[21\] VGND VGND VPWR VPWR net1721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 CPU.registerFile\[6\]\[17\] VGND VGND VPWR VPWR net1732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 CPU.registerFile\[22\]\[29\] VGND VGND VPWR VPWR net1743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold457 CPU.registerFile\[19\]\[14\] VGND VGND VPWR VPWR net1754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 CPU.registerFile\[13\]\[20\] VGND VGND VPWR VPWR net1765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09942_ _05463_ _06273_ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__nand2_1
X_14157__295 clknet_1_0__leaf__08500_ VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__inv_2
Xhold479 CPU.registerFile\[13\]\[29\] VGND VGND VPWR VPWR net1776 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__03689_ clknet_0__03689_ VGND VGND VPWR VPWR clknet_1_1__leaf__03689_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ _06202_ _06207_ _06177_ VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__o21a_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 CPU.registerFile\[11\]\[13\] VGND VGND VPWR VPWR net2399 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 CPU.registerFile\[29\]\[15\] VGND VGND VPWR VPWR net2410 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1124 CPU.registerFile\[22\]\[7\] VGND VGND VPWR VPWR net2421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 CPU.registerFile\[23\]\[1\] VGND VGND VPWR VPWR net2432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 CPU.registerFile\[9\]\[2\] VGND VGND VPWR VPWR net2443 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1157 CPU.registerFile\[26\]\[13\] VGND VGND VPWR VPWR net2454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1168 CPU.registerFile\[12\]\[5\] VGND VGND VPWR VPWR net2465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 CPU.registerFile\[9\]\[14\] VGND VGND VPWR VPWR net2476 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13626__1007 clknet_1_1__leaf__08447_ VGND VGND VPWR VPWR net1063 sky130_fd_sc_hd__inv_2
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15745__535 clknet_1_0__leaf__03652_ VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__inv_2
XFILLER_0_119_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09307_ _05658_ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09238_ _05585_ _05589_ _05587_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_889 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09169_ _05514_ _05520_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__nand2_2
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11200_ _07189_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12180_ net1312 VGND VGND VPWR VPWR _07749_ sky130_fd_sc_hd__clkbuf_4
X_15639__440 clknet_1_1__leaf__03641_ VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__inv_2
X_11131_ net1416 _07135_ VGND VGND VPWR VPWR _07146_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold980 CPU.registerFile\[14\]\[17\] VGND VGND VPWR VPWR net2277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold991 CPU.registerFile\[14\]\[10\] VGND VGND VPWR VPWR net2288 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11062_ mapped_spi_flash.cmd_addr\[4\] _07097_ _07039_ VGND VGND VPWR VPWR _07098_
+ sky130_fd_sc_hd__mux2_1
X_10013_ CPU.Jimm\[13\] _06203_ _06339_ _06204_ _06341_ VGND VGND VPWR VPWR _06342_
+ sky130_fd_sc_hd__o32a_1
X_14821_ CPU.registerFile\[27\]\[12\] CPU.registerFile\[26\]\[12\] _02768_ VGND VGND
+ VPWR VPWR _02891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14752_ _08857_ _02821_ _02823_ _08661_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__a211o_1
X_17540_ _05108_ _05109_ _05058_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__a21oi_1
X_11964_ _07613_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__clkbuf_1
X_10915_ _06974_ mapped_spi_flash.snd_bitcount\[1\] mapped_spi_flash.snd_bitcount\[0\]
+ VGND VGND VPWR VPWR _06977_ sky130_fd_sc_hd__or3b_1
X_17471_ _05016_ net2590 _05051_ _05052_ _05053_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__o221a_1
X_14683_ CPU.registerFile\[17\]\[9\] _08795_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__or2_1
X_11895_ _06624_ net2383 _07573_ VGND VGND VPWR VPWR _07577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16422_ _03692_ _04120_ _04139_ _04096_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__a211o_1
X_10846_ CPU.aluReg\[16\] CPU.aluReg\[14\] _06906_ VGND VGND VPWR VPWR _06924_ sky130_fd_sc_hd__mux2_1
X_14262__390 clknet_1_0__leaf__08510_ VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__inv_2
XFILLER_0_6_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16353_ _06109_ VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__clkbuf_4
X_19141_ clknet_leaf_10_clk _02661_ VGND VGND VPWR VPWR CPU.PC\[23\] sky130_fd_sc_hd__dfxtp_2
X_13565_ clknet_1_1__leaf__08440_ VGND VGND VPWR VPWR _08442_ sky130_fd_sc_hd__buf_1
X_10777_ _06870_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15304_ _03078_ _03359_ _03361_ _03043_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__a211o_1
XFILLER_0_109_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12516_ net1914 _07360_ _07942_ VGND VGND VPWR VPWR _07946_ sky130_fd_sc_hd__mux2_1
X_19072_ net64 _02592_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_16284_ CPU.registerFile\[16\]\[6\] _03848_ _03769_ _04004_ VGND VGND VPWR VPWR _04005_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18023_ net1034 _01551_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_15235_ CPU.registerFile\[27\]\[22\] CPU.registerFile\[26\]\[22\] _03172_ VGND VGND
+ VPWR VPWR _03295_ sky130_fd_sc_hd__mux2_1
X_12447_ _07909_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15874__619 clknet_1_1__leaf__03682_ VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__inv_2
XFILLER_0_2_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13368__862 clknet_1_0__leaf__08369_ VGND VGND VPWR VPWR net918 sky130_fd_sc_hd__inv_2
XFILLER_0_140_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15166_ _03098_ _03225_ _03227_ _02903_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__a211o_1
X_12378_ _06643_ net1804 _07870_ VGND VGND VPWR VPWR _07873_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__03643_ _03643_ VGND VGND VPWR VPWR clknet_0__03643_ sky130_fd_sc_hd__clkbuf_16
X_11329_ _07237_ VGND VGND VPWR VPWR _07260_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15097_ CPU.registerFile\[17\]\[19\] _03036_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18925_ net699 _02445_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_13972__129 clknet_1_0__leaf__08481_ VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__inv_2
XFILLER_0_157_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18856_ net630 _02376_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_17807_ net887 _01369_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_18787_ net576 _02311_ VGND VGND VPWR VPWR CPU.aluReg\[17\] sky130_fd_sc_hd__dfxtp_1
X_15999_ _05689_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__buf_4
X_17738_ net823 _01304_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17669_ per_uart.uart0.rx_bitcount\[2\] per_uart.uart0.rx_bitcount\[1\] per_uart.uart0.rx_bitcount\[0\]
+ _04986_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__a31o_1
XFILLER_0_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09023_ CPU.rs2\[22\] _05246_ _05250_ VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold210 _02286_ VGND VGND VPWR VPWR net1507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold221 mapped_spi_flash.cmd_addr\[10\] VGND VGND VPWR VPWR net1518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 _08282_ VGND VGND VPWR VPWR net1529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold243 mapped_spi_flash.rcv_data\[23\] VGND VGND VPWR VPWR net1540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 mapped_spi_ram.rcv_data\[22\] VGND VGND VPWR VPWR net1551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold265 CPU.cycles\[27\] VGND VGND VPWR VPWR net1562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold276 CPU.state\[0\] VGND VGND VPWR VPWR net1573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold287 CPU.rs2\[28\] VGND VGND VPWR VPWR net1584 sky130_fd_sc_hd__dlygate4sd3_1
X_14090__235 clknet_1_1__leaf__08493_ VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__inv_2
X_09925_ _05318_ _05748_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__nor2_1
Xhold298 CPU.rs2\[26\] VGND VGND VPWR VPWR net1595 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ _05555_ _05326_ _05327_ _05526_ _05799_ VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__a2111oi_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _06125_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__clkbuf_1
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15669__466 clknet_1_1__leaf__03645_ VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__inv_2
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _06822_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__clkbuf_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _07462_ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__clkbuf_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13237__759 clknet_1_0__leaf__08342_ VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__inv_2
XFILLER_0_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10631_ _06784_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__clkbuf_1
X_10562_ net2010 _05873_ _06739_ VGND VGND VPWR VPWR _06747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12301_ mapped_spi_ram.rcv_data\[0\] _07786_ VGND VGND VPWR VPWR _07826_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10493_ net1938 _05873_ _06702_ VGND VGND VPWR VPWR _06710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15020_ CPU.registerFile\[30\]\[17\] CPU.registerFile\[31\]\[17\] _02887_ VGND VGND
+ VPWR VPWR _03085_ sky130_fd_sc_hd__mux2_1
X_12232_ mapped_spi_ram.rcv_data\[31\] _07787_ VGND VGND VPWR VPWR _07788_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12163_ net1471 _07714_ _07736_ _07737_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11114_ net1375 _07135_ VGND VGND VPWR VPWR _07137_ sky130_fd_sc_hd__or2_1
X_16971_ CPU.registerFile\[2\]\[23\] CPU.registerFile\[3\]\[23\] _04431_ VGND VGND
+ VPWR VPWR _04675_ sky130_fd_sc_hd__mux2_1
X_12094_ _07687_ net1312 _07675_ VGND VGND VPWR VPWR _07688_ sky130_fd_sc_hd__a21oi_4
X_18710_ net499 _02234_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[10\] sky130_fd_sc_hd__dfxtp_1
X_15922_ clknet_1_1__leaf__03686_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__buf_1
X_11045_ CPU.aluIn1\[6\] CPU.Bimm\[6\] _07082_ VGND VGND VPWR VPWR _07083_ sky130_fd_sc_hd__a21oi_1
X_13862__1220 clknet_1_1__leaf__08470_ VGND VGND VPWR VPWR net1276 sky130_fd_sc_hd__inv_2
XFILLER_0_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18641_ clknet_leaf_15_clk _02165_ VGND VGND VPWR VPWR CPU.rs2\[13\] sky130_fd_sc_hd__dfxtp_1
X_14804_ _08785_ _02872_ _02874_ _08870_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__a211o_1
X_18572_ net393 net29 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_12996_ _08201_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15784_ per_uart.uart0.enable16_counter\[15\] _08359_ VGND VGND VPWR VPWR _03658_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17523_ _05075_ _05025_ _06103_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__o21bai_1
X_11947_ _07604_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__clkbuf_1
X_14735_ CPU.registerFile\[30\]\[10\] CPU.registerFile\[31\]\[10\] _08645_ VGND VGND
+ VPWR VPWR _02807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ CPU.registerFile\[5\]\[8\] CPU.registerFile\[4\]\[8\] _08864_ VGND VGND VPWR
+ VPWR _02740_ sky130_fd_sc_hd__mux2_1
X_17454_ _05038_ _05039_ _05020_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__a21oi_1
X_11878_ _06607_ net1953 _07562_ VGND VGND VPWR VPWR _07568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16405_ CPU.registerFile\[28\]\[9\] CPU.registerFile\[29\]\[9\] _04122_ VGND VGND
+ VPWR VPWR _04123_ sky130_fd_sc_hd__mux2_1
X_10829_ CPU.aluIn1\[19\] _06910_ _06881_ VGND VGND VPWR VPWR _06911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17385_ per_uart.uart0.rxd_reg\[9\] _04992_ _04993_ per_uart.uart0.rxd_reg\[8\] VGND
+ VGND VPWR VPWR _05009_ sky130_fd_sc_hd__a22o_1
X_14597_ _08415_ _08833_ _08835_ _08420_ VGND VGND VPWR VPWR _08836_ sky130_fd_sc_hd__a211o_1
X_19124_ clknet_leaf_10_clk _02644_ VGND VGND VPWR VPWR CPU.PC\[6\] sky130_fd_sc_hd__dfxtp_2
X_16336_ CPU.registerFile\[10\]\[8\] CPU.registerFile\[11\]\[8\] _03931_ VGND VGND
+ VPWR VPWR _04055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16267_ CPU.registerFile\[0\]\[6\] _03828_ _03725_ _03987_ VGND VGND VPWR VPWR _03988_
+ sky130_fd_sc_hd__o211a_1
X_19055_ net797 _02575_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08481_ clknet_0__08481_ VGND VGND VPWR VPWR clknet_1_1__leaf__08481_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13479_ CPU.Bimm\[9\] _05783_ _08416_ VGND VGND VPWR VPWR _08431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15218_ _03027_ _03276_ _03278_ _03111_ VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__a211o_1
X_18006_ net1017 _01534_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16198_ CPU.registerFile\[20\]\[4\] CPU.registerFile\[21\]\[4\] _03883_ VGND VGND
+ VPWR VPWR _03921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15149_ CPU.registerFile\[30\]\[20\] CPU.registerFile\[31\]\[20\] _02887_ VGND VGND
+ VPWR VPWR _03211_ sky130_fd_sc_hd__mux2_1
X_15774__561 clknet_1_1__leaf__03655_ VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__inv_2
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13625__1006 clknet_1_1__leaf__08447_ VGND VGND VPWR VPWR net1062 sky130_fd_sc_hd__inv_2
XFILLER_0_77_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09710_ _05912_ _06051_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__nor2_1
X_18908_ net682 _02428_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_09641_ _05981_ _05984_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__nand2_1
X_18839_ clknet_leaf_7_clk _02363_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_09572_ CPU.PC\[23\] _05915_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15857__603 clknet_1_0__leaf__03681_ VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__inv_2
XFILLER_0_143_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09006_ CPU.aluIn1\[17\] _05345_ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13955__113 clknet_1_0__leaf__08480_ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__inv_2
X_09908_ _06204_ _06240_ _06241_ _05855_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__o22a_1
X_09839_ _05555_ _05526_ VGND VGND VPWR VPWR _06175_ sky130_fd_sc_hd__nand2_4
X_12850_ _08124_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__clkbuf_1
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _07527_ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__clkbuf_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _08086_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14520_ CPU.registerFile\[30\]\[5\] CPU.registerFile\[31\]\[5\] _08645_ VGND VGND
+ VPWR VPWR _08761_ sky130_fd_sc_hd__mux2_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13551__940 clknet_1_1__leaf__08439_ VGND VGND VPWR VPWR net996 sky130_fd_sc_hd__inv_2
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _06593_ net2202 _07490_ VGND VGND VPWR VPWR _07491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ CPU.registerFile\[13\]\[3\] CPU.registerFile\[12\]\[3\] _08693_ VGND VGND
+ VPWR VPWR _08694_ sky130_fd_sc_hd__mux2_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11663_ net2547 _07309_ _07453_ VGND VGND VPWR VPWR _07454_ sky130_fd_sc_hd__mux2_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13402_ _08379_ _06472_ _00000_ VGND VGND VPWR VPWR _08380_ sky130_fd_sc_hd__mux2_1
X_10614_ _05735_ _05736_ CPU.writeBack VGND VGND VPWR VPWR _06774_ sky130_fd_sc_hd__nand3b_4
X_17170_ CPU.registerFile\[16\]\[28\] _04656_ _06149_ _04868_ VGND VGND VPWR VPWR
+ _04869_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14382_ CPU.registerFile\[5\]\[1\] CPU.registerFile\[4\]\[1\] _08576_ VGND VGND VPWR
+ VPWR _08627_ sky130_fd_sc_hd__mux2_1
X_11594_ net2198 _07309_ _07416_ VGND VGND VPWR VPWR _07417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16121_ CPU.registerFile\[19\]\[2\] CPU.registerFile\[18\]\[2\] _03767_ VGND VGND
+ VPWR VPWR _03846_ sky130_fd_sc_hd__mux2_1
X_13333_ clknet_1_1__leaf__08341_ VGND VGND VPWR VPWR _08365_ sky130_fd_sc_hd__buf_1
XFILLER_0_106_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10545_ _05736_ _05740_ CPU.Bimm\[1\] VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__and3b_1
XFILLER_0_107_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16052_ net2661 _03566_ _03778_ _03390_ VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__o211a_1
X_10476_ _05735_ CPU.Bimm\[11\] _05740_ VGND VGND VPWR VPWR _06700_ sky130_fd_sc_hd__and3b_1
X_15003_ CPU.registerFile\[0\]\[16\] _02948_ _03068_ _02791_ VGND VGND VPWR VPWR _03069_
+ sky130_fd_sc_hd__o211a_1
X_12215_ mapped_spi_ram.snd_bitcount\[1\] mapped_spi_ram.snd_bitcount\[0\] mapped_spi_ram.snd_bitcount\[2\]
+ VGND VGND VPWR VPWR _07774_ sky130_fd_sc_hd__o21ai_1
X_13195_ net1502 _08307_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__xnor2_1
X_12146_ _07715_ _07725_ VGND VGND VPWR VPWR _07726_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12077_ mapped_spi_ram.state\[2\] net1301 VGND VGND VPWR VPWR _07676_ sky130_fd_sc_hd__nor2_1
X_16954_ _04367_ _04655_ _04658_ _04410_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__a211o_1
X_11028_ _07001_ VGND VGND VPWR VPWR _07069_ sky130_fd_sc_hd__clkbuf_4
X_16885_ _04503_ _04588_ _04590_ _04509_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__a211o_1
XFILLER_0_154_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18624_ net445 _02148_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18555_ net376 _02079_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_12979_ net1961 _07332_ _08192_ VGND VGND VPWR VPWR _08193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17506_ _08335_ _06189_ _05073_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_144_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14718_ _08549_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18486_ net307 _02010_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17437_ _08311_ _06467_ _05025_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__nor3_1
XFILLER_0_145_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14649_ _08808_ _08809_ CPU.registerFile\[25\]\[8\] VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_16 _04160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_27 _04838_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 _07919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_49 clknet_1_1__leaf__08506_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17368_ _04996_ _04997_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19107_ net90 _02627_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16319_ _03749_ _03751_ CPU.registerFile\[25\]\[7\] VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19038_ net780 _02558_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08464_ clknet_0__08464_ VGND VGND VPWR VPWR clknet_1_1__leaf__08464_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15698__492 clknet_1_0__leaf__03648_ VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__inv_2
XFILLER_0_11_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__08495_ _08495_ VGND VGND VPWR VPWR clknet_0__08495_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15852__599 clknet_1_1__leaf__03680_ VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__inv_2
XFILLER_0_128_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09624_ CPU.PC\[7\] CPU.Bimm\[7\] _05913_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__and3_1
X_09555_ _05488_ _05898_ _05491_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09486_ _05793_ _05810_ VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14022__173 clknet_1_0__leaf__08487_ VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__inv_2
X_10330_ _05872_ VGND VGND VPWR VPWR _06611_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14096__241 clknet_1_0__leaf__08493_ VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__inv_2
XFILLER_0_103_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13581__966 clknet_1_0__leaf__08443_ VGND VGND VPWR VPWR net1022 sky130_fd_sc_hd__inv_2
X_10261_ _06570_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__clkbuf_1
X_12000_ _06661_ net2472 _07597_ VGND VGND VPWR VPWR _07632_ sky130_fd_sc_hd__mux2_1
X_10192_ _06140_ _06390_ _06513_ _06176_ VGND VGND VPWR VPWR _06514_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12902_ _05853_ net2381 _08145_ VGND VGND VPWR VPWR _08152_ sky130_fd_sc_hd__mux2_1
X_16670_ CPU.registerFile\[13\]\[16\] _04380_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15610__413 clknet_1_1__leaf__03639_ VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__inv_2
XFILLER_0_88_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__08484_ clknet_0__08484_ VGND VGND VPWR VPWR clknet_1_0__leaf__08484_
+ sky130_fd_sc_hd__clkbuf_16
X_12833_ _08115_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__clkbuf_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ net161 _01868_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _06620_ net2159 _08076_ VGND VGND VPWR VPWR _08078_ sky130_fd_sc_hd__mux2_1
X_15552_ CPU.registerFile\[19\]\[31\] CPU.registerFile\[18\]\[31\] _06456_ VGND VGND
+ VPWR VPWR _03603_ sky130_fd_sc_hd__mux2_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13624__1005 clknet_1_0__leaf__08447_ VGND VGND VPWR VPWR net1061 sky130_fd_sc_hd__inv_2
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ net2576 _07364_ _07475_ VGND VGND VPWR VPWR _07481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14503_ _08585_ _08586_ CPU.registerFile\[1\]\[4\] VGND VGND VPWR VPWR _08745_ sky130_fd_sc_hd__a21o_1
XFILLER_0_154_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18271_ net1282 _01799_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_15483_ CPU.registerFile\[21\]\[29\] _02752_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__or2_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _08041_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__clkbuf_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17222_ _04917_ _04918_ _03769_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__mux2_1
X_13332__831 clknet_1_1__leaf__08364_ VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__inv_2
XFILLER_0_154_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11646_ net2450 _07364_ _07438_ VGND VGND VPWR VPWR _07444_ sky130_fd_sc_hd__mux2_1
X_14434_ _08415_ _08674_ _08676_ _08420_ VGND VGND VPWR VPWR _08677_ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17153_ CPU.registerFile\[0\]\[28\] _04637_ _03741_ _04851_ VGND VGND VPWR VPWR _04852_
+ sky130_fd_sc_hd__o211a_1
X_14365_ _08607_ _08608_ _08609_ VGND VGND VPWR VPWR _08610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11577_ net1687 _07364_ _07401_ VGND VGND VPWR VPWR _07407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16104_ _03726_ _03727_ CPU.registerFile\[1\]\[2\] VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17084_ _04502_ _04772_ _04776_ _04784_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__a31o_2
X_10528_ _06728_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__clkbuf_1
Xhold809 CPU.registerFile\[12\]\[9\] VGND VGND VPWR VPWR net2106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14296_ _08537_ _08539_ _08541_ VGND VGND VPWR VPWR _08542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16035_ CPU.registerFile\[20\]\[0\] CPU.registerFile\[21\]\[0\] _03761_ VGND VGND
+ VPWR VPWR _03762_ sky130_fd_sc_hd__mux2_1
X_10459_ _06691_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13178_ net1565 _08297_ VGND VGND VPWR VPWR _08300_ sky130_fd_sc_hd__nor2_1
X_12129_ net1424 _07693_ _07712_ _07713_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__o211a_1
X_17986_ net997 _01514_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_16937_ _04502_ _04628_ _04632_ _04641_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__a31o_2
XFILLER_0_79_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16868_ CPU.registerFile\[22\]\[20\] CPU.registerFile\[23\]\[20\] _04362_ VGND VGND
+ VPWR VPWR _04575_ sky130_fd_sc_hd__mux2_1
X_18607_ net428 _02131_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_16799_ CPU.registerFile\[9\]\[19\] _04460_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__or2_1
X_09340_ _05689_ _05690_ _05691_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__a21o_1
X_18538_ net359 _02062_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09271_ _05621_ _05616_ _05622_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__o21ba_1
X_18469_ net290 _01993_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_562 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08447_ clknet_0__08447_ VGND VGND VPWR VPWR clknet_1_1__leaf__08447_
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0__08478_ _08478_ VGND VGND VPWR VPWR clknet_0__08478_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08986_ _05337_ _05331_ _05326_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__a21oi_1
X_14210__343 clknet_1_0__leaf__08505_ VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__inv_2
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09607_ CPU.PC\[4\] _05950_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__or2_1
X_09538_ CPU.PC\[4\] CPU.PC\[3\] CPU.PC\[2\] VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09469_ _05812_ _05816_ _05794_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11500_ net1679 _07362_ _07354_ VGND VGND VPWR VPWR _07363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12480_ net2326 _07324_ _07920_ VGND VGND VPWR VPWR _07927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11431_ _05785_ VGND VGND VPWR VPWR _07316_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11362_ net1828 _05805_ _07274_ VGND VGND VPWR VPWR _07278_ sky130_fd_sc_hd__mux2_1
X_13101_ mapped_spi_flash.rbusy mapped_spi_ram.rbusy CPU.state\[2\] VGND VGND VPWR
+ VPWR _08257_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10313_ _06599_ net1840 _06597_ VGND VGND VPWR VPWR _06600_ sky130_fd_sc_hd__mux2_1
X_13926__87 clknet_1_1__leaf__08477_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__inv_2
X_11293_ _07241_ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_946 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13032_ CPU.registerFile\[4\]\[28\] net1402 _08217_ VGND VGND VPWR VPWR _08221_ sky130_fd_sc_hd__mux2_1
X_10244_ _06561_ VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15835__583 clknet_1_0__leaf__03679_ VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__inv_2
X_13362__857 clknet_1_1__leaf__08368_ VGND VGND VPWR VPWR net913 sky130_fd_sc_hd__inv_2
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17840_ net920 _01402_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_10175_ _05281_ _05440_ VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__xnor2_1
X_17771_ net851 _01333_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_14983_ _06058_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__clkbuf_4
X_16722_ CPU.registerFile\[2\]\[17\] CPU.registerFile\[3\]\[17\] _04431_ VGND VGND
+ VPWR VPWR _04432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16653_ _03741_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__buf_4
Xclkbuf_1_0__f__08467_ clknet_0__08467_ VGND VGND VPWR VPWR clknet_1_0__leaf__08467_
+ sky130_fd_sc_hd__clkbuf_16
X_12816_ CPU.aluShamt\[1\] CPU.aluShamt\[0\] VGND VGND VPWR VPWR _08106_ sky130_fd_sc_hd__and2_1
X_16584_ CPU.registerFile\[10\]\[14\] CPU.registerFile\[11\]\[14\] _03931_ VGND VGND
+ VPWR VPWR _04297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18323_ net144 _01851_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_15535_ CPU.registerFile\[10\]\[30\] CPU.registerFile\[11\]\[30\] _08522_ VGND VGND
+ VPWR VPWR _03587_ sky130_fd_sc_hd__mux2_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _06603_ net2310 _08065_ VGND VGND VPWR VPWR _08069_ sky130_fd_sc_hd__mux2_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18254_ net1265 _01782_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15466_ _08533_ _03515_ _03519_ _03188_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__o211a_1
X_12678_ _08032_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17205_ _04579_ _04580_ CPU.registerFile\[17\]\[29\] VGND VGND VPWR VPWR _04903_
+ sky130_fd_sc_hd__a21o_1
X_11629_ net2229 _07347_ _07427_ VGND VGND VPWR VPWR _07435_ sky130_fd_sc_hd__mux2_1
X_14417_ _08418_ VGND VGND VPWR VPWR _08661_ sky130_fd_sc_hd__buf_2
XFILLER_0_127_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18185_ net1196 _01713_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[24\] sky130_fd_sc_hd__dfxtp_1
X_15397_ _03451_ _03452_ _08562_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17136_ _04574_ _04831_ _04835_ _04584_ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14348_ _05861_ VGND VGND VPWR VPWR _08594_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold606 CPU.registerFile\[2\]\[19\] VGND VGND VPWR VPWR net1903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 CPU.registerFile\[11\]\[8\] VGND VGND VPWR VPWR net1914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 CPU.registerFile\[10\]\[16\] VGND VGND VPWR VPWR net1925 sky130_fd_sc_hd__dlygate4sd3_1
X_15918__658 clknet_1_1__leaf__03687_ VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__inv_2
Xhold639 CPU.registerFile\[15\]\[23\] VGND VGND VPWR VPWR net1936 sky130_fd_sc_hd__dlygate4sd3_1
X_14279_ _08408_ VGND VGND VPWR VPWR _08525_ sky130_fd_sc_hd__clkbuf_8
X_17067_ net2591 _04458_ _04768_ _04663_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16018_ _03744_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__buf_4
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1306 CPU.PC\[6\] VGND VGND VPWR VPWR net2603 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1317 CPU.registerFile\[3\]\[2\] VGND VGND VPWR VPWR net2614 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ net980 _01497_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold1328 _02690_ VGND VGND VPWR VPWR net2625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1339 CPU.registerFile\[25\]\[31\] VGND VGND VPWR VPWR net2636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13339__837 clknet_1_1__leaf__08365_ VGND VGND VPWR VPWR net893 sky130_fd_sc_hd__inv_2
XFILLER_0_149_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09323_ _05564_ _05673_ _05674_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09254_ CPU.aluIn1\[12\] _05543_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09185_ CPU.aluIn1\[31\] _05525_ _05533_ _05536_ CPU.aluReg\[31\] VGND VGND VPWR
+ VPWR _05537_ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__04981_ clknet_0__04981_ VGND VGND VPWR VPWR clknet_1_0__leaf__04981_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13623__1004 clknet_1_0__leaf__08447_ VGND VGND VPWR VPWR net1060 sky130_fd_sc_hd__inv_2
X_14134__274 clknet_1_0__leaf__08498_ VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__inv_2
X_08969_ _05261_ _05311_ _05313_ _05315_ _05320_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__o311a_2
X_11980_ _06641_ net2414 _07620_ VGND VGND VPWR VPWR _07622_ sky130_fd_sc_hd__mux2_1
X_10931_ _06973_ _06990_ VGND VGND VPWR VPWR _06991_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10862_ CPU.aluReg\[12\] CPU.aluReg\[10\] _06906_ VGND VGND VPWR VPWR _06936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12601_ net2428 _07376_ _07956_ VGND VGND VPWR VPWR _07991_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10793_ _06883_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__clkbuf_1
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12532_ net2367 _07376_ _07919_ VGND VGND VPWR VPWR _07954_ sky130_fd_sc_hd__mux2_1
X_15320_ _03098_ _03375_ _03377_ _03307_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__a211o_1
X_15722__514 clknet_1_0__leaf__03650_ VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__inv_2
XFILLER_0_38_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12463_ _07917_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__clkbuf_1
X_15251_ CPU.registerFile\[5\]\[22\] CPU.registerFile\[4\]\[22\] _03105_ VGND VGND
+ VPWR VPWR _03311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17353__13 clknet_1_0__leaf__04985_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__inv_2
X_11414_ net1787 _06486_ _07296_ VGND VGND VPWR VPWR _07305_ sky130_fd_sc_hd__mux2_1
X_15182_ _03155_ _03221_ _03242_ _03243_ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__a211o_1
X_12394_ _06659_ net2321 _07847_ VGND VGND VPWR VPWR _07881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11345_ _07268_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14064_ clknet_1_1__leaf__08484_ VGND VGND VPWR VPWR _08491_ sky130_fd_sc_hd__buf_1
X_18941_ net715 _02461_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_11276_ _07231_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__clkbuf_1
X_13015_ _08211_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__clkbuf_1
X_10227_ _06521_ VGND VGND VPWR VPWR _06548_ sky130_fd_sc_hd__inv_2
X_18872_ net646 _02392_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_17823_ net903 _01385_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_10158_ _05269_ _05532_ _05535_ CPU.aluReg\[3\] _06481_ VGND VGND VPWR VPWR _06482_
+ sky130_fd_sc_hd__a221o_1
Xhold3 _01683_ VGND VGND VPWR VPWR net1300 sky130_fd_sc_hd__dlygate4sd3_1
X_17754_ net839 _01320_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_14966_ _03022_ _03032_ _02837_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__o21a_2
X_10089_ mapped_spi_ram.rcv_data\[29\] _05857_ VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_535 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16705_ CPU.registerFile\[10\]\[17\] CPU.registerFile\[11\]\[17\] _04335_ VGND VGND
+ VPWR VPWR _04415_ sky130_fd_sc_hd__mux2_1
X_17685_ CPU.mem_wdata\[2\] per_uart.uart_ctrl\[2\] _05211_ VGND VGND VPWR VPWR _05214_
+ sky130_fd_sc_hd__mux2_1
X_14897_ CPU.registerFile\[30\]\[14\] CPU.registerFile\[31\]\[14\] _02887_ VGND VGND
+ VPWR VPWR _02965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16636_ CPU.registerFile\[2\]\[15\] CPU.registerFile\[3\]\[15\] _04027_ VGND VGND
+ VPWR VPWR _04348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16567_ CPU.registerFile\[27\]\[13\] CPU.registerFile\[26\]\[13\] _04242_ VGND VGND
+ VPWR VPWR _04281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18306_ net127 _01834_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_15518_ _08521_ _03567_ _03569_ _08590_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__a211o_1
X_16498_ CPU.registerFile\[19\]\[11\] CPU.registerFile\[18\]\[11\] _03923_ VGND VGND
+ VPWR VPWR _04214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18237_ net1248 _01765_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_127_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15449_ _08581_ _03500_ _03502_ _08535_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18168_ net1179 _01696_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold403 CPU.registerFile\[5\]\[29\] VGND VGND VPWR VPWR net1700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 CPU.registerFile\[10\]\[27\] VGND VGND VPWR VPWR net1711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17119_ _03757_ _04814_ _04818_ _04476_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__o211a_1
Xhold425 CPU.registerFile\[10\]\[23\] VGND VGND VPWR VPWR net1722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 CPU.registerFile\[15\]\[2\] VGND VGND VPWR VPWR net1733 sky130_fd_sc_hd__dlygate4sd3_1
X_18099_ net1110 _01627_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold447 CPU.registerFile\[27\]\[30\] VGND VGND VPWR VPWR net1744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 CPU.registerFile\[19\]\[5\] VGND VGND VPWR VPWR net1755 sky130_fd_sc_hd__dlygate4sd3_1
X_13905__68 clknet_1_0__leaf__08475_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__inv_2
Xhold469 per_uart.uart0.rx_count16\[1\] VGND VGND VPWR VPWR net1766 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ _05461_ _06272_ _05310_ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__a21o_1
Xclkbuf_1_1__f__03688_ clknet_0__03688_ VGND VGND VPWR VPWR clknet_1_1__leaf__03688_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _06204_ _06205_ _06206_ CPU.Jimm\[13\] VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__o22a_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 CPU.registerFile\[31\]\[7\] VGND VGND VPWR VPWR net2400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 CPU.registerFile\[8\]\[9\] VGND VGND VPWR VPWR net2411 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1125 CPU.registerFile\[14\]\[16\] VGND VGND VPWR VPWR net2422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 CPU.aluShamt\[3\] VGND VGND VPWR VPWR net2433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1147 CPU.registerFile\[9\]\[16\] VGND VGND VPWR VPWR net2444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 CPU.registerFile\[14\]\[23\] VGND VGND VPWR VPWR net2455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 CPU.registerFile\[24\]\[24\] VGND VGND VPWR VPWR net2466 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09306_ _05642_ _05651_ _05657_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__and3b_1
XFILLER_0_64_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09237_ _05587_ _05588_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09168_ CPU.Jimm\[13\] CPU.Jimm\[12\] VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__nor2_8
XFILLER_0_161_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09099_ _05450_ _05265_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__nor2_2
XFILLER_0_160_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11130_ net1416 _07133_ _07145_ _07138_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold970 CPU.registerFile\[30\]\[16\] VGND VGND VPWR VPWR net2267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 CPU.registerFile\[22\]\[10\] VGND VGND VPWR VPWR net2278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold992 CPU.registerFile\[29\]\[25\] VGND VGND VPWR VPWR net2289 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ CPU.PC\[5\] _07031_ _07095_ _07096_ _05703_ VGND VGND VPWR VPWR _07097_ sky130_fd_sc_hd__o221a_1
X_10012_ net1384 _05762_ _05717_ per_uart.rx_avail _06340_ VGND VGND VPWR VPWR _06341_
+ sky130_fd_sc_hd__a221o_1
X_14820_ _02888_ _02889_ _02851_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__mux2_1
X_17405__28 clknet_1_1__leaf__05013_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__inv_2
X_14751_ CPU.registerFile\[8\]\[10\] _08776_ _02822_ _08622_ VGND VGND VPWR VPWR _02823_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11963_ _06624_ net2128 _07609_ VGND VGND VPWR VPWR _07613_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15947__684 clknet_1_0__leaf__03690_ VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__inv_2
X_10914_ mapped_spi_flash.state\[1\] VGND VGND VPWR VPWR _06976_ sky130_fd_sc_hd__inv_2
X_17470_ _07001_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__buf_2
X_11894_ _07576_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__clkbuf_1
X_14682_ _08526_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16421_ _04129_ _04137_ _04138_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__o21a_1
X_10845_ _06923_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19140_ clknet_leaf_15_clk _02660_ VGND VGND VPWR VPWR CPU.PC\[22\] sky130_fd_sc_hd__dfxtp_2
X_16352_ _03943_ _04067_ _04070_ _03730_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10776_ net2607 _06866_ _06869_ VGND VGND VPWR VPWR _06870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15303_ CPU.registerFile\[20\]\[24\] _03080_ _03360_ _03082_ VGND VGND VPWR VPWR
+ _03361_ sky130_fd_sc_hd__o211a_1
X_12515_ _07945_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19071_ net63 _02591_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_16283_ _03770_ _03771_ CPU.registerFile\[17\]\[6\] VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18022_ net1033 _01550_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_12446_ net1834 _07358_ _07906_ VGND VGND VPWR VPWR _07909_ sky130_fd_sc_hd__mux2_1
X_15234_ _03292_ _03293_ _03255_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12377_ _07872_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__clkbuf_1
X_15165_ CPU.registerFile\[8\]\[20\] _03018_ _03226_ _02864_ VGND VGND VPWR VPWR _03227_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11328_ _07259_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__03642_ _03642_ VGND VGND VPWR VPWR clknet_0__03642_ sky130_fd_sc_hd__clkbuf_16
X_15096_ _08526_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18924_ net698 _02444_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_11259_ _07222_ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__clkbuf_1
X_15692__487 clknet_1_0__leaf__03647_ VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__inv_2
X_17334__746 clknet_1_0__leaf__04983_ VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__inv_2
X_18855_ net629 _02375_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_17806_ net886 _01368_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_18786_ net575 _02310_ VGND VGND VPWR VPWR CPU.aluReg\[16\] sky130_fd_sc_hd__dfxtp_1
X_15998_ _06148_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__buf_4
X_17737_ net822 _01303_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_14949_ _03014_ _03015_ _02937_ VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__mux2_1
X_17668_ net1631 VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16619_ _04170_ _04326_ _04331_ _04180_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17599_ _05123_ _05121_ _05124_ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__or3b_1
XFILLER_0_18_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13622__1003 clknet_1_0__leaf__08447_ VGND VGND VPWR VPWR net1059 sky130_fd_sc_hd__inv_2
XFILLER_0_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09022_ _05372_ _05373_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_31_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold200 mapped_spi_flash.cmd_addr\[11\] VGND VGND VPWR VPWR net1497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 per_uart.uart0.enable16_counter\[6\] VGND VGND VPWR VPWR net1508 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold222 mapped_spi_ram.cmd_addr\[14\] VGND VGND VPWR VPWR net1519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold233 mapped_spi_flash.cmd_addr\[24\] VGND VGND VPWR VPWR net1530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 per_uart.uart0.enable16_counter\[12\] VGND VGND VPWR VPWR net1541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 mapped_spi_flash.cmd_addr\[17\] VGND VGND VPWR VPWR net1552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 mapped_spi_flash.cmd_addr\[0\] VGND VGND VPWR VPWR net1563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 CPU.rs2\[23\] VGND VGND VPWR VPWR net1574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 per_uart.uart0.tx_bitcount\[3\] VGND VGND VPWR VPWR net1585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 per_uart.uart0.enable16_counter\[7\] VGND VGND VPWR VPWR net1596 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ _05427_ _06252_ _06256_ _05517_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ _05427_ _06185_ _06186_ _06190_ _05517_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__o311a_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09786_ net2356 _06124_ _06055_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__mux2_1
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14246__375 clknet_1_0__leaf__08509_ VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__inv_2
XFILLER_0_138_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ net2553 _05853_ _06777_ VGND VGND VPWR VPWR _06784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10561_ _06746_ VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12300_ net1319 _07784_ _07825_ _07822_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13280_ net1500 _08360_ _06856_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__o21ai_1
X_10492_ _06709_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12231_ _07786_ VGND VGND VPWR VPWR _07787_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_133_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12162_ _07163_ VGND VGND VPWR VPWR _07737_ sky130_fd_sc_hd__buf_2
XFILLER_0_20_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11113_ net1375 _07133_ _07136_ _07069_ VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__o211a_1
X_16970_ _04672_ _04673_ _04557_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__mux2_1
X_12093_ net8 VGND VGND VPWR VPWR _07687_ sky130_fd_sc_hd__inv_2
X_11044_ _05570_ _05592_ VGND VGND VPWR VPWR _07082_ sky130_fd_sc_hd__nor2_1
X_18640_ clknet_leaf_15_clk _02164_ VGND VGND VPWR VPWR CPU.rs2\[12\] sky130_fd_sc_hd__dfxtp_1
X_14803_ CPU.registerFile\[0\]\[11\] _08706_ _02873_ _02791_ VGND VGND VPWR VPWR _02874_
+ sky130_fd_sc_hd__o211a_1
X_18571_ net392 net28 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_15783_ net1514 net1500 VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12995_ net1942 _07349_ _08192_ VGND VGND VPWR VPWR _08201_ sky130_fd_sc_hd__mux2_1
X_17522_ _05069_ CPU.PC\[18\] _05094_ _05095_ _05053_ VGND VGND VPWR VPWR _02656_
+ sky130_fd_sc_hd__o221a_1
X_14734_ _08837_ _02803_ _02805_ _08802_ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__a211o_1
X_15728__520 clknet_1_1__leaf__03650_ VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__inv_2
X_11946_ _06607_ net2449 _07598_ VGND VGND VPWR VPWR _07604_ sky130_fd_sc_hd__mux2_1
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15880__624 clknet_1_1__leaf__03683_ VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__inv_2
XFILLER_0_143_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17453_ _08311_ _06401_ _08331_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__or3_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14665_ CPU.registerFile\[6\]\[8\] CPU.registerFile\[7\]\[8\] _08740_ VGND VGND VPWR
+ VPWR _02739_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _07567_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16404_ _06171_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__buf_4
X_10828_ CPU.aluReg\[20\] CPU.aluReg\[18\] _06906_ VGND VGND VPWR VPWR _06910_ sky130_fd_sc_hd__mux2_1
X_17384_ _05008_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__clkbuf_1
X_14596_ CPU.registerFile\[16\]\[7\] _08412_ _08834_ _06037_ VGND VGND VPWR VPWR _08835_
+ sky130_fd_sc_hd__o211a_1
X_19123_ clknet_leaf_2_clk _02643_ VGND VGND VPWR VPWR CPU.PC\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16335_ _08513_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__buf_2
XFILLER_0_125_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10759_ _06854_ VGND VGND VPWR VPWR _06855_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_137_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19054_ net796 _02574_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__08480_ clknet_0__08480_ VGND VGND VPWR VPWR clknet_1_1__leaf__08480_
+ sky130_fd_sc_hd__clkbuf_16
X_16266_ _03985_ _03986_ CPU.registerFile\[1\]\[6\] VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__a21o_1
X_13478_ _08430_ VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18005_ net1016 _01533_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15217_ CPU.registerFile\[0\]\[21\] _02948_ _03277_ _03195_ VGND VGND VPWR VPWR _03278_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12429_ net1864 _07341_ _07895_ VGND VGND VPWR VPWR _07900_ sky130_fd_sc_hd__mux2_1
X_16197_ CPU.registerFile\[22\]\[4\] CPU.registerFile\[23\]\[4\] _03759_ VGND VGND
+ VPWR VPWR _03920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15148_ _03078_ _03207_ _03209_ _03043_ VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__a211o_1
X_15700__494 clknet_1_0__leaf__03648_ VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__inv_2
X_15079_ _03133_ _03136_ _03142_ _02784_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__o211a_1
X_18907_ net681 _02427_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09640_ CPU.PC\[13\] _05938_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__nand2_1
X_18838_ clknet_leaf_6_clk _02362_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_09571_ CPU.Iimm\[3\] _05545_ _05914_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__mux2_1
X_18769_ net558 _02293_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_830 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09005_ _05356_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13799__1162 clknet_1_1__leaf__08465_ VGND VGND VPWR VPWR net1218 sky130_fd_sc_hd__inv_2
X_09907_ _06203_ _05783_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__or2_1
X_13243__764 clknet_1_0__leaf__08343_ VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__inv_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09838_ _05692_ _05694_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__nand2_1
X_18569__26 VGND VGND VPWR VPWR _18569__26/HI net26 sky130_fd_sc_hd__conb_1
X_09769_ mapped_spi_ram.rcv_data\[10\] _05858_ _05860_ net1419 VGND VGND VPWR VPWR
+ _06108_ sky130_fd_sc_hd__a22oi_4
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ net1803 _07309_ _07526_ VGND VGND VPWR VPWR _07527_ sky130_fd_sc_hd__mux2_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12780_ _06636_ net2566 _08076_ VGND VGND VPWR VPWR _08086_ sky130_fd_sc_hd__mux2_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _07489_ VGND VGND VPWR VPWR _07490_ sky130_fd_sc_hd__buf_4
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14450_ _06061_ VGND VGND VPWR VPWR _08693_ sky130_fd_sc_hd__buf_4
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11662_ _07452_ VGND VGND VPWR VPWR _07453_ sky130_fd_sc_hd__buf_4
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13401_ _08310_ VGND VGND VPWR VPWR _08379_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10613_ _06773_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__clkbuf_1
X_11593_ _07415_ VGND VGND VPWR VPWR _07416_ sky130_fd_sc_hd__buf_4
X_14381_ CPU.registerFile\[6\]\[1\] CPU.registerFile\[7\]\[1\] _08522_ VGND VGND VPWR
+ VPWR _08626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16120_ _03843_ _03844_ _03763_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10544_ _06736_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16051_ _03692_ _03734_ _03777_ _03601_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__a211o_1
XFILLER_0_161_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10475_ _06699_ VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15002_ _02831_ _02832_ CPU.registerFile\[1\]\[16\] VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12214_ _07773_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13194_ _08309_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__clkbuf_1
X_14073__220 clknet_1_1__leaf__08491_ VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__inv_2
X_12145_ mapped_spi_ram.cmd_addr\[16\] _07061_ _07724_ VGND VGND VPWR VPWR _07725_
+ sky130_fd_sc_hd__mux2_1
X_12076_ _07672_ _07674_ VGND VGND VPWR VPWR _07675_ sky130_fd_sc_hd__nor2_2
X_16953_ CPU.registerFile\[16\]\[22\] _04656_ _04494_ _04657_ VGND VGND VPWR VPWR
+ _04658_ sky130_fd_sc_hd__o211a_1
X_13621__1002 clknet_1_0__leaf__08447_ VGND VGND VPWR VPWR net1058 sky130_fd_sc_hd__inv_2
X_11027_ _07048_ _07067_ VGND VGND VPWR VPWR _07068_ sky130_fd_sc_hd__or2_1
X_16884_ CPU.registerFile\[8\]\[21\] _04505_ _04506_ _04589_ VGND VGND VPWR VPWR _04590_
+ sky130_fd_sc_hd__o211a_1
X_18623_ net444 _02147_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18554_ net375 _02078_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12978_ _08180_ VGND VGND VPWR VPWR _08192_ sky130_fd_sc_hd__clkbuf_4
X_17505_ _05080_ _05081_ _05058_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__a21oi_1
X_14717_ _08585_ _08586_ CPU.registerFile\[1\]\[9\] VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__a21o_1
X_18485_ net306 _02009_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_11929_ _07594_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15697_ clknet_1_1__leaf__03643_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__buf_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17436_ net13 VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18583__40 VGND VGND VPWR VPWR _18583__40/HI net40 sky130_fd_sc_hd__conb_1
X_14648_ CPU.registerFile\[27\]\[8\] CPU.registerFile\[26\]\[8\] _06063_ VGND VGND
+ VPWR VPWR _02722_ sky130_fd_sc_hd__mux2_1
XANTENNA_17 _04360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_28 _04943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17367_ per_uart.uart0.rxd_reg\[3\] _04992_ _04993_ per_uart.uart0.rxd_reg\[2\] VGND
+ VGND VPWR VPWR _04997_ sky130_fd_sc_hd__a22o_1
XANTENNA_39 _08419_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14579_ _08567_ _08569_ CPU.registerFile\[9\]\[6\] VGND VGND VPWR VPWR _08819_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19106_ net89 _02626_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_16318_ CPU.registerFile\[27\]\[7\] CPU.registerFile\[26\]\[7\] _03837_ VGND VGND
+ VPWR VPWR _04038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19037_ net779 _02557_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__08463_ clknet_0__08463_ VGND VGND VPWR VPWR clknet_1_1__leaf__08463_
+ sky130_fd_sc_hd__clkbuf_16
X_16249_ _05284_ _03566_ _03970_ _03855_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__08494_ _08494_ VGND VGND VPWR VPWR clknet_0__08494_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09623_ _05948_ _05965_ _05966_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__a21o_1
X_13535__925 clknet_1_0__leaf__08438_ VGND VGND VPWR VPWR net981 sky130_fd_sc_hd__inv_2
X_09554_ _05366_ _05486_ _05490_ VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09485_ _05831_ _05808_ _05404_ _05809_ VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10260_ net1684 _06054_ _06569_ VGND VGND VPWR VPWR _06570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10191_ net1578 _05859_ _05719_ per_uart.rx_data\[1\] _06512_ VGND VGND VPWR VPWR
+ _06513_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12901_ _08151_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__08483_ clknet_0__08483_ VGND VGND VPWR VPWR clknet_1_0__leaf__08483_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _05839_ net2319 _08109_ VGND VGND VPWR VPWR _08115_ sky130_fd_sc_hd__mux2_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ net1666 _03566_ _03602_ _03390_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _08077_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__clkbuf_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13719__1091 clknet_1_1__leaf__08456_ VGND VGND VPWR VPWR net1147 sky130_fd_sc_hd__inv_2
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ CPU.registerFile\[2\]\[4\] CPU.registerFile\[3\]\[4\] _08629_ VGND VGND VPWR
+ VPWR _08744_ sky130_fd_sc_hd__mux2_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _07480_ VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__clkbuf_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ net1281 _01798_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ CPU.registerFile\[22\]\[29\] CPU.registerFile\[23\]\[29\] _08584_ VGND VGND
+ VPWR VPWR _03535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _06617_ net2530 _08040_ VGND VGND VPWR VPWR _08041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17221_ CPU.registerFile\[5\]\[30\] CPU.registerFile\[4\]\[30\] _03697_ VGND VGND
+ VPWR VPWR _04918_ sky130_fd_sc_hd__mux2_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ CPU.registerFile\[16\]\[3\] _08412_ _08675_ _06037_ VGND VGND VPWR VPWR _08676_
+ sky130_fd_sc_hd__o211a_1
X_11645_ _07443_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__clkbuf_1
X_14105__249 clknet_1_1__leaf__08494_ VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__inv_2
XFILLER_0_71_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17152_ _03748_ _03750_ CPU.registerFile\[1\]\[28\] VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__a21o_1
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14364_ _08549_ VGND VGND VPWR VPWR _08609_ sky130_fd_sc_hd__buf_4
X_11576_ _07406_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_922 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16103_ _06172_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__clkbuf_4
X_17083_ _03757_ _04779_ _04783_ _04476_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10527_ net2272 _06361_ _06724_ VGND VGND VPWR VPWR _06728_ sky130_fd_sc_hd__mux2_1
X_14295_ _08540_ VGND VGND VPWR VPWR _08541_ sky130_fd_sc_hd__clkbuf_8
X_16034_ _03736_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__buf_4
X_10458_ _06645_ net2327 _06687_ VGND VGND VPWR VPWR _06691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10389_ _06439_ VGND VGND VPWR VPWR _06651_ sky130_fd_sc_hd__clkbuf_8
X_13177_ CPU.cycles\[24\] _08297_ VGND VGND VPWR VPWR _08299_ sky130_fd_sc_hd__and2_1
X_12128_ _07163_ VGND VGND VPWR VPWR _07713_ sky130_fd_sc_hd__buf_2
X_17985_ net996 _01513_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_16936_ _04305_ _04635_ _04640_ _04476_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__o211a_1
X_12059_ CPU.registerFile\[24\]\[5\] _07366_ _07657_ VGND VGND VPWR VPWR _07664_ sky130_fd_sc_hd__mux2_1
X_15886__630 clknet_1_0__leaf__03683_ VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__inv_2
X_16867_ _03713_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__clkbuf_4
X_18606_ net427 _02130_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_15818_ _03677_ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__clkbuf_1
X_16798_ _06149_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__clkbuf_4
X_18537_ net358 _02061_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13984__140 clknet_1_0__leaf__08482_ VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__inv_2
X_09270_ CPU.aluIn1\[15\] CPU.aluIn1\[14\] CPU.aluIn1\[13\] CPU.aluIn1\[12\] _05543_
+ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__o41a_1
X_18468_ net289 _01992_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18399_ net220 _01927_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08446_ clknet_0__08446_ VGND VGND VPWR VPWR clknet_1_1__leaf__08446_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08477_ _08477_ VGND VGND VPWR VPWR clknet_0__08477_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08985_ CPU.aluIn1\[15\] _05325_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__or2_1
X_09606_ CPU.Iimm\[4\] _05547_ _05922_ _05739_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13879__1235 clknet_1_0__leaf__08472_ VGND VGND VPWR VPWR net1291 sky130_fd_sc_hd__inv_2
XFILLER_0_97_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09537_ _05547_ _05880_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__nor2_2
XFILLER_0_149_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13316__816 clknet_1_1__leaf__08363_ VGND VGND VPWR VPWR net872 sky130_fd_sc_hd__inv_2
X_09468_ _05396_ _05815_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15941__679 clknet_1_0__leaf__03689_ VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__inv_2
XFILLER_0_53_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09399_ _05412_ _05749_ VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11430_ _07315_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11361_ _07277_ VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__clkbuf_1
X_10312_ _05766_ VGND VGND VPWR VPWR _06599_ sky130_fd_sc_hd__clkbuf_4
X_13100_ _06851_ _07186_ _06856_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__o21a_1
X_11292_ net1981 _05786_ _07238_ VGND VGND VPWR VPWR _07241_ sky130_fd_sc_hd__mux2_1
X_13031_ net1383 VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__clkbuf_1
X_10243_ net1695 _05786_ _06558_ VGND VGND VPWR VPWR _06561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13249__770 clknet_1_1__leaf__08343_ VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__inv_2
X_10174_ _06392_ _06493_ _06496_ _05556_ VGND VGND VPWR VPWR _06497_ sky130_fd_sc_hd__a22o_1
X_17770_ net850 _01332_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_14982_ CPU.registerFile\[27\]\[16\] CPU.registerFile\[26\]\[16\] _02768_ VGND VGND
+ VPWR VPWR _03048_ sky130_fd_sc_hd__mux2_1
X_16721_ _06172_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__buf_4
X_14111__253 clknet_1_0__leaf__08496_ VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__inv_2
X_14185__321 clknet_1_1__leaf__08502_ VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__inv_2
X_16652_ CPU.registerFile\[20\]\[15\] CPU.registerFile\[21\]\[15\] _04287_ VGND VGND
+ VPWR VPWR _04364_ sky130_fd_sc_hd__mux2_1
X_13864_ clknet_1_1__leaf__08462_ VGND VGND VPWR VPWR _08471_ sky130_fd_sc_hd__buf_1
Xclkbuf_1_0__f__08466_ clknet_0__08466_ VGND VGND VPWR VPWR clknet_1_0__leaf__08466_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12815_ _05270_ _06861_ _06869_ _08105_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__o211a_1
X_16583_ CPU.aluIn1\[13\] _04054_ _04296_ _04259_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18322_ net143 _01850_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_15534_ _03584_ _03585_ _08541_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__mux2_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ _08068_ VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ net1264 _01781_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_15465_ _08543_ _03516_ _03518_ _03307_ VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__a211o_1
XFILLER_0_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12677_ _06601_ net2502 _08029_ VGND VGND VPWR VPWR _08032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17204_ CPU.registerFile\[19\]\[29\] CPU.registerFile\[18\]\[29\] _03745_ VGND VGND
+ VPWR VPWR _04902_ sky130_fd_sc_hd__mux2_1
X_14416_ CPU.registerFile\[8\]\[2\] _08526_ _08659_ _08622_ VGND VGND VPWR VPWR _08660_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11628_ _07434_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__clkbuf_1
X_18184_ net1195 _01712_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[23\] sky130_fd_sc_hd__dfxtp_2
X_15396_ CPU.registerFile\[5\]\[26\] CPU.registerFile\[4\]\[26\] _03105_ VGND VGND
+ VPWR VPWR _03452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17135_ _08397_ _04832_ _04834_ _08400_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__a211o_1
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14347_ _08574_ _08579_ _08591_ _08592_ VGND VGND VPWR VPWR _08593_ sky130_fd_sc_hd__o211a_1
X_11559_ _07397_ VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold607 CPU.registerFile\[20\]\[15\] VGND VGND VPWR VPWR net1904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 CPU.registerFile\[5\]\[16\] VGND VGND VPWR VPWR net1915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13564__951 clknet_1_0__leaf__08441_ VGND VGND VPWR VPWR net1007 sky130_fd_sc_hd__inv_2
XFILLER_0_122_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold629 mapped_spi_flash.rcv_data\[9\] VGND VGND VPWR VPWR net1926 sky130_fd_sc_hd__dlygate4sd3_1
X_17066_ _04545_ _04750_ _04767_ _04500_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__a211o_2
X_14278_ CPU.registerFile\[22\]\[0\] CPU.registerFile\[23\]\[0\] _08523_ VGND VGND
+ VPWR VPWR _08524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16017_ _03696_ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__buf_6
X_13229_ clknet_1_0__leaf__08341_ VGND VGND VPWR VPWR _08342_ sky130_fd_sc_hd__buf_1
XFILLER_0_122_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1307 CPU.registerFile\[8\]\[19\] VGND VGND VPWR VPWR net2604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1318 CPU.registerFile\[25\]\[2\] VGND VGND VPWR VPWR net2615 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17968_ net979 _01496_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold1329 CPU.registerFile\[9\]\[8\] VGND VGND VPWR VPWR net2626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16919_ CPU.aluIn1\[21\] _04458_ _04624_ _04259_ VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__o211a_1
X_17899_ clknet_leaf_26_clk _01427_ VGND VGND VPWR VPWR CPU.instr\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_95_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09322_ _05563_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09253_ _05600_ _05601_ _05604_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__or3b_1
XFILLER_0_8_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09184_ _05535_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13718__1090 clknet_1_1__leaf__08456_ VGND VGND VPWR VPWR net1146 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__04980_ clknet_0__04980_ VGND VGND VPWR VPWR clknet_1_0__leaf__04980_
+ sky130_fd_sc_hd__clkbuf_16
X_08968_ _05319_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08899_ _05250_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__buf_2
X_10930_ mapped_spi_flash.cmd_addr\[29\] _06983_ _06985_ mapped_spi_flash.cmd_addr\[28\]
+ VGND VGND VPWR VPWR _06990_ sky130_fd_sc_hd__a22o_1
X_10861_ _06935_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12600_ _07990_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__clkbuf_1
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10792_ CPU.aluReg\[28\] _06882_ _06869_ VGND VGND VPWR VPWR _06883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12531_ _07953_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15250_ CPU.registerFile\[6\]\[22\] CPU.registerFile\[7\]\[22\] _02982_ VGND VGND
+ VPWR VPWR _03310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12462_ net2147 _07374_ _07883_ VGND VGND VPWR VPWR _07917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11413_ _07304_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15181_ _08596_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12393_ _07880_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__clkbuf_1
X_11344_ net1948 _06465_ _07260_ VGND VGND VPWR VPWR _07268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13286__789 clknet_1_0__leaf__08345_ VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__inv_2
X_18940_ net714 _02460_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_11275_ _06653_ net2376 _07223_ VGND VGND VPWR VPWR _07231_ sky130_fd_sc_hd__mux2_1
X_13014_ net2429 _07368_ _08203_ VGND VGND VPWR VPWR _08211_ sky130_fd_sc_hd__mux2_1
X_10226_ _05530_ _06544_ _06546_ _05855_ _05799_ VGND VGND VPWR VPWR _06547_ sky130_fd_sc_hd__o2111a_1
X_18871_ net645 _02391_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_17822_ net902 _01384_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10157_ _05555_ _05269_ _05526_ _05799_ _05442_ VGND VGND VPWR VPWR _06481_ sky130_fd_sc_hd__a2111oi_1
Xhold4 mapped_spi_ram.state\[0\] VGND VGND VPWR VPWR net1301 sky130_fd_sc_hd__dlygate4sd3_1
X_14965_ _02826_ _03026_ _03031_ _02746_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__o211a_1
X_17753_ net838 _01319_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_10088_ _06414_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16704_ net2645 _04054_ _04414_ _04259_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__o211a_1
X_17684_ _05213_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__clkbuf_1
X_14896_ _06012_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__buf_4
XFILLER_0_159_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16635_ _08396_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__08449_ clknet_0__08449_ VGND VGND VPWR VPWR clknet_1_0__leaf__08449_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16566_ _04277_ _04278_ _04279_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__mux2_1
X_15924__663 clknet_1_1__leaf__03688_ VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__inv_2
X_18305_ net126 _01833_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_15517_ CPU.registerFile\[16\]\[30\] _08527_ _03568_ _08530_ VGND VGND VPWR VPWR
+ _03569_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12729_ _06653_ net2514 _08051_ VGND VGND VPWR VPWR _08059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16497_ _04211_ _04212_ _03961_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18236_ net1247 net20 VGND VGND VPWR VPWR mapped_spi_flash.div_counter\[5\] sky130_fd_sc_hd__dfxtp_1
X_15448_ CPU.registerFile\[20\]\[28\] _08523_ _03501_ _08578_ VGND VGND VPWR VPWR
+ _03502_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18167_ net1178 _01695_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[6\] sky130_fd_sc_hd__dfxtp_1
X_13488__882 clknet_1_1__leaf__08434_ VGND VGND VPWR VPWR net938 sky130_fd_sc_hd__inv_2
X_15379_ CPU.registerFile\[28\]\[26\] CPU.registerFile\[29\]\[26\] _03212_ VGND VGND
+ VPWR VPWR _03435_ sky130_fd_sc_hd__mux2_1
X_17118_ _03765_ _04815_ _04817_ _04521_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__a211o_1
Xhold404 CPU.registerFile\[19\]\[18\] VGND VGND VPWR VPWR net1701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold415 CPU.registerFile\[6\]\[16\] VGND VGND VPWR VPWR net1712 sky130_fd_sc_hd__dlygate4sd3_1
X_18098_ net1109 _01626_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xhold426 CPU.registerFile\[6\]\[18\] VGND VGND VPWR VPWR net1723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13878__1234 clknet_1_0__leaf__08472_ VGND VGND VPWR VPWR net1290 sky130_fd_sc_hd__inv_2
Xhold437 CPU.registerFile\[3\]\[9\] VGND VGND VPWR VPWR net1734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 CPU.registerFile\[5\]\[1\] VGND VGND VPWR VPWR net1745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 CPU.registerFile\[10\]\[5\] VGND VGND VPWR VPWR net1756 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17049_ CPU.registerFile\[30\]\[25\] CPU.registerFile\[31\]\[25\] _04605_ VGND VGND
+ VPWR VPWR _04751_ sky130_fd_sc_hd__mux2_1
X_09940_ _05460_ _06271_ _05451_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__a21o_1
Xclkbuf_1_1__f__03687_ clknet_0__03687_ VGND VGND VPWR VPWR clknet_1_1__leaf__03687_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _06203_ _05763_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__or2_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 CPU.registerFile\[20\]\[20\] VGND VGND VPWR VPWR net2401 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1115 CPU.registerFile\[2\]\[16\] VGND VGND VPWR VPWR net2412 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1126 CPU.registerFile\[24\]\[29\] VGND VGND VPWR VPWR net2423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 CPU.registerFile\[30\]\[1\] VGND VGND VPWR VPWR net2434 sky130_fd_sc_hd__dlygate4sd3_1
X_17311__725 clknet_1_0__leaf__04981_ VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__inv_2
Xhold1148 CPU.registerFile\[22\]\[11\] VGND VGND VPWR VPWR net2445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 CPU.registerFile\[30\]\[10\] VGND VGND VPWR VPWR net2456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09305_ _05652_ _05558_ _05655_ _05656_ _05236_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09236_ CPU.aluIn1\[4\] _05586_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09167_ _05421_ _05426_ _05518_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09098_ _05308_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold960 CPU.registerFile\[2\]\[21\] VGND VGND VPWR VPWR net2257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 CPU.registerFile\[22\]\[20\] VGND VGND VPWR VPWR net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold982 CPU.registerFile\[29\]\[27\] VGND VGND VPWR VPWR net2279 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ _05591_ _07094_ _05590_ _07023_ VGND VGND VPWR VPWR _07096_ sky130_fd_sc_hd__a31o_1
Xhold993 CPU.registerFile\[16\]\[12\] VGND VGND VPWR VPWR net2290 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10011_ mapped_spi_ram.rcv_data\[16\] _05685_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__and2_1
X_17286__702 clknet_1_1__leaf__04979_ VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__inv_2
X_14750_ _02733_ _02734_ CPU.registerFile\[9\]\[10\] VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__a21o_1
X_11962_ _07612_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__clkbuf_1
X_10913_ CPU.mem_rstrb _05859_ mapped_spi_flash.state\[2\] VGND VGND VPWR VPWR _06975_
+ sky130_fd_sc_hd__a21boi_2
XFILLER_0_98_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14681_ CPU.registerFile\[19\]\[9\] CPU.registerFile\[18\]\[9\] _02753_ VGND VGND
+ VPWR VPWR _02754_ sky130_fd_sc_hd__mux2_1
X_11893_ _06622_ net1841 _07573_ VGND VGND VPWR VPWR _07576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16420_ _06474_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__clkbuf_4
X_10844_ net2653 _06921_ _06922_ VGND VGND VPWR VPWR _06923_ sky130_fd_sc_hd__mux2_1
X_15646__446 clknet_1_0__leaf__03642_ VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__inv_2
XFILLER_0_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16351_ CPU.registerFile\[0\]\[8\] _03828_ _04068_ _04069_ VGND VGND VPWR VPWR _04070_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10775_ _06868_ VGND VGND VPWR VPWR _06869_ sky130_fd_sc_hd__buf_4
XFILLER_0_94_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14223__354 clknet_1_1__leaf__08507_ VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__inv_2
XFILLER_0_55_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15302_ CPU.registerFile\[21\]\[24\] _02752_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__or2_1
X_12514_ net1947 _07358_ _07942_ VGND VGND VPWR VPWR _07945_ sky130_fd_sc_hd__mux2_1
X_19070_ net62 _02590_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_16282_ CPU.registerFile\[19\]\[6\] CPU.registerFile\[18\]\[6\] _03923_ VGND VGND
+ VPWR VPWR _04003_ sky130_fd_sc_hd__mux2_1
X_18021_ net1032 _01549_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15233_ CPU.registerFile\[28\]\[22\] CPU.registerFile\[29\]\[22\] _03212_ VGND VGND
+ VPWR VPWR _03293_ sky130_fd_sc_hd__mux2_1
X_12445_ _07908_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15164_ _03138_ _03139_ CPU.registerFile\[9\]\[20\] VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__a21o_1
X_12376_ _06641_ net1839 _07870_ VGND VGND VPWR VPWR _07872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__03641_ _03641_ VGND VGND VPWR VPWR clknet_0__03641_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11327_ net2480 _06267_ _07249_ VGND VGND VPWR VPWR _07259_ sky130_fd_sc_hd__mux2_1
X_15095_ CPU.registerFile\[19\]\[19\] CPU.registerFile\[18\]\[19\] _03157_ VGND VGND
+ VPWR VPWR _03158_ sky130_fd_sc_hd__mux2_1
X_18923_ net697 _02443_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11258_ _06636_ net1899 _07212_ VGND VGND VPWR VPWR _07222_ sky130_fd_sc_hd__mux2_1
X_10209_ net2263 _06530_ net15 VGND VGND VPWR VPWR _06531_ sky130_fd_sc_hd__mux2_1
X_18854_ net628 _00007_ VGND VGND VPWR VPWR mapped_spi_flash.state\[3\] sky130_fd_sc_hd__dfxtp_2
X_11189_ mapped_spi_flash.rcv_bitcount\[5\] _07128_ VGND VGND VPWR VPWR _07180_ sky130_fd_sc_hd__nand2_1
X_13910__72 clknet_1_0__leaf__08476_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__inv_2
X_17805_ net885 _01367_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_18785_ net574 _02309_ VGND VGND VPWR VPWR CPU.aluReg\[15\] sky130_fd_sc_hd__dfxtp_1
X_15997_ _06172_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__buf_4
X_13684__1059 clknet_1_1__leaf__08453_ VGND VGND VPWR VPWR net1115 sky130_fd_sc_hd__inv_2
X_14948_ CPU.registerFile\[13\]\[15\] CPU.registerFile\[12\]\[15\] _02935_ VGND VGND
+ VPWR VPWR _03015_ sky130_fd_sc_hd__mux2_1
X_17736_ net821 _01302_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17667_ _05200_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__clkbuf_1
X_14879_ _08410_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16618_ _03963_ _04328_ _04330_ _04006_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__a211o_1
X_17598_ _05125_ _05153_ _05154_ _05155_ net1585 VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__a32o_1
XFILLER_0_147_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16549_ _04099_ _04260_ _04262_ _04105_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09021_ CPU.aluIn1\[23\] _05371_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18219_ net1230 _01747_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold201 _02273_ VGND VGND VPWR VPWR net1498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 _02365_ VGND VGND VPWR VPWR net1509 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold223 mapped_spi_flash.cmd_addr\[20\] VGND VGND VPWR VPWR net1520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _02287_ VGND VGND VPWR VPWR net1531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _02371_ VGND VGND VPWR VPWR net1542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 CPU.cycles\[14\] VGND VGND VPWR VPWR net1553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold267 CPU.registerFile\[31\]\[19\] VGND VGND VPWR VPWR net1564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 CPU.cycles\[5\] VGND VGND VPWR VPWR net1575 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _05427_ _06255_ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__nand2_1
Xhold289 CPU.cycles\[21\] VGND VGND VPWR VPWR net1586 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751__541 clknet_1_1__leaf__03652_ VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__inv_2
X_09854_ _05427_ _06189_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__nand2_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _06123_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__buf_4
XFILLER_0_147_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17347__8 clknet_1_0__leaf__04984_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__inv_2
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410__32 clknet_1_1__leaf__05014_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__inv_2
XFILLER_0_48_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10560_ net1729 _05853_ _06739_ VGND VGND VPWR VPWR _06746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09219_ CPU.aluIn1\[5\] CPU.Bimm\[5\] VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__nor2_1
XFILLER_0_161_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10491_ net2075 _05853_ _06702_ VGND VGND VPWR VPWR _06709_ sky130_fd_sc_hd__mux2_1
X_12230_ net8 net1298 _07782_ VGND VGND VPWR VPWR _07786_ sky130_fd_sc_hd__and3_1
XFILLER_0_161_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12161_ _07715_ _07735_ VGND VGND VPWR VPWR _07736_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11112_ net1398 _07135_ VGND VGND VPWR VPWR _07136_ sky130_fd_sc_hd__or2_1
X_12092_ _07686_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__clkbuf_1
Xhold790 CPU.registerFile\[11\]\[23\] VGND VGND VPWR VPWR net2087 sky130_fd_sc_hd__dlygate4sd3_1
X_11043_ net1491 _07054_ _07081_ _07069_ VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__o211a_1
X_14802_ _02831_ _02832_ CPU.registerFile\[1\]\[11\] VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18570_ net391 net27 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_12994_ _08200_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14733_ CPU.registerFile\[20\]\[10\] _08839_ _02804_ _08841_ VGND VGND VPWR VPWR
+ _02805_ sky130_fd_sc_hd__o211a_1
X_17521_ _08335_ _06113_ _05073_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__o21ai_1
X_11945_ _07603_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__clkbuf_1
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13877__1233 clknet_1_0__leaf__08472_ VGND VGND VPWR VPWR net1289 sky130_fd_sc_hd__inv_2
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _08379_ _05017_ _06400_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_129_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _02728_ _02731_ _02737_ _08423_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__o211a_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ _06605_ net2311 _07562_ VGND VGND VPWR VPWR _07567_ sky130_fd_sc_hd__mux2_1
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16403_ CPU.registerFile\[30\]\[9\] CPU.registerFile\[31\]\[9\] _03796_ VGND VGND
+ VPWR VPWR _04121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10827_ _06909_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17383_ _04996_ _05007_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14595_ CPU.registerFile\[17\]\[7\] _08795_ VGND VGND VPWR VPWR _08834_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16334_ CPU.aluIn1\[7\] _03566_ _04053_ _03855_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__o211a_1
X_19122_ clknet_leaf_9_clk _02642_ VGND VGND VPWR VPWR CPU.PC\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10758_ _06853_ VGND VGND VPWR VPWR _06854_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_918 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19053_ net795 _02573_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_16265_ _05690_ VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__buf_2
XFILLER_0_82_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13477_ CPU.Bimm\[8\] _05788_ _08416_ VGND VGND VPWR VPWR _08430_ sky130_fd_sc_hd__mux2_1
X_10689_ net2018 _05734_ _06816_ VGND VGND VPWR VPWR _06817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15216_ _03235_ _03236_ CPU.registerFile\[1\]\[21\] VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__a21o_1
X_18004_ net1015 _01532_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_12428_ _07899_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16196_ _03735_ _03913_ _03918_ _03755_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15147_ CPU.registerFile\[20\]\[20\] _03080_ _03208_ _03082_ VGND VGND VPWR VPWR
+ _03209_ sky130_fd_sc_hd__o211a_1
X_12359_ _06624_ net1921 _07859_ VGND VGND VPWR VPWR _07863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15078_ _03098_ _03137_ _03141_ _02903_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__a211o_1
XFILLER_0_121_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18906_ net680 _02426_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_18837_ clknet_leaf_6_clk _02361_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_09570_ _05913_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__clkbuf_4
X_18768_ net557 _02292_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18699_ net488 _02223_ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15781__567 clknet_1_0__leaf__03656_ VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__inv_2
XFILLER_0_46_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_842 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09004_ _05354_ _05355_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17317__731 clknet_1_1__leaf__04981_ VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__inv_2
XFILLER_0_111_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09906_ mapped_spi_ram.rcv_data\[21\] _05761_ _05762_ mapped_spi_flash.rcv_data\[21\]
+ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ _06172_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__clkbuf_8
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09768_ _06107_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__clkbuf_1
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _05363_ _05367_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__and2b_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _07488_ _06814_ VGND VGND VPWR VPWR _07489_ sky130_fd_sc_hd__nand2_4
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512__904 clknet_1_0__leaf__08436_ VGND VGND VPWR VPWR net960 sky130_fd_sc_hd__inv_2
XFILLER_0_83_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11661_ _06813_ _07451_ VGND VGND VPWR VPWR _07452_ sky130_fd_sc_hd__nor2_4
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13400_ _08378_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10612_ net2227 _06555_ _06738_ VGND VGND VPWR VPWR _06773_ sky130_fd_sc_hd__mux2_1
X_14380_ _08557_ _08619_ _08624_ _08423_ VGND VGND VPWR VPWR _08625_ sky130_fd_sc_hd__o211a_1
X_11592_ _07414_ _07310_ VGND VGND VPWR VPWR _07415_ sky130_fd_sc_hd__nor2_2
XFILLER_0_52_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10543_ net1972 _06555_ _06701_ VGND VGND VPWR VPWR _06736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13683__1058 clknet_1_1__leaf__08453_ VGND VGND VPWR VPWR net1114 sky130_fd_sc_hd__inv_2
X_16050_ _03756_ _03776_ _08406_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__o21a_1
XFILLER_0_106_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13262_ clknet_1_1__leaf__08341_ VGND VGND VPWR VPWR _08345_ sky130_fd_sc_hd__buf_1
XFILLER_0_107_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10474_ _06661_ net2441 _06664_ VGND VGND VPWR VPWR _06699_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15758__547 clknet_1_1__leaf__03653_ VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__inv_2
XFILLER_0_161_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15001_ CPU.registerFile\[2\]\[16\] CPU.registerFile\[3\]\[16\] _02871_ VGND VGND
+ VPWR VPWR _03067_ sky130_fd_sc_hd__mux2_1
X_12213_ _07772_ net1337 _07764_ VGND VGND VPWR VPWR _07773_ sky130_fd_sc_hd__mux2_1
X_13193_ _08307_ _08308_ VGND VGND VPWR VPWR _08309_ sky130_fd_sc_hd__and2_1
X_12144_ _07703_ VGND VGND VPWR VPWR _07724_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_130_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12075_ CPU.mem_rstrb _07673_ _05858_ VGND VGND VPWR VPWR _07674_ sky130_fd_sc_hd__o21a_1
X_16952_ _04579_ _04580_ CPU.registerFile\[17\]\[22\] VGND VGND VPWR VPWR _04657_
+ sky130_fd_sc_hd__a21o_1
X_11026_ mapped_spi_flash.cmd_addr\[9\] _07066_ _07039_ VGND VGND VPWR VPWR _07067_
+ sky130_fd_sc_hd__mux2_1
X_16883_ CPU.registerFile\[9\]\[21\] _04460_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__or2_1
X_18622_ net443 _02146_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18553_ net374 _02077_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12977_ _08191_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14229__360 clknet_1_0__leaf__08507_ VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__inv_2
X_17504_ _05055_ _06196_ _05061_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__or3_1
X_14716_ CPU.registerFile\[2\]\[9\] CPU.registerFile\[3\]\[9\] _08629_ VGND VGND VPWR
+ VPWR _02789_ sky130_fd_sc_hd__mux2_1
X_11928_ _06657_ net2032 _07584_ VGND VGND VPWR VPWR _07594_ sky130_fd_sc_hd__mux2_1
X_18484_ net305 _02008_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17435_ _08310_ _08330_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__or2_1
X_14647_ _02719_ _02720_ _08609_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__mux2_1
X_11859_ _07557_ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_18 _04642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14578_ CPU.registerFile\[10\]\[6\] CPU.registerFile\[11\]\[6\] _08564_ VGND VGND
+ VPWR VPWR _08818_ sky130_fd_sc_hd__mux2_1
XANTENNA_29 _06031_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17366_ _06854_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19105_ net88 _02625_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_16317_ _08396_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19036_ net778 _02556_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_16248_ _03692_ _03949_ _03969_ _03601_ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_1__f__08462_ clknet_0__08462_ VGND VGND VPWR VPWR clknet_1_1__leaf__08462_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__08493_ _08493_ VGND VGND VPWR VPWR clknet_0__08493_ sky130_fd_sc_hd__clkbuf_16
X_16179_ CPU.registerFile\[6\]\[4\] CPU.registerFile\[7\]\[4\] _03717_ VGND VGND VPWR
+ VPWR _03902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09622_ CPU.PC\[6\] CPU.Bimm\[6\] _05913_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__and3_1
X_09553_ _05372_ _05532_ _05534_ CPU.aluReg\[23\] VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09484_ _05384_ _05385_ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14057__205 clknet_1_0__leaf__08490_ VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__inv_2
X_13876__1232 clknet_1_0__leaf__08472_ VGND VGND VPWR VPWR net1288 sky130_fd_sc_hd__inv_2
X_10190_ mapped_spi_ram.rcv_data\[25\] _05857_ _06462_ VGND VGND VPWR VPWR _06512_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12900_ _05839_ net2136 _08145_ VGND VGND VPWR VPWR _08151_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__08482_ clknet_0__08482_ VGND VGND VPWR VPWR clknet_1_0__leaf__08482_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12831_ net2280 VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__clkbuf_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ _06339_ _03583_ _03600_ _03601_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__a211o_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12762_ _06617_ net2112 _08076_ VGND VGND VPWR VPWR _08077_ sky130_fd_sc_hd__mux2_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _08741_ _08742_ _08578_ VGND VGND VPWR VPWR _08743_ sky130_fd_sc_hd__mux2_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ net2389 _07362_ _07475_ VGND VGND VPWR VPWR _07480_ sky130_fd_sc_hd__mux2_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15481_ _08521_ _03531_ _03533_ _08590_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__a211o_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _08028_ VGND VGND VPWR VPWR _08040_ sky130_fd_sc_hd__buf_4
XFILLER_0_49_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ CPU.registerFile\[6\]\[30\] CPU.registerFile\[7\]\[30\] _03847_ VGND VGND
+ VPWR VPWR _04917_ sky130_fd_sc_hd__mux2_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14432_ CPU.registerFile\[17\]\[3\] _06456_ VGND VGND VPWR VPWR _08675_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11644_ net2248 _07362_ _07438_ VGND VGND VPWR VPWR _07443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17151_ CPU.registerFile\[2\]\[28\] CPU.registerFile\[3\]\[28\] _03759_ VGND VGND
+ VPWR VPWR _04850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14363_ CPU.registerFile\[28\]\[1\] CPU.registerFile\[29\]\[1\] _08538_ VGND VGND
+ VPWR VPWR _08608_ sky130_fd_sc_hd__mux2_1
X_11575_ net1674 _07362_ _07401_ VGND VGND VPWR VPWR _07406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16102_ CPU.registerFile\[2\]\[2\] CPU.registerFile\[3\]\[2\] _03693_ VGND VGND VPWR
+ VPWR _03827_ sky130_fd_sc_hd__mux2_1
X_17082_ _03765_ _04780_ _04782_ _04521_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__a211o_1
XFILLER_0_123_934 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10526_ _06727_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__clkbuf_1
X_14294_ _06035_ VGND VGND VPWR VPWR _08540_ sky130_fd_sc_hd__buf_4
XFILLER_0_40_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16033_ CPU.registerFile\[22\]\[0\] CPU.registerFile\[23\]\[0\] _03759_ VGND VGND
+ VPWR VPWR _03760_ sky130_fd_sc_hd__mux2_1
X_10457_ _06690_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13176_ _08297_ net1548 VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__nor2_1
X_10388_ _06650_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__clkbuf_1
X_12127_ _07696_ _07711_ VGND VGND VPWR VPWR _07712_ sky130_fd_sc_hd__or2_1
X_17984_ net995 _01512_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_16935_ _04347_ _04636_ _04639_ _04521_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__a211o_1
X_12058_ _07663_ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__clkbuf_1
X_11009_ mapped_spi_flash.cmd_addr\[11\] _07051_ _07039_ VGND VGND VPWR VPWR _07052_
+ sky130_fd_sc_hd__mux2_1
X_16866_ _04479_ _04567_ _04572_ _04446_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__o211a_1
X_18605_ net426 _02129_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_15817_ _07001_ per_uart.uart0.enable16_counter\[15\] _08359_ VGND VGND VPWR VPWR
+ _03677_ sky130_fd_sc_hd__and3_1
X_16797_ _08393_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18536_ net357 _02060_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_14162__300 clknet_1_1__leaf__08500_ VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__inv_2
X_18467_ net288 _00011_ VGND VGND VPWR VPWR mapped_spi_ram.state\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18398_ net219 _01926_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14006__159 clknet_1_0__leaf__08485_ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__inv_2
XFILLER_0_70_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19019_ net761 _02539_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[4\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__08445_ clknet_0__08445_ VGND VGND VPWR VPWR clknet_1_1__leaf__08445_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__08476_ _08476_ VGND VGND VPWR VPWR clknet_0__08476_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08984_ _05321_ _05324_ _05329_ _05334_ _05335_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_139_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09605_ CPU.Bimm\[5\] _05913_ CPU.PC\[5\] VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__a21o_1
X_13682__1057 clknet_1_1__leaf__08453_ VGND VGND VPWR VPWR net1113 sky130_fd_sc_hd__inv_2
X_09536_ _05879_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__buf_2
XFILLER_0_78_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09467_ _05400_ _05814_ _05502_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09398_ _05748_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11360_ net1759 _05786_ _07274_ VGND VGND VPWR VPWR _07277_ sky130_fd_sc_hd__mux2_1
X_10311_ _06598_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11291_ _07240_ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13030_ CPU.registerFile\[4\]\[29\] net1382 _08217_ VGND VGND VPWR VPWR _08220_ sky130_fd_sc_hd__mux2_1
X_10242_ _06560_ VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10173_ _06312_ _06393_ _06494_ _06395_ _06495_ VGND VGND VPWR VPWR _06496_ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14981_ _03045_ _03046_ _02851_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__mux2_1
X_16720_ _04427_ _04429_ _04153_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13518__910 clknet_1_1__leaf__08436_ VGND VGND VPWR VPWR net966 sky130_fd_sc_hd__inv_2
X_16651_ CPU.registerFile\[22\]\[15\] CPU.registerFile\[23\]\[15\] _04362_ VGND VGND
+ VPWR VPWR _04363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__08465_ clknet_0__08465_ VGND VGND VPWR VPWR clknet_1_0__leaf__08465_
+ sky130_fd_sc_hd__clkbuf_16
X_13968__125 clknet_1_1__leaf__08481_ VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__inv_2
X_12814_ net2599 _08104_ VGND VGND VPWR VPWR _08105_ sky130_fd_sc_hd__xor2_1
X_16582_ _04141_ _04276_ _04295_ _04096_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__a211o_1
X_18321_ net142 _01849_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_15533_ CPU.registerFile\[13\]\[30\] CPU.registerFile\[12\]\[30\] _08794_ VGND VGND
+ VPWR VPWR _03585_ sky130_fd_sc_hd__mux2_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _06601_ net2139 _08065_ VGND VGND VPWR VPWR _08068_ sky130_fd_sc_hd__mux2_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15464_ CPU.registerFile\[8\]\[28\] _08545_ _03517_ _03268_ VGND VGND VPWR VPWR _03518_
+ sky130_fd_sc_hd__o211a_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18252_ net1263 _01780_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _08031_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14415_ _08567_ _08569_ CPU.registerFile\[9\]\[2\] VGND VGND VPWR VPWR _08659_ sky130_fd_sc_hd__a21o_1
X_17203_ _04899_ _04900_ _03742_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__mux2_1
X_11627_ net2531 _07345_ _07427_ VGND VGND VPWR VPWR _07434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15395_ CPU.registerFile\[6\]\[26\] CPU.registerFile\[7\]\[26\] _08536_ VGND VGND
+ VPWR VPWR _03451_ sky130_fd_sc_hd__mux2_1
X_18183_ net1194 net1517 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14346_ _05876_ VGND VGND VPWR VPWR _08592_ sky130_fd_sc_hd__buf_4
X_17134_ CPU.registerFile\[16\]\[27\] _04656_ _04494_ _04833_ VGND VGND VPWR VPWR
+ _04834_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11558_ net1817 _07345_ _07390_ VGND VGND VPWR VPWR _07397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold608 CPU.registerFile\[17\]\[15\] VGND VGND VPWR VPWR net1905 sky130_fd_sc_hd__dlygate4sd3_1
X_17065_ _04758_ _04766_ _04542_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__o21a_1
X_10509_ _06718_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__clkbuf_1
X_14277_ _08522_ VGND VGND VPWR VPWR _08523_ sky130_fd_sc_hd__buf_4
Xhold619 CPU.registerFile\[21\]\[10\] VGND VGND VPWR VPWR net1916 sky130_fd_sc_hd__dlygate4sd3_1
X_11489_ _07355_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16016_ _03738_ _03740_ _03742_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__mux2_1
X_13228_ clknet_1_0__leaf__08340_ VGND VGND VPWR VPWR _08341_ sky130_fd_sc_hd__buf_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ net1620 _08287_ VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__xor2_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ net978 _01495_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[5\] sky130_fd_sc_hd__dfxtp_1
Xhold1308 CPU.PC\[16\] VGND VGND VPWR VPWR net2605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1319 CPU.registerFile\[25\]\[25\] VGND VGND VPWR VPWR net2616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16918_ _04545_ _04604_ _04623_ _04500_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__a211o_1
X_17898_ clknet_leaf_26_clk _01426_ VGND VGND VPWR VPWR CPU.instr\[5\] sky130_fd_sc_hd__dfxtp_4
X_16849_ CPU.registerFile\[5\]\[20\] CPU.registerFile\[4\]\[20\] _04428_ VGND VGND
+ VPWR VPWR _04556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09321_ _05626_ _05627_ _05566_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__a21o_1
X_18519_ net340 _02043_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09252_ _05602_ _05603_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09183_ _05534_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15819__569 clknet_1_0__leaf__03656_ VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__inv_2
XFILLER_0_141_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0__08459_ _08459_ VGND VGND VPWR VPWR clknet_0__08459_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08967_ _05316_ _05318_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__or2_2
X_14169__306 clknet_1_1__leaf__08501_ VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__inv_2
X_08898_ _05249_ VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10860_ net2669 _06934_ _06922_ VGND VGND VPWR VPWR _06935_ sky130_fd_sc_hd__mux2_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09519_ _05381_ _05382_ _05391_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__and3_1
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10791_ CPU.aluIn1\[28\] _06879_ _06881_ VGND VGND VPWR VPWR _06882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ net2040 _07374_ _07919_ VGND VGND VPWR VPWR _07953_ sky130_fd_sc_hd__mux2_1
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_776 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12461_ _07916_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11412_ net1778 _06465_ _07296_ VGND VGND VPWR VPWR _07304_ sky130_fd_sc_hd__mux2_1
X_15180_ _03229_ _03240_ _03241_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__o21a_2
XFILLER_0_62_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12392_ _06657_ net2490 _07870_ VGND VGND VPWR VPWR _07880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14131_ clknet_1_0__leaf__08495_ VGND VGND VPWR VPWR _08498_ sky130_fd_sc_hd__buf_1
X_11343_ _07267_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11274_ _07230_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13797__1161 clknet_1_1__leaf__08464_ VGND VGND VPWR VPWR net1217 sky130_fd_sc_hd__inv_2
XFILLER_0_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13013_ _08210_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__clkbuf_1
X_10225_ _05530_ _06545_ VGND VGND VPWR VPWR _06546_ sky130_fd_sc_hd__nand2_1
X_18870_ net644 _02390_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_17821_ net901 _01383_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_10156_ _05794_ _06477_ _06479_ VGND VGND VPWR VPWR _06480_ sky130_fd_sc_hd__o21ai_1
X_14035__185 clknet_1_0__leaf__08488_ VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__inv_2
Xhold5 _07676_ VGND VGND VPWR VPWR net1302 sky130_fd_sc_hd__dlygate4sd3_1
X_17752_ net837 _01318_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_14964_ _03027_ _03028_ _03030_ _08870_ VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__a211o_1
X_10087_ net2298 _06413_ _06293_ VGND VGND VPWR VPWR _06414_ sky130_fd_sc_hd__mux2_1
X_13594__978 clknet_1_1__leaf__08444_ VGND VGND VPWR VPWR net1034 sky130_fd_sc_hd__inv_2
X_16703_ _04141_ _04395_ _04413_ _04096_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__a211o_1
X_17683_ _05207_ _05212_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__and2_1
X_14895_ _08837_ _02959_ _02962_ _08802_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__a211o_1
X_16634_ _04344_ _04345_ _04153_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__08448_ clknet_0__08448_ VGND VGND VPWR VPWR clknet_1_0__leaf__08448_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16565_ _03741_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__buf_4
X_10989_ _07008_ _07034_ VGND VGND VPWR VPWR _07035_ sky130_fd_sc_hd__or2_1
X_17719__50 clknet_1_0__leaf__05015_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__inv_2
X_18304_ net125 _01832_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15516_ CPU.registerFile\[17\]\[30\] _08528_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12728_ _08058_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__clkbuf_1
X_16496_ CPU.registerFile\[20\]\[11\] CPU.registerFile\[21\]\[11\] _03883_ VGND VGND
+ VPWR VPWR _04212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18235_ net1246 net19 VGND VGND VPWR VPWR mapped_spi_flash.div_counter\[4\] sky130_fd_sc_hd__dfxtp_1
X_15623__425 clknet_1_1__leaf__03640_ VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__inv_2
X_12659_ _06651_ net2038 _08015_ VGND VGND VPWR VPWR _08022_ sky130_fd_sc_hd__mux2_1
X_15447_ CPU.registerFile\[21\]\[28\] _02752_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18166_ net1177 _01694_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15378_ CPU.registerFile\[30\]\[26\] CPU.registerFile\[31\]\[26\] _03291_ VGND VGND
+ VPWR VPWR _03434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17117_ CPU.registerFile\[0\]\[27\] _04637_ _04472_ _04816_ VGND VGND VPWR VPWR _04817_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14329_ CPU.registerFile\[6\]\[0\] CPU.registerFile\[7\]\[0\] _08522_ VGND VGND VPWR
+ VPWR _08575_ sky130_fd_sc_hd__mux2_1
Xhold405 CPU.registerFile\[6\]\[0\] VGND VGND VPWR VPWR net1702 sky130_fd_sc_hd__dlygate4sd3_1
X_18097_ net1108 _01625_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13681__1056 clknet_1_0__leaf__08453_ VGND VGND VPWR VPWR net1112 sky130_fd_sc_hd__inv_2
Xhold416 CPU.registerFile\[28\]\[12\] VGND VGND VPWR VPWR net1713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 CPU.registerFile\[10\]\[3\] VGND VGND VPWR VPWR net1724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold438 CPU.registerFile\[28\]\[8\] VGND VGND VPWR VPWR net1735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 CPU.registerFile\[5\]\[11\] VGND VGND VPWR VPWR net1746 sky130_fd_sc_hd__dlygate4sd3_1
X_17048_ _04502_ _04737_ _04741_ _04749_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__a31o_1
Xclkbuf_1_1__f__03686_ clknet_0__03686_ VGND VGND VPWR VPWR clknet_1_1__leaf__03686_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ mapped_spi_ram.rcv_data\[22\] _05857_ _05762_ net1416 VGND VGND VPWR VPWR
+ _06205_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1105 CPU.registerFile\[8\]\[22\] VGND VGND VPWR VPWR net2402 sky130_fd_sc_hd__dlygate4sd3_1
X_18999_ clknet_leaf_13_clk _02519_ VGND VGND VPWR VPWR CPU.aluIn1\[16\] sky130_fd_sc_hd__dfxtp_4
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 CPU.registerFile\[14\]\[25\] VGND VGND VPWR VPWR net2413 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1127 CPU.registerFile\[14\]\[9\] VGND VGND VPWR VPWR net2424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 CPU.registerFile\[11\]\[7\] VGND VGND VPWR VPWR net2435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 CPU.registerFile\[13\]\[19\] VGND VGND VPWR VPWR net2446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09304_ _05653_ _05654_ _05558_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09235_ CPU.aluIn1\[4\] _05586_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15598__402 clknet_1_0__leaf__03638_ VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__inv_2
X_09166_ _05427_ _05513_ _05517_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14140__280 clknet_1_1__leaf__08498_ VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__inv_2
XFILLER_0_90_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09097_ _05263_ _05266_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold950 CPU.registerFile\[11\]\[14\] VGND VGND VPWR VPWR net2247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 CPU.registerFile\[16\]\[0\] VGND VGND VPWR VPWR net2258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold972 CPU.registerFile\[20\]\[11\] VGND VGND VPWR VPWR net2269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 _08114_ VGND VGND VPWR VPWR net2280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 CPU.registerFile\[11\]\[26\] VGND VGND VPWR VPWR net2291 sky130_fd_sc_hd__dlygate4sd3_1
X_10010_ mapped_spi_ram.rcv_data\[0\] _05761_ _05762_ net1379 VGND VGND VPWR VPWR
+ _06339_ sky130_fd_sc_hd__a22o_4
XFILLER_0_101_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09999_ CPU.PC\[9\] _05885_ VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__xnor2_1
X_11961_ _06622_ net2141 _07609_ VGND VGND VPWR VPWR _07612_ sky130_fd_sc_hd__mux2_1
X_10912_ net1393 VGND VGND VPWR VPWR _06974_ sky130_fd_sc_hd__inv_2
X_14680_ _02752_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__buf_4
X_11892_ _07575_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13631_ clknet_1_0__leaf__08440_ VGND VGND VPWR VPWR _08448_ sky130_fd_sc_hd__buf_1
XFILLER_0_79_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10843_ _06868_ VGND VGND VPWR VPWR _06922_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16350_ _03985_ _03986_ CPU.registerFile\[1\]\[8\] VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10774_ _06864_ _06867_ _05236_ VGND VGND VPWR VPWR _06868_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_109_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13292__794 clknet_1_0__leaf__08361_ VGND VGND VPWR VPWR net850 sky130_fd_sc_hd__inv_2
X_12513_ _07944_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__clkbuf_1
X_15301_ CPU.registerFile\[22\]\[24\] CPU.registerFile\[23\]\[24\] _02998_ VGND VGND
+ VPWR VPWR _03359_ sky130_fd_sc_hd__mux2_1
X_16281_ _04000_ _04001_ _03961_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18020_ net1031 _01548_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12444_ net1764 _07356_ _07906_ VGND VGND VPWR VPWR _07908_ sky130_fd_sc_hd__mux2_1
X_15232_ CPU.registerFile\[30\]\[22\] CPU.registerFile\[31\]\[22\] _03291_ VGND VGND
+ VPWR VPWR _03292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15163_ CPU.registerFile\[10\]\[20\] CPU.registerFile\[11\]\[20\] _03183_ VGND VGND
+ VPWR VPWR _03225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12375_ _07871_ VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__03640_ _03640_ VGND VGND VPWR VPWR clknet_0__03640_ sky130_fd_sc_hd__clkbuf_16
X_11326_ _07258_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15094_ _02752_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__buf_4
X_18922_ net696 _02442_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_11257_ _07221_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10208_ net1362 VGND VGND VPWR VPWR _06530_ sky130_fd_sc_hd__clkbuf_4
X_18853_ net627 _00006_ VGND VGND VPWR VPWR mapped_spi_flash.state\[2\] sky130_fd_sc_hd__dfxtp_2
X_11188_ net1649 _07178_ _07179_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__a21boi_1
X_13602__985 clknet_1_0__leaf__08445_ VGND VGND VPWR VPWR net1041 sky130_fd_sc_hd__inv_2
X_17804_ net884 _01366_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_10139_ _05745_ _06449_ _06455_ _06463_ VGND VGND VPWR VPWR _06464_ sky130_fd_sc_hd__a211o_2
X_18784_ net573 _02308_ VGND VGND VPWR VPWR CPU.aluReg\[14\] sky130_fd_sc_hd__dfxtp_1
X_15996_ CPU.registerFile\[2\]\[0\] CPU.registerFile\[3\]\[0\] _03693_ VGND VGND VPWR
+ VPWR _03723_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17735_ net820 _01301_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_14947_ CPU.registerFile\[15\]\[15\] CPU.registerFile\[14\]\[15\] _03013_ VGND VGND
+ VPWR VPWR _03014_ sky130_fd_sc_hd__mux2_1
X_17666_ _05192_ _05198_ _05199_ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__and3_1
X_14878_ CPU.registerFile\[2\]\[13\] CPU.registerFile\[3\]\[13\] _02871_ VGND VGND
+ VPWR VPWR _02947_ sky130_fd_sc_hd__mux2_1
X_15848__595 clknet_1_1__leaf__03680_ VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__inv_2
XFILLER_0_58_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13375__869 clknet_1_1__leaf__08369_ VGND VGND VPWR VPWR net925 sky130_fd_sc_hd__inv_2
X_16617_ CPU.registerFile\[16\]\[14\] _04252_ _04090_ _04329_ VGND VGND VPWR VPWR
+ _04330_ sky130_fd_sc_hd__o211a_1
X_17597_ _05121_ _05153_ _05148_ _06973_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__o211ai_1
X_16548_ CPU.registerFile\[8\]\[13\] _04101_ _04102_ _04261_ VGND VGND VPWR VPWR _04262_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16479_ CPU.registerFile\[2\]\[11\] CPU.registerFile\[3\]\[11\] _04027_ VGND VGND
+ VPWR VPWR _04195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14198__332 clknet_1_0__leaf__08504_ VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__inv_2
X_09020_ CPU.aluIn1\[23\] _05371_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18218_ net1229 _01746_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19198_ net57 net56 VGND VGND VPWR VPWR mapped_spi_ram.div_counter\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18149_ net1160 _01677_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold202 mapped_spi_flash.cmd_addr\[19\] VGND VGND VPWR VPWR net1499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 per_uart.uart0.txd_reg\[5\] VGND VGND VPWR VPWR net1510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 mapped_spi_flash.cmd_addr\[5\] VGND VGND VPWR VPWR net1521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 per_uart.uart0.txd_reg\[2\] VGND VGND VPWR VPWR net1532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 CPU.cycles\[8\] VGND VGND VPWR VPWR net1543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold257 _08286_ VGND VGND VPWR VPWR net1554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 CPU.cycles\[24\] VGND VGND VPWR VPWR net1565 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold279 _08274_ VGND VGND VPWR VPWR net1576 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ _05321_ _06254_ VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__or2_1
X_09853_ _05328_ _06188_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__xnor2_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15593__398 clknet_1_1__leaf__08511_ VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__inv_2
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ _05764_ _06110_ _06120_ _06122_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__a211o_4
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13577__962 clknet_1_0__leaf__08443_ VGND VGND VPWR VPWR net1018 sky130_fd_sc_hd__inv_2
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13796__1160 clknet_1_1__leaf__08464_ VGND VGND VPWR VPWR net1216 sky130_fd_sc_hd__inv_2
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09218_ CPU.aluIn1\[6\] CPU.Bimm\[6\] VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__xnor2_1
X_10490_ _06708_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09149_ _05386_ _05499_ _05500_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12160_ mapped_spi_ram.cmd_addr\[11\] _07091_ _07724_ VGND VGND VPWR VPWR _07735_
+ sky130_fd_sc_hd__mux2_1
X_11111_ _07134_ VGND VGND VPWR VPWR _07135_ sky130_fd_sc_hd__clkbuf_2
X_12091_ mapped_spi_flash.div_counter\[0\] _07198_ _06855_ VGND VGND VPWR VPWR _07686_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_102_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15953__690 clknet_1_1__leaf__03690_ VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__inv_2
Xhold780 CPU.registerFile\[19\]\[0\] VGND VGND VPWR VPWR net2077 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold791 CPU.registerFile\[17\]\[31\] VGND VGND VPWR VPWR net2088 sky130_fd_sc_hd__dlygate4sd3_1
X_11042_ _07048_ _07080_ VGND VGND VPWR VPWR _07081_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14801_ CPU.registerFile\[2\]\[11\] CPU.registerFile\[3\]\[11\] _02871_ VGND VGND
+ VPWR VPWR _02872_ sky130_fd_sc_hd__mux2_1
X_12993_ net2190 _07347_ _08192_ VGND VGND VPWR VPWR _08200_ sky130_fd_sc_hd__mux2_1
X_17520_ _05092_ _05093_ _05058_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__a21oi_1
X_14732_ CPU.registerFile\[21\]\[10\] _08718_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__or2_1
X_11944_ _06605_ net2369 _07598_ VGND VGND VPWR VPWR _07603_ sky130_fd_sc_hd__mux2_1
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13680__1055 clknet_1_0__leaf__08453_ VGND VGND VPWR VPWR net1111 sky130_fd_sc_hd__inv_2
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17451_ _05035_ _05036_ _05037_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__a21oi_1
X_14663_ _08857_ _02732_ _02736_ _08661_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__a211o_1
X_11875_ _07566_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14147__286 clknet_1_0__leaf__08499_ VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__inv_2
X_16402_ _04098_ _04106_ _04110_ _04119_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__a31o_4
Xclkbuf_1_0__f__03689_ clknet_0__03689_ VGND VGND VPWR VPWR clknet_1_0__leaf__03689_
+ sky130_fd_sc_hd__clkbuf_16
X_10826_ net2656 _06908_ _06889_ VGND VGND VPWR VPWR _06909_ sky130_fd_sc_hd__mux2_1
X_17382_ per_uart.uart0.rxd_reg\[8\] _04992_ _04993_ per_uart.uart0.rxd_reg\[7\] VGND
+ VGND VPWR VPWR _05007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14594_ CPU.registerFile\[19\]\[7\] CPU.registerFile\[18\]\[7\] _06064_ VGND VGND
+ VPWR VPWR _08833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19121_ clknet_leaf_2_clk _02641_ VGND VGND VPWR VPWR CPU.PC\[3\] sky130_fd_sc_hd__dfxtp_2
X_16333_ _03692_ _04033_ _04052_ _03601_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10757_ _05703_ VGND VGND VPWR VPWR _06853_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19052_ net794 _02572_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16264_ _05689_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__clkbuf_4
X_13476_ _08429_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10688_ _06815_ VGND VGND VPWR VPWR _06816_ sky130_fd_sc_hd__buf_4
XFILLER_0_113_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18003_ net1014 _01531_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12427_ net1932 _07339_ _07895_ VGND VGND VPWR VPWR _07899_ sky130_fd_sc_hd__mux2_1
X_15215_ CPU.registerFile\[2\]\[21\] CPU.registerFile\[3\]\[21\] _03275_ VGND VGND
+ VPWR VPWR _03276_ sky130_fd_sc_hd__mux2_1
X_16195_ _03702_ _03914_ _03917_ _03803_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__a211o_1
XFILLER_0_22_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12358_ _07862_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15146_ CPU.registerFile\[21\]\[20\] _02960_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__or2_1
X_11309_ net2257 _06054_ _07249_ VGND VGND VPWR VPWR _07250_ sky130_fd_sc_hd__mux2_1
X_15735__526 clknet_1_1__leaf__03651_ VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__inv_2
X_15077_ CPU.registerFile\[8\]\[18\] _03018_ _03140_ _02864_ VGND VGND VPWR VPWR _03141_
+ sky130_fd_sc_hd__o211a_1
X_12289_ net1459 _07812_ _07819_ _07809_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__o211a_1
X_18905_ net679 _02425_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_18836_ clknet_leaf_6_clk _02360_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_18767_ net556 _02291_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[29\] sky130_fd_sc_hd__dfxtp_1
X_15979_ CPU.registerFile\[15\]\[0\] CPU.registerFile\[14\]\[0\] _03705_ VGND VGND
+ VPWR VPWR _03706_ sky130_fd_sc_hd__mux2_1
X_13761__1129 clknet_1_1__leaf__08460_ VGND VGND VPWR VPWR net1185 sky130_fd_sc_hd__inv_2
XFILLER_0_89_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18698_ net487 _02222_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_bitcount\[5\] sky130_fd_sc_hd__dfxtp_1
X_17649_ per_uart.uart0.rx_count16\[1\] per_uart.uart0.rx_count16\[0\] VGND VGND VPWR
+ VPWR _05187_ sky130_fd_sc_hd__nand2_1
X_15629__431 clknet_1_0__leaf__03640_ VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__inv_2
XFILLER_0_93_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09003_ CPU.aluIn1\[18\] _05353_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09905_ _05855_ _05550_ _05790_ CPU.cycles\[13\] _06238_ VGND VGND VPWR VPWR _06239_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14252__381 clknet_1_1__leaf__08509_ VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__inv_2
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09836_ _06171_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__clkbuf_4
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09767_ net2328 _06106_ _06055_ VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _05369_ _05521_ _05748_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__o21a_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13358__853 clknet_1_0__leaf__08368_ VGND VGND VPWR VPWR net909 sky130_fd_sc_hd__inv_2
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11660_ _05739_ _05738_ _05737_ VGND VGND VPWR VPWR _07451_ sky130_fd_sc_hd__or3b_4
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10611_ _06772_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__clkbuf_1
X_11591_ _05735_ _05736_ CPU.writeBack VGND VGND VPWR VPWR _07414_ sky130_fd_sc_hd__nand3_4
XFILLER_0_135_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10542_ _06735_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10473_ _06698_ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15000_ _03064_ _03065_ _03025_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__mux2_1
X_12212_ _07670_ _07671_ _07771_ _07749_ VGND VGND VPWR VPWR _07772_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13192_ CPU.cycles\[30\] _08305_ VGND VGND VPWR VPWR _08308_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12143_ net1412 _07714_ _07723_ _07713_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12074_ CPU.mem_wmask\[1\] CPU.mem_wmask\[0\] CPU.mem_wmask\[3\] CPU.mem_wmask\[2\]
+ VGND VGND VPWR VPWR _07673_ sky130_fd_sc_hd__or4_4
X_16951_ _03847_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__clkbuf_4
X_11025_ _07023_ _07064_ _07065_ _06853_ VGND VGND VPWR VPWR _07066_ sky130_fd_sc_hd__o211a_1
X_16882_ CPU.registerFile\[10\]\[21\] CPU.registerFile\[11\]\[21\] _04335_ VGND VGND
+ VPWR VPWR _04588_ sky130_fd_sc_hd__mux2_1
X_18621_ net442 _02145_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_15833_ clknet_1_0__leaf__03654_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__buf_1
X_18552_ net373 _02076_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_15764_ clknet_1_1__leaf__03654_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__buf_1
X_12976_ net2323 _07330_ _08181_ VGND VGND VPWR VPWR _08191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17503_ _05075_ _05025_ _06195_ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__o21bai_1
X_14715_ _02786_ _02787_ _08783_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__mux2_1
X_18483_ net304 _02007_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_11927_ _07593_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__clkbuf_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ _05016_ CPU.PC\[2\] _05021_ _05023_ _07002_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__o221a_1
X_14646_ CPU.registerFile\[28\]\[8\] CPU.registerFile\[29\]\[8\] _08538_ VGND VGND
+ VPWR VPWR _02720_ sky130_fd_sc_hd__mux2_1
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ net2635 _07370_ _07548_ VGND VGND VPWR VPWR _07557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14080__226 clknet_1_1__leaf__08492_ VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__inv_2
XFILLER_0_55_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10809_ CPU.aluReg\[24\] _06895_ _06889_ VGND VGND VPWR VPWR _06896_ sky130_fd_sc_hd__mux2_1
X_17365_ _04995_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_19 _04662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14577_ _08815_ _08816_ _08695_ VGND VGND VPWR VPWR _08817_ sky130_fd_sc_hd__mux2_1
X_11789_ _07520_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19104_ net87 _02624_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16316_ _04034_ _04035_ _03875_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17296_ clknet_1_0__leaf__03686_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__buf_1
XFILLER_0_125_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19035_ net777 _02555_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__08461_ clknet_0__08461_ VGND VGND VPWR VPWR clknet_1_1__leaf__08461_
+ sky130_fd_sc_hd__clkbuf_16
X_16247_ _03957_ _03968_ _08406_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__o21a_1
X_13459_ _06396_ VGND VGND VPWR VPWR _08418_ sky130_fd_sc_hd__buf_6
XFILLER_0_88_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__08492_ _08492_ VGND VGND VPWR VPWR clknet_0__08492_ sky130_fd_sc_hd__clkbuf_16
X_16178_ _03713_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__clkbuf_4
X_15659__457 clknet_1_0__leaf__03644_ VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__inv_2
XFILLER_0_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13608__991 clknet_1_1__leaf__08445_ VGND VGND VPWR VPWR net1047 sky130_fd_sc_hd__inv_2
X_15129_ _03190_ _03191_ _03025_ VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09621_ _05949_ _05963_ _05964_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__a21o_1
X_18819_ net608 _02343_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_09552_ _05372_ _05521_ _05748_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__o21ai_1
X_09483_ _05809_ _05814_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18574__31 VGND VGND VPWR VPWR _18574__31/HI net31 sky130_fd_sc_hd__conb_1
XFILLER_0_19_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13938__98 clknet_1_0__leaf__08478_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__inv_2
XFILLER_0_30_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09819_ _05890_ _06155_ VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_0__f__08481_ clknet_0__08481_ VGND VGND VPWR VPWR clknet_1_0__leaf__08481_
+ sky130_fd_sc_hd__clkbuf_16
X_12830_ _05825_ net2279 _08109_ VGND VGND VPWR VPWR _08114_ sky130_fd_sc_hd__mux2_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _08064_ VGND VGND VPWR VPWR _08076_ sky130_fd_sc_hd__buf_4
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ CPU.registerFile\[5\]\[4\] CPU.registerFile\[4\]\[4\] _08576_ VGND VGND VPWR
+ VPWR _08742_ sky130_fd_sc_hd__mux2_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _07479_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _08039_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__clkbuf_1
X_15480_ CPU.registerFile\[16\]\[29\] _08527_ _03532_ _08530_ VGND VGND VPWR VPWR
+ _03533_ sky130_fd_sc_hd__o211a_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _07442_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__clkbuf_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14431_ CPU.registerFile\[19\]\[3\] CPU.registerFile\[18\]\[3\] _06064_ VGND VGND
+ VPWR VPWR _08674_ sky130_fd_sc_hd__mux2_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17150_ _04847_ _04848_ _04557_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11574_ _07405_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__clkbuf_1
X_14362_ CPU.registerFile\[30\]\[1\] CPU.registerFile\[31\]\[1\] _08536_ VGND VGND
+ VPWR VPWR _08607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16101_ _03824_ _03825_ _03720_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10525_ net2204 _06337_ _06724_ VGND VGND VPWR VPWR _06727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17081_ CPU.registerFile\[0\]\[26\] _04637_ _04472_ _04781_ VGND VGND VPWR VPWR _04782_
+ sky130_fd_sc_hd__o211a_1
X_14293_ CPU.registerFile\[28\]\[0\] CPU.registerFile\[29\]\[0\] _08538_ VGND VGND
+ VPWR VPWR _08539_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13639__1019 clknet_1_0__leaf__08448_ VGND VGND VPWR VPWR net1075 sky130_fd_sc_hd__inv_2
XFILLER_0_40_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13760__1128 clknet_1_1__leaf__08460_ VGND VGND VPWR VPWR net1184 sky130_fd_sc_hd__inv_2
X_16032_ _06172_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__buf_4
X_14259__387 clknet_1_1__leaf__08510_ VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__inv_2
X_10456_ _06643_ net2424 _06687_ VGND VGND VPWR VPWR _06690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13175_ CPU.cycles\[22\] _08295_ net1547 VGND VGND VPWR VPWR _08298_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10387_ _06649_ net1983 _06639_ VGND VGND VPWR VPWR _06650_ sky130_fd_sc_hd__mux2_1
X_12126_ mapped_spi_ram.cmd_addr\[21\] _05667_ _07704_ VGND VGND VPWR VPWR _07711_
+ sky130_fd_sc_hd__mux2_1
X_17983_ net994 _01511_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_16934_ CPU.registerFile\[0\]\[22\] _04637_ _04472_ _04638_ VGND VGND VPWR VPWR _04639_
+ sky130_fd_sc_hd__o211a_1
X_12057_ CPU.registerFile\[24\]\[6\] _07364_ _07657_ VGND VGND VPWR VPWR _07663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11008_ _07023_ _07049_ _07050_ _06853_ VGND VGND VPWR VPWR _07051_ sky130_fd_sc_hd__o211a_1
X_16865_ _04441_ _04568_ _04571_ _04208_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__a211o_1
X_18604_ net425 _02128_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_15816_ _08359_ _03676_ _03660_ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__a21oi_1
X_16796_ CPU.registerFile\[10\]\[19\] CPU.registerFile\[11\]\[19\] _04335_ VGND VGND
+ VPWR VPWR _04504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18535_ net356 _02059_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12959_ _08182_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18466_ net287 _00010_ VGND VGND VPWR VPWR mapped_spi_ram.state\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13945__104 clknet_1_1__leaf__08479_ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__inv_2
X_14629_ _08585_ _08586_ CPU.registerFile\[1\]\[7\] VGND VGND VPWR VPWR _08868_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18397_ net218 _01925_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17279_ _08397_ _04972_ _04974_ _08400_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__a211o_1
X_15893__636 clknet_1_1__leaf__03684_ VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__inv_2
XFILLER_0_130_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19018_ net760 _02538_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__08444_ clknet_0__08444_ VGND VGND VPWR VPWR clknet_1_1__leaf__08444_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__08475_ _08475_ VGND VGND VPWR VPWR clknet_0__08475_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13541__931 clknet_1_1__leaf__08438_ VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__inv_2
XFILLER_0_11_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08983_ CPU.aluIn1\[13\] _05322_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__or2_2
X_13991__146 clknet_1_0__leaf__08483_ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__inv_2
XFILLER_0_139_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09604_ CPU.Bimm\[6\] _05913_ CPU.PC\[6\] VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__a21o_1
X_09535_ _05547_ CPU.instr\[2\] _05878_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__and3b_1
XFILLER_0_149_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09466_ _05386_ _05813_ _05500_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09397_ _05747_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10310_ _06593_ net2025 _06597_ VGND VGND VPWR VPWR _06598_ sky130_fd_sc_hd__mux2_1
X_11290_ net1909 _05767_ _07238_ VGND VGND VPWR VPWR _07240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10241_ net1714 _05767_ _06558_ VGND VGND VPWR VPWR _06560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10172_ mapped_spi_ram.rcv_data\[10\] _05857_ _05859_ net1419 VGND VGND VPWR VPWR
+ _06495_ sky130_fd_sc_hd__a22o_2
XFILLER_0_100_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14980_ CPU.registerFile\[28\]\[16\] CPU.registerFile\[29\]\[16\] _02808_ VGND VGND
+ VPWR VPWR _03046_ sky130_fd_sc_hd__mux2_1
X_13931_ clknet_1_1__leaf__08473_ VGND VGND VPWR VPWR _08478_ sky130_fd_sc_hd__buf_1
X_16650_ _03736_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__buf_4
Xclkbuf_1_0__f__08464_ clknet_0__08464_ VGND VGND VPWR VPWR clknet_1_0__leaf__08464_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15688__483 clknet_1_0__leaf__03647_ VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__inv_2
X_12813_ CPU.aluShamt\[1\] CPU.aluShamt\[0\] VGND VGND VPWR VPWR _08104_ sky130_fd_sc_hd__nor2_1
X_16581_ _04285_ _04294_ _04138_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18320_ net141 _01848_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15532_ CPU.registerFile\[15\]\[30\] CPU.registerFile\[14\]\[30\] _08560_ VGND VGND
+ VPWR VPWR _03584_ sky130_fd_sc_hd__mux2_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _08067_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__clkbuf_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13256__776 clknet_1_1__leaf__08344_ VGND VGND VPWR VPWR net832 sky130_fd_sc_hd__inv_2
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ net1262 _01779_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_15463_ _08546_ _08547_ CPU.registerFile\[9\]\[28\] VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__a21o_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _06599_ net2558 _08029_ VGND VGND VPWR VPWR _08031_ sky130_fd_sc_hd__mux2_1
X_17202_ CPU.registerFile\[20\]\[29\] CPU.registerFile\[21\]\[29\] _03737_ VGND VGND
+ VPWR VPWR _04900_ sky130_fd_sc_hd__mux2_1
X_14414_ CPU.registerFile\[10\]\[2\] CPU.registerFile\[11\]\[2\] _08564_ VGND VGND
+ VPWR VPWR _08658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11626_ _07433_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__clkbuf_1
X_18182_ net1193 _01710_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[21\] sky130_fd_sc_hd__dfxtp_1
X_15394_ _03133_ _03445_ _03449_ _03188_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17133_ _04579_ _04580_ CPU.registerFile\[17\]\[27\] VGND VGND VPWR VPWR _04833_
+ sky130_fd_sc_hd__a21o_1
X_14345_ _08581_ _08583_ _08589_ _08590_ VGND VGND VPWR VPWR _08591_ sky130_fd_sc_hd__a211o_1
X_11557_ _07396_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold609 CPU.registerFile\[18\]\[7\] VGND VGND VPWR VPWR net1906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17064_ _04574_ _04761_ _04765_ _04584_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__o211a_1
X_10508_ net2239 _06145_ _06713_ VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__mux2_1
X_11488_ net1746 _07353_ _07354_ VGND VGND VPWR VPWR _07355_ sky130_fd_sc_hd__mux2_1
X_14276_ _08409_ VGND VGND VPWR VPWR _08522_ sky130_fd_sc_hd__clkbuf_8
X_13917__79 clknet_1_1__leaf__08476_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__inv_2
XFILLER_0_123_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14192__327 clknet_1_1__leaf__08503_ VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__inv_2
X_16015_ _03741_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__buf_4
X_10439_ _06626_ net2277 _06676_ VGND VGND VPWR VPWR _06681_ sky130_fd_sc_hd__mux2_1
X_13227_ clknet_1_0__leaf__08339_ VGND VGND VPWR VPWR _08340_ sky130_fd_sc_hd__buf_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ _08287_ _08288_ VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__nor2_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ net1326 _07694_ _07696_ VGND VGND VPWR VPWR _07700_ sky130_fd_sc_hd__a21o_1
X_13089_ net1363 VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__clkbuf_1
X_17966_ net977 _01494_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1309 CPU.registerFile\[1\]\[4\] VGND VGND VPWR VPWR net2606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16917_ _04614_ _04622_ _04542_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__o21a_1
X_17897_ clknet_leaf_25_clk _01425_ VGND VGND VPWR VPWR CPU.instr\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_109_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16848_ CPU.registerFile\[6\]\[20\] CPU.registerFile\[7\]\[20\] _04426_ VGND VGND
+ VPWR VPWR _04555_ sky130_fd_sc_hd__mux2_1
X_14012__164 clknet_1_1__leaf__08486_ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__inv_2
X_16779_ _04441_ _04483_ _04487_ _04208_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13571__957 clknet_1_0__leaf__08442_ VGND VGND VPWR VPWR net1013 sky130_fd_sc_hd__inv_2
XFILLER_0_87_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09320_ _05667_ _05671_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__or2_2
X_18518_ net339 _02042_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09251_ CPU.aluIn1\[9\] CPU.Bimm\[9\] VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18449_ net270 _01977_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09182_ CPU.Jimm\[13\] _05530_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__nor2_8
XFILLER_0_141_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15901__643 clknet_1_0__leaf__03685_ VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__inv_2
XFILLER_0_145_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15600__404 clknet_1_0__leaf__03638_ VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__inv_2
XFILLER_0_114_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__08458_ _08458_ VGND VGND VPWR VPWR clknet_0__08458_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08966_ CPU.aluIn1\[12\] _05317_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__and2b_1
X_17417__39 clknet_1_0__leaf__05014_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__inv_2
XFILLER_0_75_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08897_ CPU.Bimm\[12\] _05248_ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__or2_2
X_13638__1018 clknet_1_0__leaf__08448_ VGND VGND VPWR VPWR net1074 sky130_fd_sc_hd__inv_2
XFILLER_0_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09518_ _05391_ _05497_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__xor2_1
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10790_ _06880_ VGND VGND VPWR VPWR _06881_ sky130_fd_sc_hd__buf_4
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09449_ _05775_ _05794_ _05795_ _05797_ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__o31a_1
XFILLER_0_93_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12460_ net1727 _07372_ _07906_ VGND VGND VPWR VPWR _07916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11411_ _07303_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12391_ _07879_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__clkbuf_1
X_13548__937 clknet_1_1__leaf__08439_ VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__inv_2
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11342_ net2458 _06440_ _07260_ VGND VGND VPWR VPWR _07267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11273_ _06651_ net2506 _07223_ VGND VGND VPWR VPWR _07230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13012_ net2062 _07366_ _08203_ VGND VGND VPWR VPWR _08210_ sky130_fd_sc_hd__mux2_1
X_10224_ _05417_ _06544_ _05419_ VGND VGND VPWR VPWR _06545_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_120_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17820_ net900 _01382_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_10155_ _05443_ _05433_ _05441_ _06478_ VGND VGND VPWR VPWR _06479_ sky130_fd_sc_hd__a31o_1
X_17751_ net836 _01317_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold6 _07835_ VGND VGND VPWR VPWR net1303 sky130_fd_sc_hd__clkbuf_2
X_14963_ CPU.registerFile\[0\]\[15\] _02948_ _03029_ _02791_ VGND VGND VPWR VPWR _03030_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10086_ _06412_ VGND VGND VPWR VPWR _06413_ sky130_fd_sc_hd__buf_4
XFILLER_0_89_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16702_ _04403_ _04412_ _04138_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__o21a_1
X_17682_ CPU.mem_wdata\[0\] per_uart.uart0.rx_ack _05211_ VGND VGND VPWR VPWR _05212_
+ sky130_fd_sc_hd__mux2_1
X_14894_ CPU.registerFile\[20\]\[14\] _08839_ _02961_ _08841_ VGND VGND VPWR VPWR
+ _02962_ sky130_fd_sc_hd__o211a_1
X_16633_ CPU.registerFile\[5\]\[15\] CPU.registerFile\[4\]\[15\] _04024_ VGND VGND
+ VPWR VPWR _04345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__08447_ clknet_0__08447_ VGND VGND VPWR VPWR clknet_1_0__leaf__08447_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_947 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16564_ CPU.registerFile\[28\]\[13\] CPU.registerFile\[29\]\[13\] _04122_ VGND VGND
+ VPWR VPWR _04278_ sky130_fd_sc_hd__mux2_1
X_13776_ clknet_1_0__leaf__08462_ VGND VGND VPWR VPWR _08463_ sky130_fd_sc_hd__buf_1
X_10988_ mapped_spi_flash.cmd_addr\[14\] _07033_ _07009_ VGND VGND VPWR VPWR _07034_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18303_ net124 _01831_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_15515_ CPU.registerFile\[19\]\[30\] CPU.registerFile\[18\]\[30\] _06456_ VGND VGND
+ VPWR VPWR _03567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12727_ _06651_ net2628 _08051_ VGND VGND VPWR VPWR _08058_ sky130_fd_sc_hd__mux2_1
X_16495_ CPU.registerFile\[22\]\[11\] CPU.registerFile\[23\]\[11\] _03958_ VGND VGND
+ VPWR VPWR _04211_ sky130_fd_sc_hd__mux2_1
X_18234_ net1245 net18 VGND VGND VPWR VPWR mapped_spi_flash.div_counter\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15446_ CPU.registerFile\[22\]\[28\] CPU.registerFile\[23\]\[28\] _08584_ VGND VGND
+ VPWR VPWR _03500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12658_ _08021_ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11609_ _07424_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__clkbuf_1
X_18165_ net1176 _01693_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15377_ _03078_ _03430_ _03432_ _08535_ VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__a211o_1
XFILLER_0_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12589_ net2541 _07364_ _07979_ VGND VGND VPWR VPWR _07985_ sky130_fd_sc_hd__mux2_1
X_14200__334 clknet_1_0__leaf__08504_ VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__inv_2
XFILLER_0_26_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_16
X_17116_ _03748_ _03750_ CPU.registerFile\[1\]\[27\] VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14328_ _06013_ VGND VGND VPWR VPWR _08574_ sky130_fd_sc_hd__clkbuf_4
X_18096_ net1107 _01624_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold406 CPU.registerFile\[27\]\[28\] VGND VGND VPWR VPWR net1703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold417 CPU.registerFile\[19\]\[30\] VGND VGND VPWR VPWR net1714 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold428 CPU.registerFile\[3\]\[30\] VGND VGND VPWR VPWR net1725 sky130_fd_sc_hd__dlygate4sd3_1
X_17047_ _03757_ _04744_ _04748_ _04476_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold439 CPU.registerFile\[5\]\[5\] VGND VGND VPWR VPWR net1736 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__03685_ clknet_0__03685_ VGND VGND VPWR VPWR clknet_1_1__leaf__03685_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18998_ clknet_leaf_12_clk _02518_ VGND VGND VPWR VPWR CPU.aluIn1\[15\] sky130_fd_sc_hd__dfxtp_2
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 CPU.registerFile\[30\]\[6\] VGND VGND VPWR VPWR net2403 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 CPU.registerFile\[23\]\[10\] VGND VGND VPWR VPWR net2414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1128 CPU.registerFile\[16\]\[8\] VGND VGND VPWR VPWR net2425 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17949_ net960 _01477_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[19\] sky130_fd_sc_hd__dfxtp_1
Xhold1139 CPU.registerFile\[1\]\[10\] VGND VGND VPWR VPWR net2436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09303_ _05653_ _05654_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15825__574 clknet_1_0__leaf__03678_ VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__inv_2
X_13352__848 clknet_1_0__leaf__08367_ VGND VGND VPWR VPWR net904 sky130_fd_sc_hd__inv_2
XFILLER_0_35_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09234_ CPU.Iimm\[4\] CPU.Bimm\[4\] CPU.instr\[5\] VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09165_ _05516_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09096_ _05429_ _05447_ _05296_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_31_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold940 CPU.registerFile\[7\]\[20\] VGND VGND VPWR VPWR net2237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold951 CPU.registerFile\[7\]\[7\] VGND VGND VPWR VPWR net2248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 CPU.registerFile\[8\]\[25\] VGND VGND VPWR VPWR net2259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold973 CPU.registerFile\[8\]\[0\] VGND VGND VPWR VPWR net2270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold984 CPU.registerFile\[26\]\[19\] VGND VGND VPWR VPWR net2281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 CPU.registerFile\[7\]\[0\] VGND VGND VPWR VPWR net2292 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09998_ _06327_ _05971_ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__xnor2_1
X_08949_ _05296_ _05300_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11960_ _07611_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10911_ _06854_ VGND VGND VPWR VPWR _06973_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11891_ _06620_ net2268 _07573_ VGND VGND VPWR VPWR _07575_ sky130_fd_sc_hd__mux2_1
X_10842_ CPU.aluIn1\[16\] _06920_ _06914_ VGND VGND VPWR VPWR _06921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10773_ CPU.aluWr _05770_ VGND VGND VPWR VPWR _06867_ sky130_fd_sc_hd__nand2_1
X_15300_ _03156_ _03355_ _03357_ _03163_ VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__a211o_1
X_12512_ net1802 _07356_ _07942_ VGND VGND VPWR VPWR _07944_ sky130_fd_sc_hd__mux2_1
X_16280_ CPU.registerFile\[20\]\[6\] CPU.registerFile\[21\]\[6\] _03883_ VGND VGND
+ VPWR VPWR _04001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15231_ _08409_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__buf_4
XFILLER_0_125_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12443_ _07907_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15162_ _03222_ _03223_ _02937_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__mux2_1
X_12374_ _06638_ net2304 _07870_ VGND VGND VPWR VPWR _07871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13329__828 clknet_1_1__leaf__08364_ VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__inv_2
X_11325_ net2080 _06245_ _07249_ VGND VGND VPWR VPWR _07258_ sky130_fd_sc_hd__mux2_1
X_15093_ _08414_ VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__clkbuf_4
X_11256_ _06634_ net1987 _07212_ VGND VGND VPWR VPWR _07221_ sky130_fd_sc_hd__mux2_1
X_18921_ net695 _02441_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_13874__1231 clknet_1_0__leaf__08471_ VGND VGND VPWR VPWR net1287 sky130_fd_sc_hd__inv_2
XFILLER_0_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10207_ CPU.cycles\[1\] _05759_ _06515_ _06518_ _06528_ VGND VGND VPWR VPWR _06529_
+ sky130_fd_sc_hd__a2111o_1
X_11187_ net7 _07178_ _06855_ VGND VGND VPWR VPWR _07179_ sky130_fd_sc_hd__o21a_1
X_18852_ net626 _00005_ VGND VGND VPWR VPWR mapped_spi_flash.state\[1\] sky130_fd_sc_hd__dfxtp_4
X_10138_ _05855_ _06459_ _06461_ _06462_ _06176_ VGND VGND VPWR VPWR _06463_ sky130_fd_sc_hd__o221a_1
X_17803_ net883 _01365_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_18783_ net572 _02307_ VGND VGND VPWR VPWR CPU.aluReg\[13\] sky130_fd_sc_hd__dfxtp_1
X_15995_ _08396_ VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__buf_4
X_17734_ net819 _01300_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_14946_ _06061_ VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__buf_4
X_10069_ mapped_spi_ram.rcv_data\[14\] _05857_ _05859_ mapped_spi_flash.rcv_data\[14\]
+ VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__a22o_4
X_17665_ per_uart.uart0.rx_bitcount\[1\] _05195_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__nand2_1
X_14877_ _02944_ _02945_ _08783_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16616_ _04175_ _04176_ CPU.registerFile\[17\]\[14\] VGND VGND VPWR VPWR _04329_
+ sky130_fd_sc_hd__a21o_1
X_17596_ _05237_ net1585 VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16547_ CPU.registerFile\[9\]\[13\] _04056_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16478_ _04192_ _04193_ _04153_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14124__265 clknet_1_0__leaf__08497_ VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__inv_2
X_18217_ net1228 net1413 VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[18\] sky130_fd_sc_hd__dfxtp_1
X_15429_ _08543_ _03481_ _03483_ _03307_ VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19197_ net107 net55 VGND VGND VPWR VPWR mapped_spi_ram.div_counter\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18148_ net1159 _01676_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold203 per_uart.uart0.enable16_counter\[0\] VGND VGND VPWR VPWR net1500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 _02678_ VGND VGND VPWR VPWR net1511 sky130_fd_sc_hd__dlygate4sd3_1
X_13637__1017 clknet_1_0__leaf__08448_ VGND VGND VPWR VPWR net1073 sky130_fd_sc_hd__inv_2
XFILLER_0_123_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18079_ net1090 _01607_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[21\] sky130_fd_sc_hd__dfxtp_1
Xhold225 mapped_spi_flash.cmd_addr\[13\] VGND VGND VPWR VPWR net1522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 _02675_ VGND VGND VPWR VPWR net1533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _08278_ VGND VGND VPWR VPWR net1544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 mapped_spi_flash.snd_bitcount\[5\] VGND VGND VPWR VPWR net1555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 mapped_spi_ram.rcv_data\[16\] VGND VGND VPWR VPWR net1566 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _05320_ _06253_ VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ _05334_ _06187_ _05331_ VGND VGND VPWR VPWR _06188_ sky130_fd_sc_hd__a21oi_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15712__505 clknet_1_0__leaf__03649_ VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__inv_2
X_14018__170 clknet_1_0__leaf__08486_ VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__inv_2
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _05912_ _06121_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__nor2_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15606__410 clknet_1_1__leaf__03638_ VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__inv_2
XFILLER_0_118_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09217_ CPU.aluIn1\[6\] CPU.Bimm\[6\] _05568_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__nand3_1
XFILLER_0_72_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09148_ _05383_ CPU.aluIn1\[25\] VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__and2b_1
XFILLER_0_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09079_ _05287_ CPU.aluIn1\[4\] VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__or2b_1
XFILLER_0_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11110_ _07129_ _07131_ VGND VGND VPWR VPWR _07134_ sky130_fd_sc_hd__and2_2
XFILLER_0_102_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12090_ _07685_ VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__clkbuf_1
Xhold770 CPU.registerFile\[21\]\[2\] VGND VGND VPWR VPWR net2067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 CPU.registerFile\[26\]\[11\] VGND VGND VPWR VPWR net2078 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ mapped_spi_flash.cmd_addr\[7\] _07079_ _07039_ VGND VGND VPWR VPWR _07080_
+ sky130_fd_sc_hd__mux2_1
Xhold792 CPU.registerFile\[23\]\[9\] VGND VGND VPWR VPWR net2089 sky130_fd_sc_hd__dlygate4sd3_1
X_14800_ _08525_ VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__buf_4
X_12992_ _08199_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__clkbuf_1
X_14731_ CPU.registerFile\[22\]\[10\] CPU.registerFile\[23\]\[10\] _08756_ VGND VGND
+ VPWR VPWR _02803_ sky130_fd_sc_hd__mux2_1
X_11943_ _07602_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__clkbuf_1
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _08255_ net2388 _06973_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__o21ai_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ CPU.registerFile\[8\]\[8\] _08776_ _02735_ _08622_ VGND VGND VPWR VPWR _02736_
+ sky130_fd_sc_hd__o211a_1
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ _06603_ net2209 _07562_ VGND VGND VPWR VPWR _07566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _03901_ _04113_ _04118_ _04072_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_0__f__03688_ clknet_0__03688_ VGND VGND VPWR VPWR clknet_1_0__leaf__03688_
+ sky130_fd_sc_hd__clkbuf_16
X_10825_ CPU.aluIn1\[20\] _06907_ _06881_ VGND VGND VPWR VPWR _06908_ sky130_fd_sc_hd__mux2_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17381_ _05006_ VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14593_ CPU.mem_wdata\[6\] _08514_ _08832_ _08751_ VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19120_ clknet_leaf_10_clk _02640_ VGND VGND VPWR VPWR CPU.PC\[2\] sky130_fd_sc_hd__dfxtp_2
X_16332_ _04043_ _04051_ _08406_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10756_ mapped_spi_flash.state\[2\] net1652 VGND VGND VPWR VPWR _06852_ sky130_fd_sc_hd__or2b_1
XFILLER_0_153_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19051_ net793 _02571_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16263_ CPU.registerFile\[2\]\[6\] CPU.registerFile\[3\]\[6\] _03693_ VGND VGND VPWR
+ VPWR _03984_ sky130_fd_sc_hd__mux2_1
X_13475_ CPU.Bimm\[7\] _05822_ _08416_ VGND VGND VPWR VPWR _08429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10687_ _06813_ _06814_ VGND VGND VPWR VPWR _06815_ sky130_fd_sc_hd__nor2b_4
X_18002_ net1013 _01530_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15214_ _08525_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__buf_4
X_12426_ _07898_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__clkbuf_1
X_16194_ CPU.registerFile\[24\]\[4\] _03915_ _03747_ _03916_ VGND VGND VPWR VPWR _03917_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15145_ CPU.registerFile\[22\]\[20\] CPU.registerFile\[23\]\[20\] _02998_ VGND VGND
+ VPWR VPWR _03207_ sky130_fd_sc_hd__mux2_1
X_12357_ _06622_ net2446 _07859_ VGND VGND VPWR VPWR _07862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11308_ _07237_ VGND VGND VPWR VPWR _07249_ sky130_fd_sc_hd__buf_4
X_15076_ _03138_ _03139_ CPU.registerFile\[9\]\[18\] VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__a21o_1
X_12288_ mapped_spi_ram.rcv_data\[6\] _07813_ VGND VGND VPWR VPWR _07819_ sky130_fd_sc_hd__or2_1
X_18904_ net678 _02424_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_13381__874 clknet_1_1__leaf__08370_ VGND VGND VPWR VPWR net930 sky130_fd_sc_hd__inv_2
X_11239_ _07200_ VGND VGND VPWR VPWR _07212_ sky130_fd_sc_hd__buf_4
X_18835_ net624 _02359_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_15978_ _03704_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__buf_4
X_18766_ net555 _02290_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14929_ CPU.registerFile\[16\]\[15\] _02755_ _02995_ _02757_ VGND VGND VPWR VPWR
+ _02996_ sky130_fd_sc_hd__o211a_1
X_18697_ net486 net1447 VGND VGND VPWR VPWR mapped_spi_flash.rcv_bitcount\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17648_ net2622 _05185_ _05186_ _03659_ _06858_ VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__o221a_1
X_17579_ per_uart.uart0.tx_count16\[3\] _03659_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14206__340 clknet_1_1__leaf__08504_ VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__inv_2
XFILLER_0_85_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09002_ CPU.aluIn1\[18\] _05353_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15937__675 clknet_1_1__leaf__03689_ VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__inv_2
XFILLER_0_111_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09904_ _05910_ _06235_ _06237_ _05881_ VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09835_ _05689_ _05690_ VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__nand2_8
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09766_ _06105_ VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__buf_4
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09697_ CPU.PC\[21\] _05893_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__xnor2_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13873__1230 clknet_1_0__leaf__08471_ VGND VGND VPWR VPWR net1286 sky130_fd_sc_hd__inv_2
X_10610_ net2161 _06530_ _06738_ VGND VGND VPWR VPWR _06772_ sky130_fd_sc_hd__mux2_1
X_15682__478 clknet_1_1__leaf__03646_ VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__inv_2
X_17324__737 clknet_1_1__leaf__04982_ VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__inv_2
X_11590_ _07413_ VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10541_ net2049 _06530_ _06701_ VGND VGND VPWR VPWR _06735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10472_ _06659_ net2331 _06664_ VGND VGND VPWR VPWR _06698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12211_ mapped_spi_ram.snd_bitcount\[3\] _07770_ _07758_ VGND VGND VPWR VPWR _07771_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13191_ CPU.cycles\[30\] _08305_ VGND VGND VPWR VPWR _08307_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12142_ _07715_ _07722_ VGND VGND VPWR VPWR _07723_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12073_ net1307 VGND VGND VPWR VPWR _07672_ sky130_fd_sc_hd__inv_2
X_16950_ CPU.registerFile\[19\]\[22\] CPU.registerFile\[18\]\[22\] _04327_ VGND VGND
+ VPWR VPWR _04655_ sky130_fd_sc_hd__mux2_1
X_11024_ CPU.PC\[10\] _05643_ VGND VGND VPWR VPWR _07065_ sky130_fd_sc_hd__or2_1
X_16881_ CPU.aluIn1\[20\] _04458_ _04587_ _04259_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__o211a_1
X_18620_ net441 _02144_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_15763_ clknet_1_1__leaf__08339_ VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__buf_1
X_18551_ net372 _02075_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_12975_ _08190_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14714_ CPU.registerFile\[5\]\[9\] CPU.registerFile\[4\]\[9\] _08864_ VGND VGND VPWR
+ VPWR _02787_ sky130_fd_sc_hd__mux2_1
X_17502_ _05069_ CPU.PC\[14\] _05078_ _05079_ _05053_ VGND VGND VPWR VPWR _02652_
+ sky130_fd_sc_hd__o221a_1
X_18482_ net303 _02006_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11926_ _06655_ net1830 _07584_ VGND VGND VPWR VPWR _07593_ sky130_fd_sc_hd__mux2_1
X_13636__1016 clknet_1_0__leaf__08448_ VGND VGND VPWR VPWR net1072 sky130_fd_sc_hd__inv_2
XFILLER_0_86_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _05022_ _06498_ _08256_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__o21ai_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ CPU.registerFile\[30\]\[8\] CPU.registerFile\[31\]\[8\] _08645_ VGND VGND
+ VPWR VPWR _02719_ sky130_fd_sc_hd__mux2_1
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _07556_ VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__clkbuf_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10808_ CPU.aluIn1\[24\] _06894_ _06881_ VGND VGND VPWR VPWR _06895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17364_ _06992_ _04994_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__and2_1
X_14576_ CPU.registerFile\[13\]\[6\] CPU.registerFile\[12\]\[6\] _08693_ VGND VGND
+ VPWR VPWR _08816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11788_ _06653_ net2024 _07512_ VGND VGND VPWR VPWR _07520_ sky130_fd_sc_hd__mux2_1
X_16315_ CPU.registerFile\[28\]\[7\] CPU.registerFile\[29\]\[7\] _03739_ VGND VGND
+ VPWR VPWR _04035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19103_ net86 _02623_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_17299__714 clknet_1_0__leaf__04980_ VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__inv_2
X_10739_ net2238 _06386_ _06838_ VGND VGND VPWR VPWR _06843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19034_ net776 _02554_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_16246_ _03758_ _03962_ _03967_ _03775_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__08460_ clknet_0__08460_ VGND VGND VPWR VPWR clknet_1_1__leaf__08460_
+ sky130_fd_sc_hd__clkbuf_16
X_13458_ _08417_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__08491_ _08491_ VGND VGND VPWR VPWR clknet_0__08491_ sky130_fd_sc_hd__clkbuf_16
X_12409_ _07889_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__clkbuf_1
X_16177_ _03703_ _03897_ _03899_ _03714_ VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__a211o_1
XFILLER_0_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13389_ _06390_ _06391_ _08372_ VGND VGND VPWR VPWR _08373_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15128_ CPU.registerFile\[5\]\[19\] CPU.registerFile\[4\]\[19\] _03105_ VGND VGND
+ VPWR VPWR _03191_ sky130_fd_sc_hd__mux2_1
X_14236__366 clknet_1_1__leaf__08508_ VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__inv_2
X_15059_ _03078_ _03120_ _03122_ _03043_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__a211o_1
X_09620_ CPU.PC\[5\] CPU.Bimm\[5\] _05913_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__and3_1
X_18818_ net607 _02342_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09551_ CPU.PC\[23\] _05894_ VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__xnor2_1
X_18749_ net538 net1498 VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09482_ _05399_ _05521_ _05748_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15870__615 clknet_1_0__leaf__03682_ VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__inv_2
XFILLER_0_100_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15718__511 clknet_1_1__leaf__03649_ VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__inv_2
XFILLER_0_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09818_ CPU.PC\[15\] _05889_ CPU.PC\[16\] VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_1_0__f__08480_ clknet_0__08480_ VGND VGND VPWR VPWR clknet_1_0__leaf__08480_
+ sky130_fd_sc_hd__clkbuf_16
X_09749_ _05349_ _05521_ _05748_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__o21a_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _08075_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__clkbuf_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ net2353 _07360_ _07475_ VGND VGND VPWR VPWR _07479_ sky130_fd_sc_hd__mux2_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _06615_ net2536 _08029_ VGND VGND VPWR VPWR _08039_ sky130_fd_sc_hd__mux2_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ CPU.mem_wdata\[2\] _08514_ _08673_ _07822_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__o211a_1
X_11642_ net2034 _07360_ _07438_ VGND VGND VPWR VPWR _07442_ sky130_fd_sc_hd__mux2_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14361_ _08521_ _08603_ _08605_ _08533_ VGND VGND VPWR VPWR _08606_ sky130_fd_sc_hd__a211o_1
X_11573_ net1720 _07360_ _07401_ VGND VGND VPWR VPWR _07405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16100_ CPU.registerFile\[5\]\[2\] CPU.registerFile\[4\]\[2\] _03704_ VGND VGND VPWR
+ VPWR _03825_ sky130_fd_sc_hd__mux2_1
X_17080_ _03748_ _03750_ CPU.registerFile\[1\]\[26\] VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__a21o_1
X_10524_ _06726_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__clkbuf_1
X_14292_ _08409_ VGND VGND VPWR VPWR _08538_ sky130_fd_sc_hd__buf_4
XFILLER_0_107_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16031_ _03757_ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10455_ _06689_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13174_ CPU.cycles\[22\] CPU.cycles\[23\] _08295_ VGND VGND VPWR VPWR _08297_ sky130_fd_sc_hd__and3_1
X_10386_ _06412_ VGND VGND VPWR VPWR _06649_ sky130_fd_sc_hd__clkbuf_8
X_12125_ net1425 _07693_ _07710_ _07175_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__o211a_1
X_17982_ net993 _01510_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_16933_ _04389_ _04390_ CPU.registerFile\[1\]\[22\] VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__a21o_1
X_12056_ _07662_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11007_ CPU.PC\[12\] _07031_ VGND VGND VPWR VPWR _07050_ sky130_fd_sc_hd__or2_1
X_16864_ CPU.registerFile\[24\]\[20\] _04319_ _04569_ _04570_ VGND VGND VPWR VPWR
+ _04571_ sky130_fd_sc_hd__o211a_1
X_18603_ net424 _02127_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15815_ net1598 _08357_ net1603 VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__o21ai_1
X_16795_ _08397_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18534_ net355 _02058_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12958_ net1882 _07309_ _08181_ VGND VGND VPWR VPWR _08182_ sky130_fd_sc_hd__mux2_1
X_11909_ _07561_ VGND VGND VPWR VPWR _07584_ sky130_fd_sc_hd__buf_4
X_18465_ net286 _00009_ VGND VGND VPWR VPWR mapped_spi_ram.state\[1\] sky130_fd_sc_hd__dfxtp_1
X_12889_ _08144_ VGND VGND VPWR VPWR _08145_ sky130_fd_sc_hd__buf_4
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15665__462 clknet_1_0__leaf__03645_ VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__inv_2
X_14628_ CPU.registerFile\[2\]\[7\] CPU.registerFile\[3\]\[7\] _08629_ VGND VGND VPWR
+ VPWR _08867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18396_ net217 _01924_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14559_ CPU.registerFile\[22\]\[6\] CPU.registerFile\[23\]\[6\] _08756_ VGND VGND
+ VPWR VPWR _08799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13233__755 clknet_1_1__leaf__08342_ VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__inv_2
XFILLER_0_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17278_ CPU.registerFile\[16\]\[31\] _04656_ _06149_ _04973_ VGND VGND VPWR VPWR
+ _04974_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19017_ net759 _02537_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_16229_ CPU.registerFile\[28\]\[5\] CPU.registerFile\[29\]\[5\] _03739_ VGND VGND
+ VPWR VPWR _03951_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__08443_ clknet_0__08443_ VGND VGND VPWR VPWR clknet_1_1__leaf__08443_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__08474_ _08474_ VGND VGND VPWR VPWR clknet_0__08474_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08982_ _05333_ VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__inv_2
X_09603_ CPU.Bimm\[7\] _05913_ CPU.PC\[7\] VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09534_ CPU.instr\[4\] CPU.instr\[6\] _05422_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__and3b_1
XFILLER_0_94_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09465_ _05391_ _05497_ _05499_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__a21o_1
X_14063__211 clknet_1_1__leaf__08490_ VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__inv_2
XFILLER_0_149_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09396_ _05746_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_47_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10240_ _06559_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13635__1015 clknet_1_1__leaf__08448_ VGND VGND VPWR VPWR net1071 sky130_fd_sc_hd__inv_2
X_10171_ _05691_ _06311_ VGND VGND VPWR VPWR _06494_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_0__f__08463_ clknet_0__08463_ VGND VGND VPWR VPWR clknet_1_0__leaf__08463_
+ sky130_fd_sc_hd__clkbuf_16
X_12812_ _05268_ _06861_ _08102_ _08103_ _06869_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__o221a_1
X_16580_ _04170_ _04289_ _04293_ _04180_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__o211a_1
X_15531_ _08592_ _03570_ _03574_ _03582_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _06599_ net2538 _08065_ VGND VGND VPWR VPWR _08067_ sky130_fd_sc_hd__mux2_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14265__392 clknet_1_0__leaf__08511_ VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__inv_2
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ net1261 _01778_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_15462_ CPU.registerFile\[10\]\[28\] CPU.registerFile\[11\]\[28\] _03183_ VGND VGND
+ VPWR VPWR _03516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _08030_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ CPU.registerFile\[22\]\[29\] CPU.registerFile\[23\]\[29\] _03761_ VGND VGND
+ VPWR VPWR _04899_ sky130_fd_sc_hd__mux2_1
X_14413_ _08655_ _08656_ _08562_ VGND VGND VPWR VPWR _08657_ sky130_fd_sc_hd__mux2_1
X_11625_ net2390 _07343_ _07427_ VGND VGND VPWR VPWR _07433_ sky130_fd_sc_hd__mux2_1
X_18181_ net1192 _01709_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[20\] sky130_fd_sc_hd__dfxtp_1
X_15393_ _03098_ _03446_ _03448_ _03307_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17132_ CPU.registerFile\[19\]\[27\] CPU.registerFile\[18\]\[27\] _03745_ VGND VGND
+ VPWR VPWR _04832_ sky130_fd_sc_hd__mux2_1
X_14344_ _08418_ VGND VGND VPWR VPWR _08590_ sky130_fd_sc_hd__buf_4
XFILLER_0_123_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11556_ net1712 _07343_ _07390_ VGND VGND VPWR VPWR _07396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17063_ _08397_ _04762_ _04764_ _04410_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10507_ _06717_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__clkbuf_1
X_14275_ _08520_ VGND VGND VPWR VPWR _08521_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11487_ _07311_ VGND VGND VPWR VPWR _07354_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16014_ _06148_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__clkbuf_4
X_13525__916 clknet_1_1__leaf__08437_ VGND VGND VPWR VPWR net972 sky130_fd_sc_hd__inv_2
XFILLER_0_150_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13226_ clknet_leaf_20_clk VGND VGND VPWR VPWR _08339_ sky130_fd_sc_hd__buf_1
X_10438_ _06680_ VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ net1571 _08285_ VGND VGND VPWR VPWR _08288_ sky130_fd_sc_hd__nor2_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _06637_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__clkbuf_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ net1372 _07693_ _07699_ _07175_ VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ CPU.registerFile\[4\]\[1\] net1362 _08216_ VGND VGND VPWR VPWR _08250_ sky130_fd_sc_hd__mux2_1
X_17965_ net976 _01493_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12039_ _07653_ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__clkbuf_1
X_16916_ _04574_ _04617_ _04621_ _04584_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__o211a_1
X_17896_ clknet_leaf_25_clk _01424_ VGND VGND VPWR VPWR CPU.instr\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16847_ _04419_ _04551_ _04553_ _04383_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__a211o_1
X_16778_ CPU.registerFile\[24\]\[18\] _04319_ _04165_ _04486_ VGND VGND VPWR VPWR
+ _04487_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18517_ net338 _02041_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09250_ CPU.aluIn1\[9\] CPU.Bimm\[9\] VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__or2_1
X_18448_ net269 _01976_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09181_ _05532_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18379_ net200 _01907_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__08457_ _08457_ VGND VGND VPWR VPWR clknet_0__08457_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08965_ CPU.rs2\[12\] _05246_ _05250_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__o21ai_2
X_08896_ _05240_ _05241_ _05243_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09517_ _05856_ _05861_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09448_ _05793_ _05796_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__nand2_1
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09379_ _05555_ _05728_ _05730_ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_35_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11410_ net1730 _06440_ _07296_ VGND VGND VPWR VPWR _07303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12390_ _06655_ net2037 _07870_ VGND VGND VPWR VPWR _07879_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15876__621 clknet_1_1__leaf__03682_ VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__inv_2
X_11341_ _07266_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11272_ _07229_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__clkbuf_1
X_13011_ _08209_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__clkbuf_1
X_10223_ _05417_ _06541_ _06543_ VGND VGND VPWR VPWR _06544_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_101_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13974__131 clknet_1_0__leaf__08481_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__inv_2
X_13922__83 clknet_1_0__leaf__08477_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__inv_2
X_10154_ _05794_ _05444_ VGND VGND VPWR VPWR _06478_ sky130_fd_sc_hd__nand2_1
X_17750_ net835 _01316_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_14962_ _02831_ _02832_ CPU.registerFile\[1\]\[15\] VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__a21o_1
Xhold7 _07844_ VGND VGND VPWR VPWR net1304 sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ _06176_ net1376 _06403_ _06411_ VGND VGND VPWR VPWR _06412_ sky130_fd_sc_hd__a211o_2
X_16701_ _04170_ _04406_ _04411_ _04180_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17681_ _05708_ _05209_ _05210_ _07673_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__nand4_4
X_14893_ CPU.registerFile\[21\]\[14\] _02960_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__or2_1
X_16632_ CPU.registerFile\[6\]\[15\] CPU.registerFile\[7\]\[15\] _04022_ VGND VGND
+ VPWR VPWR _04344_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__08446_ clknet_0__08446_ VGND VGND VPWR VPWR clknet_1_0__leaf__08446_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13775_ clknet_1_0__leaf__08340_ VGND VGND VPWR VPWR _08462_ sky130_fd_sc_hd__buf_1
X_16563_ CPU.registerFile\[30\]\[13\] CPU.registerFile\[31\]\[13\] _04201_ VGND VGND
+ VPWR VPWR _04277_ sky130_fd_sc_hd__mux2_1
X_10987_ _07023_ _07030_ _07032_ _06853_ VGND VGND VPWR VPWR _07033_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18302_ net123 _01830_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_12726_ _08057_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__clkbuf_1
X_15514_ _08513_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__buf_2
XFILLER_0_29_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16494_ _04075_ _04204_ _04209_ _04042_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18233_ net1244 net17 VGND VGND VPWR VPWR mapped_spi_flash.div_counter\[2\] sky130_fd_sc_hd__dfxtp_1
X_15445_ _03156_ _03496_ _03498_ _03163_ VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__a211o_1
X_12657_ _06649_ net2007 _08015_ VGND VGND VPWR VPWR _08021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11608_ net1799 _07326_ _07416_ VGND VGND VPWR VPWR _07424_ sky130_fd_sc_hd__mux2_1
X_18164_ net1175 _01692_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[3\] sky130_fd_sc_hd__dfxtp_1
X_15376_ CPU.registerFile\[20\]\[26\] _03080_ _03431_ _03082_ VGND VGND VPWR VPWR
+ _03432_ sky130_fd_sc_hd__o211a_1
X_12588_ _07984_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14327_ _08557_ _08563_ _08572_ _08423_ VGND VGND VPWR VPWR _08573_ sky130_fd_sc_hd__o211a_1
X_17115_ CPU.registerFile\[2\]\[27\] CPU.registerFile\[3\]\[27\] _03759_ VGND VGND
+ VPWR VPWR _04815_ sky130_fd_sc_hd__mux2_1
X_11539_ net1857 _07326_ _07379_ VGND VGND VPWR VPWR _07387_ sky130_fd_sc_hd__mux2_1
X_18095_ net1106 _01623_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold407 CPU.registerFile\[31\]\[5\] VGND VGND VPWR VPWR net1704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 CPU.registerFile\[10\]\[29\] VGND VGND VPWR VPWR net1715 sky130_fd_sc_hd__dlygate4sd3_1
X_15777__563 clknet_1_1__leaf__03656_ VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__inv_2
X_17046_ _03765_ _04745_ _04747_ _04521_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__a211o_1
XFILLER_0_111_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold429 CPU.registerFile\[28\]\[7\] VGND VGND VPWR VPWR net1726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03684_ clknet_0__03684_ VGND VGND VPWR VPWR clknet_1_1__leaf__03684_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13209_ _05752_ _05773_ _05830_ VGND VGND VPWR VPWR _08323_ sky130_fd_sc_hd__or3_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13306__807 clknet_1_1__leaf__08362_ VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__inv_2
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ clknet_leaf_13_clk _02517_ VGND VGND VPWR VPWR CPU.aluIn1\[14\] sky130_fd_sc_hd__dfxtp_4
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 CPU.registerFile\[14\]\[19\] VGND VGND VPWR VPWR net2404 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ net959 _01476_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[18\] sky130_fd_sc_hd__dfxtp_1
Xhold1118 CPU.registerFile\[20\]\[10\] VGND VGND VPWR VPWR net2415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 CPU.registerFile\[29\]\[31\] VGND VGND VPWR VPWR net2426 sky130_fd_sc_hd__dlygate4sd3_1
X_17879_ clknet_leaf_18_clk _00029_ VGND VGND VPWR VPWR CPU.cycles\[22\] sky130_fd_sc_hd__dfxtp_1
X_13495__889 clknet_1_0__leaf__08434_ VGND VGND VPWR VPWR net945 sky130_fd_sc_hd__inv_2
X_17422__43 clknet_1_1__leaf__05015_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__inv_2
XFILLER_0_49_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13634__1014 clknet_1_1__leaf__08448_ VGND VGND VPWR VPWR net1070 sky130_fd_sc_hd__inv_2
X_13239__761 clknet_1_0__leaf__08342_ VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__inv_2
XFILLER_0_76_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09302_ CPU.aluIn1\[23\] _05545_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09233_ _05573_ _05583_ _05584_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09164_ _05514_ _05515_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__nor2_2
XFILLER_0_72_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09095_ _05430_ _05446_ _05300_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__a21o_1
Xhold930 CPU.registerFile\[18\]\[0\] VGND VGND VPWR VPWR net2227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 CPU.registerFile\[20\]\[7\] VGND VGND VPWR VPWR net2238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__08509_ _08509_ VGND VGND VPWR VPWR clknet_0__08509_ sky130_fd_sc_hd__clkbuf_16
Xhold952 CPU.registerFile\[29\]\[6\] VGND VGND VPWR VPWR net2249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 CPU.registerFile\[9\]\[22\] VGND VGND VPWR VPWR net2260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold974 CPU.registerFile\[14\]\[4\] VGND VGND VPWR VPWR net2271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 CPU.registerFile\[29\]\[30\] VGND VGND VPWR VPWR net2282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 CPU.registerFile\[26\]\[22\] VGND VGND VPWR VPWR net2293 sky130_fd_sc_hd__dlygate4sd3_1
X_09997_ _05972_ _05945_ VGND VGND VPWR VPWR _06327_ sky130_fd_sc_hd__and2b_1
X_08948_ _05298_ _05299_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__nor2_2
X_10910_ _06972_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__clkbuf_1
X_11890_ _07574_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10841_ CPU.aluReg\[17\] CPU.aluReg\[15\] _06906_ VGND VGND VPWR VPWR _06920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10772_ CPU.aluIn1\[31\] _06861_ _06863_ _06865_ VGND VGND VPWR VPWR _06866_ sky130_fd_sc_hd__o22a_1
XFILLER_0_137_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12511_ _07943_ VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15230_ _03078_ _03287_ _03289_ _03043_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__a211o_1
XFILLER_0_137_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12442_ net1718 _07353_ _07906_ VGND VGND VPWR VPWR _07907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15161_ CPU.registerFile\[13\]\[20\] CPU.registerFile\[12\]\[20\] _02935_ VGND VGND
+ VPWR VPWR _03223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12373_ _07847_ VGND VGND VPWR VPWR _07870_ sky130_fd_sc_hd__buf_4
XFILLER_0_22_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14041__191 clknet_1_1__leaf__08488_ VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__inv_2
X_17293__709 clknet_1_0__leaf__04979_ VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__inv_2
X_11324_ _07257_ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__clkbuf_1
X_15092_ _06339_ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__clkbuf_4
X_18920_ net694 _02440_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_11255_ _07220_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__clkbuf_1
X_10206_ _06524_ _06525_ _06526_ _06527_ _05541_ VGND VGND VPWR VPWR _06528_ sky130_fd_sc_hd__o41a_2
X_18851_ net625 _00004_ VGND VGND VPWR VPWR mapped_spi_flash.state\[0\] sky130_fd_sc_hd__dfxtp_1
X_11186_ _07176_ _07177_ VGND VGND VPWR VPWR _07178_ sky130_fd_sc_hd__nor2_1
X_17802_ net882 _01364_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_10137_ _06390_ _06391_ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__nand2_1
X_18782_ net571 _02306_ VGND VGND VPWR VPWR CPU.aluReg\[12\] sky130_fd_sc_hd__dfxtp_1
X_15994_ _03718_ _03719_ _03720_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__mux2_1
X_17733_ net818 _01299_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_10068_ _05693_ _06393_ VGND VGND VPWR VPWR _06395_ sky130_fd_sc_hd__nor2_2
X_14945_ _02798_ _02997_ _03002_ _03011_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__a31o_1
X_17664_ per_uart.uart0.rx_bitcount\[1\] _05195_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__or2_1
X_14876_ CPU.registerFile\[5\]\[13\] CPU.registerFile\[4\]\[13\] _08864_ VGND VGND
+ VPWR VPWR _02945_ sky130_fd_sc_hd__mux2_1
X_16615_ CPU.registerFile\[19\]\[14\] CPU.registerFile\[18\]\[14\] _04327_ VGND VGND
+ VPWR VPWR _04328_ sky130_fd_sc_hd__mux2_1
X_17595_ per_uart.uart0.tx_bitcount\[1\] per_uart.uart0.tx_bitcount\[0\] per_uart.uart0.tx_bitcount\[2\]
+ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16546_ CPU.registerFile\[10\]\[13\] CPU.registerFile\[11\]\[13\] _03931_ VGND VGND
+ VPWR VPWR _04260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12709_ _08048_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16477_ CPU.registerFile\[5\]\[11\] CPU.registerFile\[4\]\[11\] _04024_ VGND VGND
+ VPWR VPWR _04193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18216_ net1227 _01744_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15428_ CPU.registerFile\[8\]\[27\] _08545_ _03482_ _03268_ VGND VGND VPWR VPWR _03483_
+ sky130_fd_sc_hd__o211a_1
X_19196_ net106 net54 VGND VGND VPWR VPWR mapped_spi_ram.div_counter\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18147_ net1158 _01675_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_15359_ CPU.registerFile\[6\]\[25\] CPU.registerFile\[7\]\[25\] _08536_ VGND VGND
+ VPWR VPWR _03416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold204 _01321_ VGND VGND VPWR VPWR net1501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 mapped_spi_flash.cmd_addr\[9\] VGND VGND VPWR VPWR net1512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18078_ net1089 _01606_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[20\] sky130_fd_sc_hd__dfxtp_1
Xhold226 mapped_spi_ram.rcv_data\[24\] VGND VGND VPWR VPWR net1523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 mapped_spi_flash.cmd_addr\[6\] VGND VGND VPWR VPWR net1534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold248 mapped_spi_flash.cmd_addr\[2\] VGND VGND VPWR VPWR net1545 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ _05261_ _05311_ _05313_ _05315_ VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__o31a_1
Xhold259 mapped_spi_ram.rcv_data\[18\] VGND VGND VPWR VPWR net1556 sky130_fd_sc_hd__dlygate4sd3_1
X_17029_ _04723_ _04731_ _04542_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__o21a_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09851_ _05321_ _05324_ _05335_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__o21a_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _05929_ _05994_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__xnor2_1
X_13901__64 clknet_1_1__leaf__08475_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__inv_2
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503__896 clknet_1_0__leaf__08435_ VGND VGND VPWR VPWR net952 sky130_fd_sc_hd__inv_2
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_918 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09216_ CPU.aluIn1\[7\] CPU.Bimm\[7\] VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14099__243 clknet_1_0__leaf__08494_ VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__inv_2
X_09147_ _05387_ CPU.aluIn1\[24\] VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09078_ _05285_ _05284_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__or2b_1
XFILLER_0_20_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold760 CPU.registerFile\[17\]\[19\] VGND VGND VPWR VPWR net2057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 CPU.registerFile\[18\]\[27\] VGND VGND VPWR VPWR net2068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 CPU.registerFile\[18\]\[30\] VGND VGND VPWR VPWR net2079 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ _07023_ _07077_ _07078_ _06853_ VGND VGND VPWR VPWR _07079_ sky130_fd_sc_hd__o211a_1
X_15914__654 clknet_1_1__leaf__03687_ VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__inv_2
Xhold793 CPU.registerFile\[14\]\[18\] VGND VGND VPWR VPWR net2090 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12991_ net2218 _07345_ _08192_ VGND VGND VPWR VPWR _08199_ sky130_fd_sc_hd__mux2_1
X_11942_ _06603_ net2510 _07598_ VGND VGND VPWR VPWR _07602_ sky130_fd_sc_hd__mux2_1
X_14730_ _02751_ _02799_ _02801_ _02759_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _02733_ _02734_ CPU.registerFile\[9\]\[8\] VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__a21o_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _07565_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18595__52 VGND VGND VPWR VPWR _18595__52/HI net52 sky130_fd_sc_hd__conb_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16400_ _03943_ _04114_ _04116_ _04117_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_0__f__03687_ clknet_0__03687_ VGND VGND VPWR VPWR clknet_1_0__leaf__03687_
+ sky130_fd_sc_hd__clkbuf_16
X_10824_ CPU.aluReg\[21\] CPU.aluReg\[19\] _06906_ VGND VGND VPWR VPWR _06907_ sky130_fd_sc_hd__mux2_1
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17380_ _04996_ _05005_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__and2_1
X_14592_ _08425_ _08814_ _08831_ _08597_ VGND VGND VPWR VPWR _08832_ sky130_fd_sc_hd__a211o_1
X_13335__833 clknet_1_0__leaf__08365_ VGND VGND VPWR VPWR net889 sky130_fd_sc_hd__inv_2
X_17401__24 clknet_1_0__leaf__05013_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__inv_2
XFILLER_0_94_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16331_ _03758_ _04046_ _04050_ _03775_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15960__696 clknet_1_0__leaf__03691_ VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__inv_2
X_10755_ mapped_spi_flash.state\[2\] CPU.mem_rstrb _05860_ VGND VGND VPWR VPWR _06851_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_109_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16262_ _03981_ _03982_ _03720_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19050_ net792 _02570_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_13474_ _08428_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10686_ _05737_ _05738_ _05739_ VGND VGND VPWR VPWR _06814_ sky130_fd_sc_hd__and3b_2
X_15213_ _03272_ _03273_ _03025_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__mux2_1
X_17301__716 clknet_1_1__leaf__04980_ VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__inv_2
X_18001_ net1012 _01529_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12425_ net1935 _07337_ _07895_ VGND VGND VPWR VPWR _07898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16193_ _03749_ _03751_ CPU.registerFile\[25\]\[4\] VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15144_ _03156_ _03203_ _03205_ _03163_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__a211o_1
X_12356_ _07861_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11307_ _07248_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15075_ _06059_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__clkbuf_4
X_12287_ net1458 _07812_ _07818_ _07809_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18903_ net677 _02423_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_13633__1013 clknet_1_1__leaf__08448_ VGND VGND VPWR VPWR net1069 sky130_fd_sc_hd__inv_2
X_11238_ _07211_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18834_ net623 _02358_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_11169_ net1643 _07134_ VGND VGND VPWR VPWR _07168_ sky130_fd_sc_hd__or2_1
X_18765_ net554 _02289_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[27\] sky130_fd_sc_hd__dfxtp_1
X_15977_ _03696_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14928_ CPU.registerFile\[17\]\[15\] _08795_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__or2_1
X_18696_ net485 net1445 VGND VGND VPWR VPWR mapped_spi_flash.rcv_bitcount\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17647_ net2622 net2673 VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__nand2_1
X_14859_ _08525_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17578_ _05140_ VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14048__197 clknet_1_0__leaf__08489_ VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__inv_2
XFILLER_0_129_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16529_ _04080_ _04081_ CPU.registerFile\[25\]\[12\] VGND VGND VPWR VPWR _04244_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09001_ CPU.rs2\[18\] _05246_ _05250_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__o21a_1
X_19179_ clknet_leaf_0_clk _02699_ VGND VGND VPWR VPWR per_uart.rx_error sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09903_ _05888_ _06236_ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__or2_1
X_15636__437 clknet_1_0__leaf__03641_ VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__inv_2
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09834_ _06170_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__clkbuf_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _05764_ _06086_ _06102_ _06104_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__a211o_4
X_09696_ _05856_ _06037_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__nand2_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10540_ _06734_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10471_ _06697_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12210_ mapped_spi_ram.snd_bitcount\[2\] mapped_spi_ram.snd_bitcount\[1\] mapped_spi_ram.snd_bitcount\[0\]
+ VGND VGND VPWR VPWR _07770_ sky130_fd_sc_hd__or3_1
X_13190_ _08305_ net1550 VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12141_ mapped_spi_ram.cmd_addr\[17\] _07051_ _07704_ VGND VGND VPWR VPWR _07722_
+ sky130_fd_sc_hd__mux2_1
X_12072_ CPU.mem_rstrb _05858_ VGND VGND VPWR VPWR _07671_ sky130_fd_sc_hd__and2_2
Xhold590 CPU.registerFile\[22\]\[12\] VGND VGND VPWR VPWR net1887 sky130_fd_sc_hd__dlygate4sd3_1
X_11023_ _05599_ _07056_ VGND VGND VPWR VPWR _07064_ sky130_fd_sc_hd__xnor2_1
X_16880_ _04545_ _04564_ _04586_ _04500_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__a211o_1
X_18550_ net371 _02074_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_12974_ net2315 _07328_ _08181_ VGND VGND VPWR VPWR _08190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1290 CPU.registerFile\[24\]\[26\] VGND VGND VPWR VPWR net2587 sky130_fd_sc_hd__dlygate4sd3_1
X_17501_ _08335_ _06212_ _05073_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__o21ai_1
X_14713_ CPU.registerFile\[6\]\[9\] CPU.registerFile\[7\]\[9\] _08740_ VGND VGND VPWR
+ VPWR _02786_ sky130_fd_sc_hd__mux2_1
X_18481_ net302 _02005_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_11925_ _07592_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__clkbuf_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _08334_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__buf_2
XFILLER_0_129_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ net2594 _07368_ _07548_ VGND VGND VPWR VPWR _07556_ sky130_fd_sc_hd__mux2_1
X_14644_ _08837_ _08879_ _02717_ _08802_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__a211o_1
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10807_ CPU.aluReg\[25\] CPU.aluReg\[23\] _06872_ VGND VGND VPWR VPWR _06894_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14575_ CPU.registerFile\[15\]\[6\] CPU.registerFile\[14\]\[6\] _08771_ VGND VGND
+ VPWR VPWR _08815_ sky130_fd_sc_hd__mux2_1
X_17363_ per_uart.uart0.rxd_reg\[2\] _04992_ _04993_ per_uart.uart0.rxd_reg\[1\] VGND
+ VGND VPWR VPWR _04994_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11787_ _07519_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__clkbuf_1
X_19102_ net85 _02622_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16314_ CPU.registerFile\[30\]\[7\] CPU.registerFile\[31\]\[7\] _03796_ VGND VGND
+ VPWR VPWR _04034_ sky130_fd_sc_hd__mux2_1
X_10738_ _06842_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19033_ net775 _02553_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13457_ CPU.Iimm\[1\] _08415_ _08416_ VGND VGND VPWR VPWR _08417_ sky130_fd_sc_hd__mux2_1
X_16245_ _03963_ _03964_ _03966_ _06142_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__a211o_1
X_10669_ _06804_ VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12408_ net1711 _07320_ _07884_ VGND VGND VPWR VPWR _07889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__08490_ _08490_ VGND VGND VPWR VPWR clknet_0__08490_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_112_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16176_ CPU.registerFile\[12\]\[4\] _03707_ _03708_ _03898_ VGND VGND VPWR VPWR _03899_
+ sky130_fd_sc_hd__o211a_1
X_13388_ _05538_ _05539_ _08371_ _05422_ VGND VGND VPWR VPWR _08372_ sky130_fd_sc_hd__and4b_1
XFILLER_0_140_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15127_ CPU.registerFile\[6\]\[19\] CPU.registerFile\[7\]\[19\] _02982_ VGND VGND
+ VPWR VPWR _03190_ sky130_fd_sc_hd__mux2_1
X_12339_ _07852_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__clkbuf_1
X_15058_ CPU.registerFile\[20\]\[18\] _03080_ _03121_ _03082_ VGND VGND VPWR VPWR
+ _03122_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14009_ clknet_1_0__leaf__08484_ VGND VGND VPWR VPWR _08486_ sky130_fd_sc_hd__buf_1
X_18817_ net606 _02341_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_09550_ CPU.PC\[22\] CPU.PC\[21\] _05893_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__and3_1
X_18748_ net537 _02272_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09481_ _05555_ _05827_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__or2_1
X_18679_ net468 _02203_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13615__997 clknet_1_0__leaf__08446_ VGND VGND VPWR VPWR net1053 sky130_fd_sc_hd__inv_2
XFILLER_0_59_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09817_ _05912_ _06153_ VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__nor2_1
X_17330__742 clknet_1_0__leaf__04983_ VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__inv_2
X_09748_ _05892_ _06087_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__or2_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _05377_ _05747_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__nor2_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _07478_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__clkbuf_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _08038_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18565__22 VGND VGND VPWR VPWR _18565__22/HI net22 sky130_fd_sc_hd__conb_1
XFILLER_0_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _07441_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__clkbuf_1
X_13632__1012 clknet_1_1__leaf__08448_ VGND VGND VPWR VPWR net1068 sky130_fd_sc_hd__inv_2
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14360_ CPU.registerFile\[20\]\[1\] _08527_ _08604_ _08530_ VGND VGND VPWR VPWR _08605_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11572_ _07404_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13311_ clknet_1_1__leaf__08341_ VGND VGND VPWR VPWR _08363_ sky130_fd_sc_hd__buf_1
X_10523_ net2474 _06316_ _06724_ VGND VGND VPWR VPWR _06726_ sky130_fd_sc_hd__mux2_1
X_14291_ CPU.registerFile\[30\]\[0\] CPU.registerFile\[31\]\[0\] _08536_ VGND VGND
+ VPWR VPWR _08537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16030_ _03712_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__buf_4
XFILLER_0_122_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10454_ _06641_ net2288 _06687_ VGND VGND VPWR VPWR _06689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13173_ net1614 _08295_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__xor2_1
X_10385_ _06648_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__clkbuf_1
X_12124_ _07696_ _07709_ VGND VGND VPWR VPWR _07710_ sky130_fd_sc_hd__or2_1
X_17981_ net992 _01509_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_15771__558 clknet_1_1__leaf__03655_ VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__inv_2
X_16932_ _06172_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__clkbuf_4
X_12055_ CPU.registerFile\[24\]\[7\] _07362_ _07657_ VGND VGND VPWR VPWR _07662_ sky130_fd_sc_hd__mux2_1
X_11006_ _05608_ _07026_ VGND VGND VPWR VPWR _07049_ sky130_fd_sc_hd__xnor2_1
X_16863_ _04484_ _04485_ CPU.registerFile\[25\]\[20\] VGND VGND VPWR VPWR _04570_
+ sky130_fd_sc_hd__a21o_1
X_18602_ net423 _02126_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_15814_ _08358_ _03675_ _03660_ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__a21oi_1
X_16794_ _08403_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18533_ net354 _02057_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12957_ _08180_ VGND VGND VPWR VPWR _08181_ sky130_fd_sc_hd__buf_4
X_13808__1171 clknet_1_0__leaf__08465_ VGND VGND VPWR VPWR net1227 sky130_fd_sc_hd__inv_2
X_18464_ net285 _00008_ VGND VGND VPWR VPWR mapped_spi_ram.state\[0\] sky130_fd_sc_hd__dfxtp_1
X_11908_ _07583_ VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__clkbuf_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _06595_ _07199_ VGND VGND VPWR VPWR _08144_ sky130_fd_sc_hd__nand2_4
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14627_ _08863_ _08865_ _08783_ VGND VGND VPWR VPWR _08866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11839_ net2193 _07351_ _07537_ VGND VGND VPWR VPWR _07547_ sky130_fd_sc_hd__mux2_1
X_18395_ net216 _01923_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14558_ _08415_ _08793_ _08797_ _08420_ VGND VGND VPWR VPWR _08798_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__08511_ clknet_0__08511_ VGND VGND VPWR VPWR clknet_1_1__leaf__08511_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13509_ clknet_1_0__leaf__08366_ VGND VGND VPWR VPWR _08436_ sky130_fd_sc_hd__buf_1
XFILLER_0_153_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17277_ _03749_ _03751_ CPU.registerFile\[17\]\[31\] VGND VGND VPWR VPWR _04973_
+ sky130_fd_sc_hd__a21o_1
X_14489_ _08515_ _08716_ _08721_ _08730_ VGND VGND VPWR VPWR _08731_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19016_ net758 _02536_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[1\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__08442_ clknet_0__08442_ VGND VGND VPWR VPWR clknet_1_1__leaf__08442_
+ sky130_fd_sc_hd__clkbuf_16
X_16228_ CPU.registerFile\[30\]\[5\] CPU.registerFile\[31\]\[5\] _03796_ VGND VGND
+ VPWR VPWR _03950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08473_ _08473_ VGND VGND VPWR VPWR clknet_0__08473_ sky130_fd_sc_hd__clkbuf_16
X_16159_ _03736_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__buf_4
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08981_ _05331_ _05332_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__or2_2
XFILLER_0_139_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09602_ CPU.Bimm\[8\] _05914_ CPU.PC\[8\] VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__a21o_1
X_09533_ _05856_ _05876_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15748__538 clknet_1_1__leaf__03652_ VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__inv_2
X_09464_ _05396_ _05811_ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09395_ CPU.Jimm\[12\] _05527_ VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10170_ mapped_spi_flash.rcv_data\[26\] _05859_ _05719_ per_uart.rx_data\[2\] _06492_
+ VGND VGND VPWR VPWR _06493_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__08462_ clknet_0__08462_ VGND VGND VPWR VPWR clknet_1_0__leaf__08462_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12811_ _06859_ VGND VGND VPWR VPWR _08103_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ _06013_ _03577_ _03581_ _08422_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__o211a_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _08066_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15461_ _03513_ _03514_ _08541_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__mux2_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _06593_ net2636 _08029_ VGND VGND VPWR VPWR _08030_ sky130_fd_sc_hd__mux2_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _03714_ _04893_ _04897_ _08403_ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14412_ CPU.registerFile\[13\]\[2\] CPU.registerFile\[12\]\[2\] _08560_ VGND VGND
+ VPWR VPWR _08656_ sky130_fd_sc_hd__mux2_1
X_11624_ _07432_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__clkbuf_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18180_ net1191 net1557 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[19\] sky130_fd_sc_hd__dfxtp_1
X_15392_ CPU.registerFile\[8\]\[26\] _08545_ _03447_ _03268_ VGND VGND VPWR VPWR _03448_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17131_ _04829_ _04830_ _03742_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__mux2_1
X_11555_ _07395_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__clkbuf_1
X_14343_ CPU.registerFile\[0\]\[0\] _08584_ _08587_ _08588_ VGND VGND VPWR VPWR _08589_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10506_ net2214 _06124_ _06713_ VGND VGND VPWR VPWR _06717_ sky130_fd_sc_hd__mux2_1
X_14274_ _06418_ VGND VGND VPWR VPWR _08520_ sky130_fd_sc_hd__clkbuf_8
X_17062_ CPU.registerFile\[16\]\[25\] _04656_ _04494_ _04763_ VGND VGND VPWR VPWR
+ _04764_ sky130_fd_sc_hd__o211a_1
X_11486_ _06291_ VGND VGND VPWR VPWR _07353_ sky130_fd_sc_hd__buf_4
X_16013_ CPU.registerFile\[28\]\[0\] CPU.registerFile\[29\]\[0\] _03739_ VGND VGND
+ VPWR VPWR _03740_ sky130_fd_sc_hd__mux2_1
X_13225_ net2659 _08332_ _08338_ _07822_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__o211a_1
X_10437_ _06624_ net2090 _06676_ VGND VGND VPWR VPWR _06680_ sky130_fd_sc_hd__mux2_1
X_15853__600 clknet_1_1__leaf__03680_ VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__inv_2
XFILLER_0_0_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13156_ CPU.cycles\[15\] _08285_ VGND VGND VPWR VPWR _08287_ sky130_fd_sc_hd__and2_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _06636_ net1957 _06618_ VGND VGND VPWR VPWR _06637_ sky130_fd_sc_hd__mux2_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ net1371 _07694_ _07696_ VGND VGND VPWR VPWR _07699_ sky130_fd_sc_hd__a21o_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17964_ net975 _01492_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_13087_ net1423 VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__clkbuf_1
X_10299_ net1779 _06508_ _06580_ VGND VGND VPWR VPWR _06590_ sky130_fd_sc_hd__mux2_1
X_12038_ CPU.registerFile\[24\]\[15\] _07345_ _07646_ VGND VGND VPWR VPWR _07653_
+ sky130_fd_sc_hd__mux2_1
X_16915_ _04367_ _04618_ _04620_ _04410_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__a211o_1
X_13951__110 clknet_1_0__leaf__08479_ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__inv_2
X_17895_ clknet_leaf_22_clk _01423_ VGND VGND VPWR VPWR CPU.instr\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16846_ CPU.registerFile\[12\]\[20\] _04421_ _04422_ _04552_ VGND VGND VPWR VPWR
+ _04553_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16777_ _04484_ _04485_ CPU.registerFile\[25\]\[18\] VGND VGND VPWR VPWR _04486_
+ sky130_fd_sc_hd__a21o_1
X_18516_ net337 _02040_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15589__394 clknet_1_0__leaf__08511_ VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__inv_2
XFILLER_0_75_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18447_ net268 _01975_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09180_ _05531_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18378_ net199 _01906_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17329_ clknet_1_1__leaf__03686_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__buf_1
XFILLER_0_126_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14093__238 clknet_1_1__leaf__08493_ VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__inv_2
Xclkbuf_0__08456_ _08456_ VGND VGND VPWR VPWR clknet_0__08456_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08964_ CPU.rs2\[12\] _05246_ _05250_ CPU.aluIn1\[12\] VGND VGND VPWR VPWR _05316_
+ sky130_fd_sc_hd__o211a_1
X_08895_ _05246_ VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09516_ mapped_spi_ram.rcv_data\[0\] _05858_ _05860_ net1379 VGND VGND VPWR VPWR
+ _05861_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_67_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09447_ _05410_ _05506_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__xor2_1
XFILLER_0_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09378_ _05422_ _05538_ _05729_ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__nor3_1
XFILLER_0_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11340_ net2652 _06413_ _07260_ VGND VGND VPWR VPWR _07266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11271_ _06649_ net2403 _07223_ VGND VGND VPWR VPWR _07229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13907__70 clknet_1_0__leaf__08475_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__inv_2
XFILLER_0_132_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13010_ net2349 _07364_ _08203_ VGND VGND VPWR VPWR _08209_ sky130_fd_sc_hd__mux2_1
X_10222_ _05413_ _05506_ _06542_ _05419_ VGND VGND VPWR VPWR _06543_ sky130_fd_sc_hd__a31o_1
X_13807__1170 clknet_1_0__leaf__08465_ VGND VGND VPWR VPWR net1226 sky130_fd_sc_hd__inv_2
XFILLER_0_101_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10153_ _05283_ _05443_ VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__xnor2_1
X_14961_ CPU.registerFile\[2\]\[15\] CPU.registerFile\[3\]\[15\] _02871_ VGND VGND
+ VPWR VPWR _03028_ sky130_fd_sc_hd__mux2_1
X_10084_ _06408_ _06410_ _05745_ VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__o21a_1
Xhold8 _01684_ VGND VGND VPWR VPWR net1305 sky130_fd_sc_hd__dlygate4sd3_1
X_16700_ _04367_ _04407_ _04409_ _04410_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__a211o_1
X_17680_ _05715_ _05704_ VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__nor2_1
X_14892_ _06062_ VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__buf_2
X_16631_ _04015_ _04340_ _04342_ _03979_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_0__f__08445_ clknet_0__08445_ VGND VGND VPWR VPWR clknet_1_0__leaf__08445_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16562_ _04098_ _04263_ _04267_ _04275_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__a31o_2
X_10986_ CPU.PC\[15\] _07031_ VGND VGND VPWR VPWR _07032_ sky130_fd_sc_hd__or2_1
X_18301_ net122 _01829_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_15513_ net1589 _03201_ _03565_ _03390_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__o211a_1
X_12725_ _06649_ CPU.registerFile\[25\]\[6\] _08051_ VGND VGND VPWR VPWR _08057_ sky130_fd_sc_hd__mux2_1
X_16493_ _04037_ _04205_ _04207_ _04208_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__a211o_1
XFILLER_0_139_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18232_ net1243 _01760_ VGND VGND VPWR VPWR mapped_spi_flash.div_counter\[1\] sky130_fd_sc_hd__dfxtp_1
X_15444_ CPU.registerFile\[16\]\[28\] _03159_ _03497_ _03161_ VGND VGND VPWR VPWR
+ _03498_ sky130_fd_sc_hd__o211a_1
X_12656_ _08020_ VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11607_ _07423_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__clkbuf_1
X_18163_ net1174 net1470 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12587_ net2286 _07362_ _07979_ VGND VGND VPWR VPWR _07984_ sky130_fd_sc_hd__mux2_1
X_15375_ CPU.registerFile\[21\]\[26\] _02752_ VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17114_ _04812_ _04813_ _04557_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__mux2_1
X_14326_ _08520_ _08565_ _08571_ _08419_ VGND VGND VPWR VPWR _08572_ sky130_fd_sc_hd__a211o_1
X_18094_ net1105 _01622_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_11538_ _07386_ VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold408 _08174_ VGND VGND VPWR VPWR net1705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold419 CPU.registerFile\[6\]\[11\] VGND VGND VPWR VPWR net1716 sky130_fd_sc_hd__dlygate4sd3_1
X_17045_ CPU.registerFile\[0\]\[25\] _04637_ _04472_ _04746_ VGND VGND VPWR VPWR _04747_
+ sky130_fd_sc_hd__o211a_1
X_11469_ net2001 _07341_ _07333_ VGND VGND VPWR VPWR _07342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03683_ clknet_0__03683_ VGND VGND VPWR VPWR clknet_1_1__leaf__03683_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13208_ _05796_ _05845_ _05901_ _08321_ VGND VGND VPWR VPWR _08322_ sky130_fd_sc_hd__or4_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13139_ CPU.cycles\[7\] CPU.cycles\[8\] _08275_ VGND VGND VPWR VPWR _08277_ sky130_fd_sc_hd__and3_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ clknet_leaf_14_clk _02516_ VGND VGND VPWR VPWR CPU.aluIn1\[13\] sky130_fd_sc_hd__dfxtp_4
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1108 CPU.registerFile\[12\]\[1\] VGND VGND VPWR VPWR net2405 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17947_ net958 _01475_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[17\] sky130_fd_sc_hd__dfxtp_1
Xhold1119 CPU.registerFile\[31\]\[23\] VGND VGND VPWR VPWR net2416 sky130_fd_sc_hd__dlygate4sd3_1
X_17878_ clknet_leaf_17_clk _00028_ VGND VGND VPWR VPWR CPU.cycles\[21\] sky130_fd_sc_hd__dfxtp_1
X_17407__30 clknet_1_1__leaf__05013_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__inv_2
XFILLER_0_45_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16829_ CPU.registerFile\[19\]\[19\] CPU.registerFile\[18\]\[19\] _04327_ VGND VGND
+ VPWR VPWR _04537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09301_ _05645_ _05648_ _05646_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09232_ CPU.aluIn1\[3\] _05572_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09163_ CPU.Jimm\[13\] CPU.Jimm\[12\] VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__or2_4
XFILLER_0_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09094_ _05431_ _05445_ _05286_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__a21o_1
X_14101__245 clknet_1_0__leaf__08494_ VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__inv_2
X_13508__901 clknet_1_1__leaf__08435_ VGND VGND VPWR VPWR net957 sky130_fd_sc_hd__inv_2
XFILLER_0_102_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold920 CPU.registerFile\[21\]\[0\] VGND VGND VPWR VPWR net2217 sky130_fd_sc_hd__dlygate4sd3_1
X_13958__116 clknet_1_0__leaf__08480_ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__inv_2
Xhold931 CPU.registerFile\[11\]\[12\] VGND VGND VPWR VPWR net2228 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__08508_ _08508_ VGND VGND VPWR VPWR clknet_0__08508_ sky130_fd_sc_hd__clkbuf_16
Xhold942 CPU.registerFile\[17\]\[17\] VGND VGND VPWR VPWR net2239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 CPU.registerFile\[14\]\[22\] VGND VGND VPWR VPWR net2250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 CPU.registerFile\[8\]\[14\] VGND VGND VPWR VPWR net2261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 CPU.registerFile\[17\]\[8\] VGND VGND VPWR VPWR net2272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 CPU.registerFile\[16\]\[22\] VGND VGND VPWR VPWR net2283 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__08439_ _08439_ VGND VGND VPWR VPWR clknet_0__08439_ sky130_fd_sc_hd__clkbuf_16
Xhold997 CPU.registerFile\[6\]\[28\] VGND VGND VPWR VPWR net2294 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__08339_ clknet_0__08339_ VGND VGND VPWR VPWR clknet_1_1__leaf__08339_
+ sky130_fd_sc_hd__clkbuf_16
X_09996_ _05265_ _05769_ _05770_ net1331 _06325_ VGND VGND VPWR VPWR _06326_ sky130_fd_sc_hd__a221o_2
XFILLER_0_86_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08947_ CPU.aluIn1\[6\] _05297_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10840_ _06919_ VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__clkbuf_1
X_10771_ CPU.aluReg\[30\] _05799_ _05770_ _06864_ VGND VGND VPWR VPWR _06865_ sky130_fd_sc_hd__a31o_1
XFILLER_0_109_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12510_ net1782 _07353_ _07942_ VGND VGND VPWR VPWR _07943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12441_ _07883_ VGND VGND VPWR VPWR _07906_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12372_ _07869_ VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__clkbuf_1
X_15160_ CPU.registerFile\[15\]\[20\] CPU.registerFile\[14\]\[20\] _03013_ VGND VGND
+ VPWR VPWR _03222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11323_ net2545 _06224_ _07249_ VGND VGND VPWR VPWR _07257_ sky130_fd_sc_hd__mux2_1
X_15091_ net1650 _02797_ _03154_ _02993_ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14076__222 clknet_1_1__leaf__08492_ VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__inv_2
X_14042_ clknet_1_0__leaf__08484_ VGND VGND VPWR VPWR _08489_ sky130_fd_sc_hd__buf_1
X_11254_ _06632_ net1920 _07212_ VGND VGND VPWR VPWR _07220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10205_ _05280_ _05533_ _05536_ net1361 VGND VGND VPWR VPWR _06527_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18850_ clknet_leaf_6_clk _02374_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11185_ mapped_spi_flash.div_counter\[0\] mapped_spi_flash.div_counter\[1\] VGND
+ VGND VPWR VPWR _07177_ sky130_fd_sc_hd__xnor2_1
X_17801_ net881 _01363_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_10136_ net1390 _05860_ _05719_ per_uart.rx_data\[4\] _06460_ VGND VGND VPWR VPWR
+ _06461_ sky130_fd_sc_hd__a221o_1
X_18781_ net570 _02305_ VGND VGND VPWR VPWR CPU.aluReg\[11\] sky130_fd_sc_hd__dfxtp_1
X_15993_ _06534_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__clkbuf_4
X_17732_ net817 _01298_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_10067_ _05691_ _06205_ VGND VGND VPWR VPWR _06394_ sky130_fd_sc_hd__or2_1
X_14944_ _02964_ _03005_ _03010_ _08851_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__o211a_1
X_17663_ _05197_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__clkbuf_1
X_14875_ CPU.registerFile\[6\]\[13\] CPU.registerFile\[7\]\[13\] _08740_ VGND VGND
+ VPWR VPWR _02944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16614_ _03744_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__buf_4
X_17594_ _05151_ _05152_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16545_ CPU.aluIn1\[12\] _04054_ _04258_ _04259_ VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10969_ _07008_ _07017_ VGND VGND VPWR VPWR _07018_ sky130_fd_sc_hd__or2_1
X_12708_ _06632_ net2570 _08040_ VGND VGND VPWR VPWR _08048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16476_ CPU.registerFile\[6\]\[11\] CPU.registerFile\[7\]\[11\] _04022_ VGND VGND
+ VPWR VPWR _04192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18215_ net1226 _01743_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15427_ _03138_ _03139_ CPU.registerFile\[9\]\[27\] VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__a21o_1
X_13312__812 clknet_1_0__leaf__08363_ VGND VGND VPWR VPWR net868 sky130_fd_sc_hd__inv_2
X_19195_ net105 net53 VGND VGND VPWR VPWR mapped_spi_ram.div_counter\[2\] sky130_fd_sc_hd__dfxtp_1
X_12639_ _08011_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18146_ net1157 _01674_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15358_ _03133_ _03410_ _03414_ _03188_ VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold205 CPU.cycles\[31\] VGND VGND VPWR VPWR net1502 sky130_fd_sc_hd__dlygate4sd3_1
X_14309_ _08535_ _08542_ _08553_ _08554_ VGND VGND VPWR VPWR _08555_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18077_ net1088 _01605_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15289_ CPU.registerFile\[2\]\[23\] CPU.registerFile\[3\]\[23\] _03275_ VGND VGND
+ VPWR VPWR _03348_ sky130_fd_sc_hd__mux2_1
Xhold216 mapped_spi_flash.cmd_addr\[4\] VGND VGND VPWR VPWR net1513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 mapped_spi_ram.rcv_data\[20\] VGND VGND VPWR VPWR net1524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 mapped_spi_ram.rcv_data\[23\] VGND VGND VPWR VPWR net1535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17028_ _04574_ _04726_ _04730_ _04584_ VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__o211a_1
Xhold249 mapped_spi_flash.cmd_addr\[21\] VGND VGND VPWR VPWR net1546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09850_ _05328_ _05470_ _06184_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__and3_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ CPU.Jimm\[18\] _05550_ _05790_ CPU.cycles\[18\] _06119_ VGND VGND VPWR VPWR
+ _06120_ sky130_fd_sc_hd__a221o_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ net753 _02499_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15831__580 clknet_1_1__leaf__03678_ VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__inv_2
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09215_ CPU.aluIn1\[7\] CPU.Bimm\[7\] VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14025__176 clknet_1_0__leaf__08487_ VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__inv_2
XFILLER_0_8_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09146_ _05386_ _05391_ _05400_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__and3_1
X_13584__969 clknet_1_1__leaf__08443_ VGND VGND VPWR VPWR net1025 sky130_fd_sc_hd__inv_2
XFILLER_0_121_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09077_ _05297_ CPU.aluIn1\[6\] VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__or2b_1
XFILLER_0_130_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold750 CPU.registerFile\[7\]\[19\] VGND VGND VPWR VPWR net2047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 CPU.registerFile\[12\]\[21\] VGND VGND VPWR VPWR net2058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 CPU.registerFile\[11\]\[15\] VGND VGND VPWR VPWR net2069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 CPU.registerFile\[2\]\[13\] VGND VGND VPWR VPWR net2080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 CPU.registerFile\[15\]\[8\] VGND VGND VPWR VPWR net2091 sky130_fd_sc_hd__dlygate4sd3_1
X_09979_ _05912_ _06306_ _06309_ VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__o21ai_1
X_15613__416 clknet_1_0__leaf__03639_ VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__inv_2
X_12990_ _08198_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11941_ _07601_ VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__clkbuf_1
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _06059_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__clkbuf_4
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _06601_ net1743 _07562_ VGND VGND VPWR VPWR _07565_ sky130_fd_sc_hd__mux2_1
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03686_ clknet_0__03686_ VGND VGND VPWR VPWR clknet_1_0__leaf__03686_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10823_ _06871_ VGND VGND VPWR VPWR _06906_ sky130_fd_sc_hd__clkbuf_4
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14591_ _08822_ _08830_ _08594_ VGND VGND VPWR VPWR _08831_ sky130_fd_sc_hd__o21a_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16330_ _03963_ _04047_ _04049_ _04006_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__a211o_1
X_13542_ clknet_1_0__leaf__08366_ VGND VGND VPWR VPWR _08439_ sky130_fd_sc_hd__buf_1
X_10754_ _06850_ VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16261_ CPU.registerFile\[5\]\[6\] CPU.registerFile\[4\]\[6\] _03704_ VGND VGND VPWR
+ VPWR _03982_ sky130_fd_sc_hd__mux2_1
X_13695__1069 clknet_1_1__leaf__08454_ VGND VGND VPWR VPWR net1125 sky130_fd_sc_hd__inv_2
X_13473_ CPU.Bimm\[6\] _05827_ _08416_ VGND VGND VPWR VPWR _08428_ sky130_fd_sc_hd__mux2_1
X_10685_ _06812_ VGND VGND VPWR VPWR _06813_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_125_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18000_ net1011 _01528_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_15212_ CPU.registerFile\[5\]\[21\] CPU.registerFile\[4\]\[21\] _03105_ VGND VGND
+ VPWR VPWR _03273_ sky130_fd_sc_hd__mux2_1
X_12424_ _07897_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__clkbuf_1
X_16192_ _03847_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15143_ CPU.registerFile\[16\]\[20\] _03159_ _03204_ _03161_ VGND VGND VPWR VPWR
+ _03205_ sky130_fd_sc_hd__o211a_1
X_12355_ _06620_ net1765 _07859_ VGND VGND VPWR VPWR _07861_ sky130_fd_sc_hd__mux2_1
X_11306_ net1979 _06032_ _07238_ VGND VGND VPWR VPWR _07248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15074_ _06058_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__clkbuf_4
X_12286_ net1454 _07813_ VGND VGND VPWR VPWR _07818_ sky130_fd_sc_hd__or2_1
X_11237_ _06615_ net2064 _07201_ VGND VGND VPWR VPWR _07211_ sky130_fd_sc_hd__mux2_1
X_18902_ net676 _02422_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11168_ net1346 _07160_ _07167_ _07164_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__o211a_1
X_18833_ net622 _02357_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_15889__632 clknet_1_1__leaf__03684_ VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__inv_2
X_10119_ _05290_ _06429_ VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__xor2_1
X_18764_ net553 _02288_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[26\] sky130_fd_sc_hd__dfxtp_1
X_15976_ _03702_ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__clkbuf_4
X_11099_ _07009_ _07114_ VGND VGND VPWR VPWR _07124_ sky130_fd_sc_hd__nor2_1
X_17715_ _05234_ VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__clkbuf_1
X_14927_ CPU.registerFile\[19\]\[15\] CPU.registerFile\[18\]\[15\] _02753_ VGND VGND
+ VPWR VPWR _02994_ sky130_fd_sc_hd__mux2_1
X_14130__271 clknet_1_0__leaf__08497_ VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__inv_2
X_18695_ net484 _02219_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_bitcount\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17646_ _04986_ per_uart.uart0.uart_rxd2 _03659_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__a21oi_4
X_14858_ CPU.registerFile\[27\]\[13\] CPU.registerFile\[26\]\[13\] _02768_ VGND VGND
+ VPWR VPWR _02927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13987__142 clknet_1_0__leaf__08483_ VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__inv_2
X_13809_ clknet_1_0__leaf__08462_ VGND VGND VPWR VPWR _08466_ sky130_fd_sc_hd__buf_1
X_17577_ _04996_ _05139_ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__and2_1
X_14789_ CPU.registerFile\[13\]\[11\] CPU.registerFile\[12\]\[11\] _08693_ VGND VGND
+ VPWR VPWR _02860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16528_ CPU.registerFile\[27\]\[12\] CPU.registerFile\[26\]\[12\] _04242_ VGND VGND
+ VPWR VPWR _04243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16459_ _03750_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09000_ _05351_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19178_ clknet_leaf_6_clk _02698_ VGND VGND VPWR VPWR per_uart.uart0.rx_bitcount\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18129_ net1140 _01657_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09902_ CPU.PC\[12\] _05887_ CPU.PC\[13\] VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03649_ clknet_0__03649_ VGND VGND VPWR VPWR clknet_1_1__leaf__03649_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_158_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09833_ net2220 _06169_ _06055_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__mux2_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13282__785 clknet_1_1__leaf__08345_ VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__inv_2
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14213__346 clknet_1_0__leaf__08505_ VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__inv_2
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _05912_ _06103_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__nor2_1
X_09695_ _06036_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14107__251 clknet_1_1__leaf__08494_ VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__inv_2
XFILLER_0_36_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10470_ _06657_ net2442 _06687_ VGND VGND VPWR VPWR _06697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09129_ _05477_ _05479_ _05480_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12140_ net1426 _07714_ _07721_ _07713_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__o211a_1
X_15838__586 clknet_1_0__leaf__03679_ VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__inv_2
XFILLER_0_103_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12071_ net1307 VGND VGND VPWR VPWR _07670_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold580 CPU.registerFile\[19\]\[19\] VGND VGND VPWR VPWR net1877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 CPU.registerFile\[13\]\[6\] VGND VGND VPWR VPWR net1888 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ net1497 _07054_ _07063_ _07014_ VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__o211a_1
X_14188__323 clknet_1_1__leaf__08503_ VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__inv_2
X_12973_ _08189_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__clkbuf_1
X_13892__56 clknet_1_1__leaf__08474_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__inv_2
Xhold1280 CPU.registerFile\[25\]\[16\] VGND VGND VPWR VPWR net2577 sky130_fd_sc_hd__dlygate4sd3_1
X_17500_ _05076_ _05077_ _05020_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__a21oi_1
Xhold1291 CPU.registerFile\[9\]\[7\] VGND VGND VPWR VPWR net2588 sky130_fd_sc_hd__dlygate4sd3_1
X_14712_ _02728_ _02778_ _02783_ _02784_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__o211a_1
X_18480_ net301 _02004_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_11924_ _06653_ net2188 _07584_ VGND VGND VPWR VPWR _07592_ sky130_fd_sc_hd__mux2_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _05018_ _05019_ _05020_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__a21oi_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ CPU.registerFile\[20\]\[8\] _08839_ _08880_ _08841_ VGND VGND VPWR VPWR _02717_
+ sky130_fd_sc_hd__o211a_1
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _07555_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__clkbuf_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10806_ _06893_ VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__clkbuf_1
X_17362_ per_uart.uart0.rx_ack _04992_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__nor2_4
X_14574_ _08515_ _08798_ _08803_ _08813_ VGND VGND VPWR VPWR _08814_ sky130_fd_sc_hd__a31o_1
X_11786_ _06651_ net1992 _07512_ VGND VGND VPWR VPWR _07519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19101_ net84 _02621_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16313_ _08404_ _04014_ _04021_ _04032_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__a31o_2
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10737_ net1955 _06361_ _06838_ VGND VGND VPWR VPWR _06842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19032_ net774 _02552_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_16244_ CPU.registerFile\[16\]\[5\] _03848_ _03769_ _03965_ VGND VGND VPWR VPWR _03966_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13456_ _08265_ VGND VGND VPWR VPWR _08416_ sky130_fd_sc_hd__buf_4
XFILLER_0_125_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10668_ CPU.registerFile\[1\]\[7\] _06386_ _06799_ VGND VGND VPWR VPWR _06804_ sky130_fd_sc_hd__mux2_1
X_13567__953 clknet_1_0__leaf__08442_ VGND VGND VPWR VPWR net1009 sky130_fd_sc_hd__inv_2
X_12407_ _07888_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16175_ CPU.registerFile\[13\]\[4\] _03709_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__or2_1
X_10599_ _06766_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13387_ CPU.state\[1\] _05703_ VGND VGND VPWR VPWR _08371_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15126_ _03133_ _03182_ _03187_ _03188_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__o211a_1
X_12338_ _06603_ net1937 _07848_ VGND VGND VPWR VPWR _07852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15057_ CPU.registerFile\[21\]\[18\] _02960_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__or2_1
X_12269_ mapped_spi_ram.rcv_data\[14\] _07800_ VGND VGND VPWR VPWR _07808_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18816_ net605 _02340_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_18747_ net536 _02271_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[9\] sky130_fd_sc_hd__dfxtp_1
X_09480_ mapped_spi_ram.rcv_data\[2\] _05685_ _05698_ mapped_spi_flash.rcv_data\[2\]
+ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__a22o_1
X_18678_ net467 _02202_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17629_ net1663 VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15943__681 clknet_1_0__leaf__03689_ VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__inv_2
XFILLER_0_86_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17392__16 clknet_1_0__leaf__04985_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__inv_2
XFILLER_0_160_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15642__442 clknet_1_0__leaf__03642_ VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__inv_2
XFILLER_0_160_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14137__277 clknet_1_0__leaf__08498_ VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__inv_2
X_09816_ _06152_ _05990_ VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__xnor2_1
X_13694__1068 clknet_1_1__leaf__08454_ VGND VGND VPWR VPWR net1124 sky130_fd_sc_hd__inv_2
X_09747_ CPU.PC\[18\] _05891_ CPU.PC\[19\] VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__a21oi_1
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _06017_ _06018_ _06020_ _05516_ VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15725__517 clknet_1_1__leaf__03650_ VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__inv_2
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11640_ net1986 _07358_ _07438_ VGND VGND VPWR VPWR _07441_ sky130_fd_sc_hd__mux2_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_866 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11571_ net2074 _07358_ _07401_ VGND VGND VPWR VPWR _07404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18580__37 VGND VGND VPWR VPWR _18580__37/HI net37 sky130_fd_sc_hd__conb_1
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10522_ _06725_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__clkbuf_1
X_14290_ _08409_ VGND VGND VPWR VPWR _08536_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_134_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10453_ _06688_ VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10384_ _06647_ net1849 _06639_ VGND VGND VPWR VPWR _06648_ sky130_fd_sc_hd__mux2_1
X_13172_ _08295_ _08296_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12123_ mapped_spi_ram.cmd_addr\[22\] _05671_ _07704_ VGND VGND VPWR VPWR _07709_
+ sky130_fd_sc_hd__mux2_2
X_17980_ net991 _01508_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_16931_ CPU.registerFile\[2\]\[22\] CPU.registerFile\[3\]\[22\] _04431_ VGND VGND
+ VPWR VPWR _04636_ sky130_fd_sc_hd__mux2_1
X_12054_ _07661_ VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__clkbuf_1
X_11005_ _06982_ VGND VGND VPWR VPWR _07048_ sky130_fd_sc_hd__clkbuf_2
X_16862_ _06148_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__clkbuf_4
X_18601_ net422 _02125_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_15813_ net1598 _08357_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__nand2_1
X_16793_ CPU.aluIn1\[18\] _04458_ _04501_ _04259_ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__o211a_1
X_18532_ net353 _02056_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12956_ _07414_ _06775_ VGND VGND VPWR VPWR _08180_ sky130_fd_sc_hd__nor2_2
XFILLER_0_158_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18463_ net284 _01991_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_11907_ _06636_ net1887 _07573_ VGND VGND VPWR VPWR _07583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15675_ clknet_1_0__leaf__03643_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__buf_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _08143_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ CPU.registerFile\[5\]\[7\] CPU.registerFile\[4\]\[7\] _08864_ VGND VGND VPWR
+ VPWR _08865_ sky130_fd_sc_hd__mux2_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _07546_ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__clkbuf_1
X_18394_ net215 _01922_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ CPU.registerFile\[16\]\[6\] _08412_ _08796_ _06037_ VGND VGND VPWR VPWR _08797_
+ sky130_fd_sc_hd__o211a_1
X_11769_ _06634_ net2300 _07501_ VGND VGND VPWR VPWR _07510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__08510_ clknet_0__08510_ VGND VGND VPWR VPWR clknet_1_1__leaf__08510_
+ sky130_fd_sc_hd__clkbuf_16
X_17276_ CPU.registerFile\[19\]\[31\] CPU.registerFile\[18\]\[31\] _03745_ VGND VGND
+ VPWR VPWR _04972_ sky130_fd_sc_hd__mux2_1
X_14488_ _08722_ _08725_ _08729_ _08554_ VGND VGND VPWR VPWR _08730_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_858 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19015_ net757 _02535_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_16227_ _08404_ _03935_ _03939_ _03948_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__a31o_2
XFILLER_0_130_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08441_ clknet_0__08441_ VGND VGND VPWR VPWR clknet_1_1__leaf__08441_
+ sky130_fd_sc_hd__clkbuf_16
X_13439_ _08402_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08472_ _08472_ VGND VGND VPWR VPWR clknet_0__08472_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13348__844 clknet_1_1__leaf__08367_ VGND VGND VPWR VPWR net900 sky130_fd_sc_hd__inv_2
X_16158_ CPU.registerFile\[22\]\[3\] CPU.registerFile\[23\]\[3\] _03759_ VGND VGND
+ VPWR VPWR _03882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15109_ _06062_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__buf_4
XFILLER_0_11_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16089_ _03692_ _03795_ _03814_ _03601_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__a211o_1
X_08980_ CPU.aluIn1\[14\] _05330_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__nor2_1
X_09601_ CPU.Bimm\[9\] _05914_ CPU.PC\[9\] VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__a21o_1
X_09532_ _05875_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09463_ _05399_ _05810_ VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09394_ _05744_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__buf_4
XFILLER_0_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13288__791 clknet_1_0__leaf__08345_ VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__inv_2
XFILLER_0_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14070__217 clknet_1_1__leaf__08491_ VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__08461_ clknet_0__08461_ VGND VGND VPWR VPWR clknet_1_0__leaf__08461_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12810_ CPU.aluShamt\[2\] CPU.aluShamt\[1\] CPU.aluShamt\[0\] net2433 VGND VGND VPWR
+ VPWR _08102_ sky130_fd_sc_hd__o31a_1
XFILLER_0_158_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _06593_ net2056 _08065_ VGND VGND VPWR VPWR _08066_ sky130_fd_sc_hd__mux2_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15460_ CPU.registerFile\[13\]\[28\] CPU.registerFile\[12\]\[28\] _08794_ VGND VGND
+ VPWR VPWR _03514_ sky130_fd_sc_hd__mux2_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _08028_ VGND VGND VPWR VPWR _08029_ sky130_fd_sc_hd__buf_4
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ CPU.registerFile\[15\]\[2\] CPU.registerFile\[14\]\[2\] _08558_ VGND VGND
+ VPWR VPWR _08655_ sky130_fd_sc_hd__mux2_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11623_ net2236 _07341_ _07427_ VGND VGND VPWR VPWR _07432_ sky130_fd_sc_hd__mux2_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15391_ _03138_ _03139_ CPU.registerFile\[9\]\[26\] VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__a21o_1
XFILLER_0_154_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_22_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_16
X_17130_ CPU.registerFile\[20\]\[27\] CPU.registerFile\[21\]\[27\] _03737_ VGND VGND
+ VPWR VPWR _04830_ sky130_fd_sc_hd__mux2_1
X_14342_ _08549_ VGND VGND VPWR VPWR _08588_ sky130_fd_sc_hd__buf_4
X_11554_ net1732 _07341_ _07390_ VGND VGND VPWR VPWR _07395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_858 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17061_ _04579_ _04580_ CPU.registerFile\[17\]\[25\] VGND VGND VPWR VPWR _04763_
+ sky130_fd_sc_hd__a21o_1
X_10505_ _06716_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__clkbuf_1
X_14273_ _08415_ _08516_ _08518_ _08420_ VGND VGND VPWR VPWR _08519_ sky130_fd_sc_hd__a211o_1
X_11485_ _07352_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16012_ _03736_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__clkbuf_8
X_13224_ _08335_ _06522_ _08336_ _08337_ _08332_ VGND VGND VPWR VPWR _08338_ sky130_fd_sc_hd__o221ai_1
X_10436_ _06679_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17337__749 clknet_1_1__leaf__04983_ VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__inv_2
X_13155_ _08285_ net1554 VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__nor2_1
X_10367_ _06266_ VGND VGND VPWR VPWR _06636_ sky130_fd_sc_hd__buf_4
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12106_ net1365 _07693_ _07698_ _07175_ VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__o211a_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ CPU.registerFile\[4\]\[2\] _06507_ _08239_ VGND VGND VPWR VPWR _08249_ sky130_fd_sc_hd__mux2_1
X_17963_ net974 _01491_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_10298_ _06589_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__clkbuf_1
X_12037_ _07652_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__clkbuf_1
X_16914_ CPU.registerFile\[16\]\[21\] _04252_ _04494_ _04619_ VGND VGND VPWR VPWR
+ _04620_ sky130_fd_sc_hd__o211a_1
X_17894_ clknet_leaf_9_clk _01422_ VGND VGND VPWR VPWR CPU.aluWr sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16845_ CPU.registerFile\[13\]\[20\] _04380_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__or2_1
X_16776_ _05690_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18515_ net336 _02039_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12939_ _08171_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__clkbuf_1
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18446_ net267 _01974_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14609_ _08808_ _08809_ CPU.registerFile\[25\]\[7\] VGND VGND VPWR VPWR _08848_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18377_ net198 _01905_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13693__1067 clknet_1_1__leaf__08454_ VGND VGND VPWR VPWR net1123 sky130_fd_sc_hd__inv_2
X_17259_ CPU.registerFile\[2\]\[31\] CPU.registerFile\[3\]\[31\] _03759_ VGND VGND
+ VPWR VPWR _04955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__08455_ _08455_ VGND VGND VPWR VPWR clknet_0__08455_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15754__543 clknet_1_0__leaf__03653_ VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__inv_2
X_08963_ _05314_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08894_ _05245_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__clkbuf_4
X_14249__378 clknet_1_1__leaf__08509_ VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__inv_2
X_09515_ _05859_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_149_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09446_ _05410_ _05402_ _05407_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__and3_1
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09377_ CPU.instr\[6\] _05243_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11270_ _07228_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__clkbuf_1
X_10221_ _05420_ _05410_ _05408_ VGND VGND VPWR VPWR _06542_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10152_ _06392_ _06472_ _06475_ _05555_ VGND VGND VPWR VPWR _06476_ sky130_fd_sc_hd__a22o_1
X_14960_ _08580_ VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__clkbuf_4
X_10083_ _05298_ _05769_ _05770_ CPU.aluReg\[6\] _06409_ VGND VGND VPWR VPWR _06410_
+ sky130_fd_sc_hd__a221o_1
Xhold9 mapped_spi_ram.rcv_bitcount\[4\] VGND VGND VPWR VPWR net1306 sky130_fd_sc_hd__dlygate4sd3_1
X_14891_ CPU.registerFile\[22\]\[14\] CPU.registerFile\[23\]\[14\] _08756_ VGND VGND
+ VPWR VPWR _02959_ sky130_fd_sc_hd__mux2_1
X_16630_ CPU.registerFile\[12\]\[15\] _04017_ _04018_ _04341_ VGND VGND VPWR VPWR
+ _04342_ sky130_fd_sc_hd__o211a_1
X_13842_ clknet_1_1__leaf__08462_ VGND VGND VPWR VPWR _08469_ sky130_fd_sc_hd__buf_1
X_15883__627 clknet_1_0__leaf__03683_ VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__08444_ clknet_0__08444_ VGND VGND VPWR VPWR clknet_1_0__leaf__08444_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16561_ _03901_ _04270_ _04274_ _04072_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__o211a_1
X_10985_ _05643_ VGND VGND VPWR VPWR _07031_ sky130_fd_sc_hd__buf_2
X_18300_ net121 _01828_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_15512_ _06339_ _03547_ _03564_ _03243_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__a211o_2
X_12724_ _08056_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__clkbuf_1
X_16492_ _06141_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18231_ net1242 _01759_ VGND VGND VPWR VPWR mapped_spi_flash.div_counter\[0\] sky130_fd_sc_hd__dfxtp_1
X_15443_ CPU.registerFile\[17\]\[28\] _08528_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__or2_1
X_12655_ _06647_ net1945 _08015_ VGND VGND VPWR VPWR _08020_ sky130_fd_sc_hd__mux2_1
X_13981__137 clknet_1_0__leaf__08482_ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__inv_2
XFILLER_0_38_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11606_ net1998 _07324_ _07416_ VGND VGND VPWR VPWR _07423_ sky130_fd_sc_hd__mux2_1
X_18162_ net1173 _01690_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15374_ CPU.registerFile\[22\]\[26\] CPU.registerFile\[23\]\[26\] _08584_ VGND VGND
+ VPWR VPWR _03430_ sky130_fd_sc_hd__mux2_1
X_12586_ _07983_ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17113_ CPU.registerFile\[5\]\[27\] CPU.registerFile\[4\]\[27\] _03697_ VGND VGND
+ VPWR VPWR _04813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14325_ CPU.registerFile\[8\]\[0\] _08526_ _08570_ _06036_ VGND VGND VPWR VPWR _08571_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18093_ net1104 _01621_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_11537_ net1773 _07324_ _07379_ VGND VGND VPWR VPWR _07386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17044_ _04389_ _04390_ CPU.registerFile\[1\]\[25\] VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__a21o_1
Xhold409 CPU.registerFile\[28\]\[23\] VGND VGND VPWR VPWR net1706 sky130_fd_sc_hd__dlygate4sd3_1
X_15703__497 clknet_1_1__leaf__03648_ VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__inv_2
XFILLER_0_34_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11468_ _06144_ VGND VGND VPWR VPWR _07341_ sky130_fd_sc_hd__buf_4
Xclkbuf_1_1__f__03682_ clknet_0__03682_ VGND VGND VPWR VPWR clknet_1_1__leaf__03682_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13207_ _06018_ _06096_ _08312_ _08320_ VGND VGND VPWR VPWR _08321_ sky130_fd_sc_hd__or4_1
X_10419_ _06670_ VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11399_ _07297_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ net1622 _08275_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__xor2_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ clknet_leaf_14_clk _02515_ VGND VGND VPWR VPWR CPU.aluIn1\[12\] sky130_fd_sc_hd__dfxtp_4
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ net1397 VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__clkbuf_1
X_17946_ net957 _01474_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[16\] sky130_fd_sc_hd__dfxtp_1
Xhold1109 CPU.registerFile\[3\]\[24\] VGND VGND VPWR VPWR net2406 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_16
X_17877_ clknet_leaf_17_clk _00027_ VGND VGND VPWR VPWR CPU.cycles\[20\] sky130_fd_sc_hd__dfxtp_1
X_16828_ _04534_ _04535_ _04365_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16759_ CPU.registerFile\[6\]\[18\] CPU.registerFile\[7\]\[18\] _04426_ VGND VGND
+ VPWR VPWR _04468_ sky130_fd_sc_hd__mux2_1
X_09300_ CPU.PC\[23\] VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09231_ _05575_ _05581_ _05582_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18429_ net250 _01957_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09162_ CPU.Jimm\[14\] VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__buf_4
XFILLER_0_56_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09093_ _05432_ _05444_ _05290_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold910 CPU.registerFile\[3\]\[25\] VGND VGND VPWR VPWR net2207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 CPU.registerFile\[3\]\[15\] VGND VGND VPWR VPWR net2218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold932 CPU.registerFile\[7\]\[14\] VGND VGND VPWR VPWR net2229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08507_ _08507_ VGND VGND VPWR VPWR clknet_0__08507_ sky130_fd_sc_hd__clkbuf_16
X_15678__474 clknet_1_0__leaf__03646_ VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__inv_2
XFILLER_0_40_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold943 CPU.registerFile\[6\]\[5\] VGND VGND VPWR VPWR net2240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold954 CPU.registerFile\[27\]\[24\] VGND VGND VPWR VPWR net2251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold965 CPU.registerFile\[21\]\[28\] VGND VGND VPWR VPWR net2262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 CPU.registerFile\[8\]\[1\] VGND VGND VPWR VPWR net2273 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__08438_ _08438_ VGND VGND VPWR VPWR clknet_0__08438_ sky130_fd_sc_hd__clkbuf_16
Xhold987 CPU.registerFile\[29\]\[29\] VGND VGND VPWR VPWR net2284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 CPU.registerFile\[16\]\[17\] VGND VGND VPWR VPWR net2295 sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ _05818_ _06320_ _06323_ _06324_ _05308_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__a32o_1
X_13246__767 clknet_1_1__leaf__08343_ VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__inv_2
Xclkbuf_0__08369_ _08369_ VGND VGND VPWR VPWR clknet_0__08369_ sky130_fd_sc_hd__clkbuf_16
X_08946_ CPU.aluIn1\[6\] _05297_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__and2_1
X_14182__318 clknet_1_1__leaf__08502_ VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__inv_2
X_10770_ CPU.aluShamt\[4\] _06859_ VGND VGND VPWR VPWR _06864_ sky130_fd_sc_hd__nor2_2
XFILLER_0_66_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09429_ _05776_ _05777_ _05778_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12440_ _07905_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12371_ _06636_ net1825 _07859_ VGND VGND VPWR VPWR _07869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11322_ _07256_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15090_ _02750_ _03132_ _03153_ _02839_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__a211o_1
XFILLER_0_132_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14002__155 clknet_1_1__leaf__08485_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__inv_2
XFILLER_0_160_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11253_ _07219_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__clkbuf_1
X_13561__948 clknet_1_0__leaf__08441_ VGND VGND VPWR VPWR net1004 sky130_fd_sc_hd__inv_2
X_10204_ _05274_ _05528_ VGND VGND VPWR VPWR _06526_ sky130_fd_sc_hd__and2_1
X_11184_ mapped_spi_flash.div_counter\[3\] mapped_spi_flash.div_counter\[2\] mapped_spi_flash.div_counter\[5\]
+ mapped_spi_flash.div_counter\[4\] VGND VGND VPWR VPWR _07176_ sky130_fd_sc_hd__or4_1
X_17800_ net880 _01362_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_10135_ mapped_spi_ram.rcv_data\[28\] _05857_ VGND VGND VPWR VPWR _06460_ sky130_fd_sc_hd__and2_1
X_18780_ net569 _02304_ VGND VGND VPWR VPWR CPU.aluReg\[10\] sky130_fd_sc_hd__dfxtp_1
X_15992_ CPU.registerFile\[5\]\[0\] CPU.registerFile\[4\]\[0\] _03704_ VGND VGND VPWR
+ VPWR _03719_ sky130_fd_sc_hd__mux2_1
X_17731_ net816 _01297_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_14943_ _03006_ _03007_ _03009_ _02814_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__a211o_2
X_10066_ _05526_ _05696_ VGND VGND VPWR VPWR _06393_ sky130_fd_sc_hd__nor2_2
X_13692__1066 clknet_1_0__leaf__08454_ VGND VGND VPWR VPWR net1122 sky130_fd_sc_hd__inv_2
XFILLER_0_82_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17662_ _05195_ _05192_ _05196_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__and3b_1
X_14874_ _02728_ _02938_ _02942_ _02784_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16613_ _04324_ _04325_ _03961_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17593_ per_uart.uart0.tx_bitcount\[1\] per_uart.uart0.tx_bitcount\[0\] _05147_ VGND
+ VGND VPWR VPWR _05152_ sky130_fd_sc_hd__and3_1
XFILLER_0_159_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16544_ _06855_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__buf_2
XFILLER_0_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10968_ mapped_spi_flash.cmd_addr\[17\] _05663_ _07009_ VGND VGND VPWR VPWR _07017_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12707_ _08047_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__clkbuf_1
X_16475_ _04015_ _04188_ _04190_ _03979_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__a211o_1
X_13687_ clknet_1_1__leaf__08451_ VGND VGND VPWR VPWR _08454_ sky130_fd_sc_hd__buf_1
X_10899_ CPU.aluReg\[3\] CPU.aluReg\[1\] _06939_ VGND VGND VPWR VPWR _06964_ sky130_fd_sc_hd__mux2_1
X_13630__1011 clknet_1_1__leaf__08447_ VGND VGND VPWR VPWR net1067 sky130_fd_sc_hd__inv_2
X_15426_ CPU.registerFile\[10\]\[27\] CPU.registerFile\[11\]\[27\] _03183_ VGND VGND
+ VPWR VPWR _03481_ sky130_fd_sc_hd__mux2_1
X_18214_ net1225 _01742_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[15\] sky130_fd_sc_hd__dfxtp_1
X_19194_ net104 net1481 VGND VGND VPWR VPWR mapped_spi_ram.div_counter\[1\] sky130_fd_sc_hd__dfxtp_1
X_12638_ _06630_ net1878 _08004_ VGND VGND VPWR VPWR _08011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18145_ net1156 _01673_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_15357_ _03098_ _03411_ _03413_ _03307_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__a211o_1
X_12569_ _07974_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14308_ _08422_ VGND VGND VPWR VPWR _08554_ sky130_fd_sc_hd__buf_4
XFILLER_0_103_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18076_ net1087 _01604_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_15288_ _03345_ _03346_ _03025_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__mux2_1
Xhold206 _00039_ VGND VGND VPWR VPWR net1503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 per_uart.uart0.enable16_counter\[1\] VGND VGND VPWR VPWR net1514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold228 mapped_spi_flash.cmd_addr\[16\] VGND VGND VPWR VPWR net1525 sky130_fd_sc_hd__dlygate4sd3_1
X_17027_ _04367_ _04727_ _04729_ _04410_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__a211o_1
XFILLER_0_150_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold239 mapped_spi_ram.rcv_data\[15\] VGND VGND VPWR VPWR net1536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _05881_ _06111_ _06118_ _05540_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_147_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18978_ net752 _02498_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ net940 _01457_ VGND VGND VPWR VPWR CPU.aluShamt\[4\] sky130_fd_sc_hd__dfxtp_1
X_13538__928 clknet_1_1__leaf__08438_ VGND VGND VPWR VPWR net984 sky130_fd_sc_hd__inv_2
XFILLER_0_48_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09214_ _05564_ _05565_ VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09145_ _05366_ _05486_ _05489_ _05496_ VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09076_ _05293_ CPU.aluIn1\[7\] VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__or2b_1
XFILLER_0_102_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold740 CPU.registerFile\[13\]\[3\] VGND VGND VPWR VPWR net2037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 CPU.registerFile\[12\]\[25\] VGND VGND VPWR VPWR net2048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 CPU.registerFile\[11\]\[19\] VGND VGND VPWR VPWR net2059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 CPU.registerFile\[8\]\[27\] VGND VGND VPWR VPWR net2070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 CPU.registerFile\[9\]\[27\] VGND VGND VPWR VPWR net2081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 CPU.registerFile\[2\]\[23\] VGND VGND VPWR VPWR net2092 sky130_fd_sc_hd__dlygate4sd3_1
X_09978_ CPU.cycles\[10\] _05553_ _06197_ _06308_ VGND VGND VPWR VPWR _06309_ sky130_fd_sc_hd__o2bb2a_1
X_08929_ CPU.aluIn1\[0\] _05274_ _05276_ _05280_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__a31o_1
X_11940_ _06601_ net2245 _07598_ VGND VGND VPWR VPWR _07601_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _07564_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__clkbuf_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03685_ clknet_0__03685_ VGND VGND VPWR VPWR clknet_1_0__leaf__03685_
+ sky130_fd_sc_hd__clkbuf_16
X_10822_ _06905_ VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__clkbuf_1
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _08574_ _08825_ _08829_ _08592_ VGND VGND VPWR VPWR _08830_ sky130_fd_sc_hd__o211a_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10753_ net2477 _06555_ _06815_ VGND VGND VPWR VPWR _06850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16260_ CPU.registerFile\[6\]\[6\] CPU.registerFile\[7\]\[6\] _03717_ VGND VGND VPWR
+ VPWR _03981_ sky130_fd_sc_hd__mux2_1
X_13472_ _08427_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__clkbuf_1
X_10684_ CPU.Bimm\[1\] CPU.Bimm\[11\] CPU.writeBack VGND VGND VPWR VPWR _06812_ sky130_fd_sc_hd__or3b_1
XFILLER_0_152_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15211_ CPU.registerFile\[6\]\[21\] CPU.registerFile\[7\]\[21\] _02982_ VGND VGND
+ VPWR VPWR _03272_ sky130_fd_sc_hd__mux2_1
X_12423_ net1742 _07335_ _07895_ VGND VGND VPWR VPWR _07897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16191_ CPU.registerFile\[27\]\[4\] CPU.registerFile\[26\]\[4\] _03837_ VGND VGND
+ VPWR VPWR _03914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15142_ CPU.registerFile\[17\]\[20\] _03036_ VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__or2_1
X_12354_ _07860_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__clkbuf_1
X_11305_ _07247_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__clkbuf_1
X_15073_ CPU.registerFile\[10\]\[18\] CPU.registerFile\[11\]\[18\] _02779_ VGND VGND
+ VPWR VPWR _03137_ sky130_fd_sc_hd__mux2_1
X_12285_ net1454 _07812_ _07817_ _07809_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18901_ net675 _02421_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11236_ _07210_ VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__clkbuf_1
X_18832_ net621 _02356_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_11167_ _05679_ _07132_ VGND VGND VPWR VPWR _07167_ sky130_fd_sc_hd__nand2_1
X_10118_ _05290_ _05432_ _05444_ _06442_ VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__a31o_1
X_18763_ net552 net1531 VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[25\] sky130_fd_sc_hd__dfxtp_1
X_15975_ _08396_ VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__clkbuf_8
X_11098_ _07118_ _07123_ _07120_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17714_ _07001_ _05233_ VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__and2_1
X_14926_ net1636 _02797_ _02992_ _02993_ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__o211a_1
X_10049_ _05555_ _05294_ _05295_ _05526_ _05799_ VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__a2111oi_1
X_18694_ net483 _02218_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_bitcount\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14165__302 clknet_1_0__leaf__08501_ VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__inv_2
X_17645_ net2624 _08360_ _05184_ _07002_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__o211a_1
X_14857_ _02924_ _02925_ _02851_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__mux2_1
X_18586__43 VGND VGND VPWR VPWR _18586__43/HI net43 sky130_fd_sc_hd__conb_1
X_14788_ CPU.registerFile\[15\]\[11\] CPU.registerFile\[14\]\[11\] _08771_ VGND VGND
+ VPWR VPWR _02859_ sky130_fd_sc_hd__mux2_1
X_17576_ per_uart.uart0.tx_count16\[1\] per_uart.uart0.tx_count16\[0\] _05137_ _05138_
+ per_uart.uart0.tx_count16\[2\] VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__a32o_1
XFILLER_0_147_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16527_ _03744_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16458_ _03748_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15409_ _03156_ _03461_ _03463_ _03163_ VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__a211o_1
X_19177_ clknet_leaf_6_clk net1632 VGND VGND VPWR VPWR per_uart.uart0.rx_bitcount\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16389_ CPU.registerFile\[15\]\[9\] CPU.registerFile\[14\]\[9\] _03705_ VGND VGND
+ VPWR VPWR _04107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18128_ net1139 _01656_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18059_ net1070 _01587_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09901_ _05939_ _05979_ VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03648_ clknet_0__03648_ VGND VGND VPWR VPWR clknet_1_1__leaf__03648_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09832_ _06168_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__buf_4
Xclkbuf_0__03679_ _03679_ VGND VGND VPWR VPWR clknet_0__03679_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_158_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _05925_ _05995_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__xnor2_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13850__1209 clknet_1_1__leaf__08469_ VGND VGND VPWR VPWR net1265 sky130_fd_sc_hd__inv_2
X_09694_ _06035_ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__clkbuf_8
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13319__819 clknet_1_1__leaf__08363_ VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__inv_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13590__974 clknet_1_1__leaf__08444_ VGND VGND VPWR VPWR net1030 sky130_fd_sc_hd__inv_2
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15920__660 clknet_1_0__leaf__03687_ VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__inv_2
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09128_ _05345_ CPU.aluIn1\[17\] VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__and2b_1
X_13691__1065 clknet_1_0__leaf__08454_ VGND VGND VPWR VPWR net1121 sky130_fd_sc_hd__inv_2
XFILLER_0_60_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09059_ _05402_ _05407_ _05408_ _05410_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_32_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12070_ _07669_ VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__clkbuf_1
Xhold570 CPU.registerFile\[27\]\[4\] VGND VGND VPWR VPWR net1867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 CPU.registerFile\[27\]\[15\] VGND VGND VPWR VPWR net1878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 CPU.registerFile\[17\]\[30\] VGND VGND VPWR VPWR net1889 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ _07048_ _07062_ VGND VGND VPWR VPWR _07063_ sky130_fd_sc_hd__or2_1
X_14114__256 clknet_1_0__leaf__08496_ VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__inv_2
X_12972_ net2406 _07326_ _08181_ VGND VGND VPWR VPWR _08189_ sky130_fd_sc_hd__mux2_1
Xhold1270 CPU.registerFile\[20\]\[2\] VGND VGND VPWR VPWR net2567 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_466 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14711_ _08422_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__clkbuf_4
Xhold1281 CPU.registerFile\[9\]\[9\] VGND VGND VPWR VPWR net2578 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11923_ _07591_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__clkbuf_1
Xhold1292 CPU.registerFile\[23\]\[5\] VGND VGND VPWR VPWR net2589 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17430_ _05880_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__buf_2
X_14642_ CPU.registerFile\[21\]\[8\] _08718_ VGND VGND VPWR VPWR _08880_ sky130_fd_sc_hd__or2_1
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ net2562 _07366_ _07548_ VGND VGND VPWR VPWR _07555_ sky130_fd_sc_hd__mux2_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ CPU.aluReg\[25\] _06892_ _06889_ VGND VGND VPWR VPWR _06893_ sky130_fd_sc_hd__mux2_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14573_ _08722_ _08806_ _08812_ _08554_ VGND VGND VPWR VPWR _08813_ sky130_fd_sc_hd__o211a_1
X_17361_ _03659_ _04989_ _04990_ _04991_ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_95_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11785_ _07518_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__clkbuf_1
X_19100_ net83 _02620_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_16312_ _03901_ _04026_ _04031_ _03732_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__o211a_1
X_10736_ _06841_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__clkbuf_1
X_14008__161 clknet_1_0__leaf__08485_ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__inv_2
XFILLER_0_137_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19031_ net773 _02551_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16243_ _03770_ _03771_ CPU.registerFile\[17\]\[5\] VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__a21o_1
X_13455_ _08414_ VGND VGND VPWR VPWR _08415_ sky130_fd_sc_hd__clkbuf_4
X_13772__1139 clknet_1_0__leaf__08461_ VGND VGND VPWR VPWR net1195 sky130_fd_sc_hd__inv_2
X_10667_ _06803_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__clkbuf_1
X_14160__298 clknet_1_1__leaf__08500_ VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__inv_2
XFILLER_0_125_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12406_ net1675 _07318_ _07884_ VGND VGND VPWR VPWR _07888_ sky130_fd_sc_hd__mux2_1
X_16174_ CPU.registerFile\[15\]\[4\] CPU.registerFile\[14\]\[4\] _03705_ VGND VGND
+ VPWR VPWR _03897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10598_ net1906 _06386_ _06761_ VGND VGND VPWR VPWR _06766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15125_ _08422_ VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12337_ _07851_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15056_ CPU.registerFile\[22\]\[18\] CPU.registerFile\[23\]\[18\] _02998_ VGND VGND
+ VPWR VPWR _03120_ sky130_fd_sc_hd__mux2_1
X_12268_ net1496 _07799_ _07807_ _07796_ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__o211a_1
X_11219_ _06593_ net1974 _07201_ VGND VGND VPWR VPWR _07202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12199_ net8 net14 VGND VGND VPWR VPWR _07761_ sky130_fd_sc_hd__nand2_1
X_18815_ net604 _02339_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_18746_ net535 _02270_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[8\] sky130_fd_sc_hd__dfxtp_1
X_14909_ CPU.registerFile\[10\]\[14\] CPU.registerFile\[11\]\[14\] _02779_ VGND VGND
+ VPWR VPWR _02977_ sky130_fd_sc_hd__mux2_1
X_18677_ net466 _02201_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_17628_ per_uart.rx_data\[3\] net1662 _05170_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17559_ net6 _05121_ _05126_ _05237_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__a211o_1
XFILLER_0_128_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17721__1 clknet_1_0__leaf__08341_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__inv_2
XFILLER_0_144_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09815_ _05937_ _05986_ _05935_ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__a21o_1
X_09746_ _05856_ _06085_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__nand2_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _06017_ _06019_ VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__nand2_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13371__865 clknet_1_0__leaf__08369_ VGND VGND VPWR VPWR net921 sky130_fd_sc_hd__inv_2
X_11570_ _07403_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10521_ net2525 _06292_ _06724_ VGND VGND VPWR VPWR _06725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13240_ clknet_1_0__leaf__08341_ VGND VGND VPWR VPWR _08343_ sky130_fd_sc_hd__buf_1
XFILLER_0_45_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10452_ _06638_ net2529 _06687_ VGND VGND VPWR VPWR _06688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13171_ net1586 _08293_ VGND VGND VPWR VPWR _08296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10383_ _06385_ VGND VGND VPWR VPWR _06647_ sky130_fd_sc_hd__buf_4
XFILLER_0_131_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12122_ net1334 _07693_ _07708_ _07175_ VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__o211a_1
X_16930_ _04633_ _04634_ _04557_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__mux2_1
X_12053_ CPU.registerFile\[24\]\[8\] _07360_ _07657_ VGND VGND VPWR VPWR _07661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11004_ net1522 _07007_ _07047_ _07014_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__o211a_1
X_16861_ CPU.registerFile\[27\]\[20\] CPU.registerFile\[26\]\[20\] _04242_ VGND VGND
+ VPWR VPWR _04568_ sky130_fd_sc_hd__mux2_1
X_18600_ net421 _02124_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_15812_ _08357_ _03674_ _03661_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__a21oi_1
X_16792_ _04141_ _04478_ _04499_ _04500_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__a211o_1
X_18531_ net352 _02055_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_12955_ net1618 VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11906_ _07582_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18462_ net283 _01990_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15927__666 clknet_1_1__leaf__03688_ VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__inv_2
X_12886_ _06555_ net2104 _08108_ VGND VGND VPWR VPWR _08143_ sky130_fd_sc_hd__mux2_1
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14625_ _06062_ VGND VGND VPWR VPWR _08864_ sky130_fd_sc_hd__buf_4
X_11837_ net2583 _07349_ _07537_ VGND VGND VPWR VPWR _07546_ sky130_fd_sc_hd__mux2_1
X_18393_ net214 _01921_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ CPU.registerFile\[17\]\[6\] _08795_ VGND VGND VPWR VPWR _08796_ sky130_fd_sc_hd__or2_1
X_11768_ _07509_ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10719_ _06832_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14487_ _08543_ _08726_ _08728_ _08552_ VGND VGND VPWR VPWR _08729_ sky130_fd_sc_hd__a211o_1
X_17275_ _04969_ _04970_ _03742_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11699_ _07472_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__clkbuf_1
X_19014_ clknet_leaf_12_clk _02534_ VGND VGND VPWR VPWR CPU.aluIn1\[31\] sky130_fd_sc_hd__dfxtp_1
X_16226_ _03901_ _03942_ _03947_ _03732_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_1__f__08440_ clknet_0__08440_ VGND VGND VPWR VPWR clknet_1_1__leaf__08440_
+ sky130_fd_sc_hd__clkbuf_16
X_13438_ CPU.Jimm\[17\] _08401_ _08388_ VGND VGND VPWR VPWR _08402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__08471_ _08471_ VGND VGND VPWR VPWR clknet_0__08471_ sky130_fd_sc_hd__clkbuf_16
X_16157_ _03735_ _03876_ _03880_ _03755_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15108_ _03169_ _03170_ _02851_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__mux2_1
X_16088_ _03805_ _03813_ _08406_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15039_ CPU.registerFile\[6\]\[17\] CPU.registerFile\[7\]\[17\] _02982_ VGND VGND
+ VPWR VPWR _03104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17314__728 clknet_1_1__leaf__04981_ VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__inv_2
X_15672__469 clknet_1_1__leaf__03645_ VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__inv_2
X_09600_ CPU.Bimm\[10\] _05914_ CPU.PC\[10\] VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09531_ _05722_ _05723_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__and2_2
X_18729_ net518 _02253_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[29\] sky130_fd_sc_hd__dfxtp_1
X_13690__1064 clknet_1_0__leaf__08454_ VGND VGND VPWR VPWR net1120 sky130_fd_sc_hd__inv_2
X_09462_ _05385_ _05388_ _05808_ _05809_ _05403_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__o311a_1
XFILLER_0_65_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09393_ _05540_ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__clkbuf_4
X_14143__282 clknet_1_0__leaf__08499_ VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__inv_2
XFILLER_0_7_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13934__94 clknet_1_1__leaf__08478_ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__inv_2
XFILLER_0_10_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15731__522 clknet_1_0__leaf__03651_ VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__inv_2
X_17289__705 clknet_1_1__leaf__04979_ VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__inv_2
X_13596__980 clknet_1_0__leaf__08444_ VGND VGND VPWR VPWR net1036 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__08460_ clknet_0__08460_ VGND VGND VPWR VPWR clknet_1_0__leaf__08460_
+ sky130_fd_sc_hd__clkbuf_16
X_13771__1138 clknet_1_0__leaf__08461_ VGND VGND VPWR VPWR net1194 sky130_fd_sc_hd__inv_2
X_09729_ _05367_ _06069_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__nand2_1
X_12740_ _08064_ VGND VGND VPWR VPWR _08065_ sky130_fd_sc_hd__buf_4
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15649__449 clknet_1_1__leaf__03642_ VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__inv_2
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19196__54 VGND VGND VPWR VPWR _19196__54/HI net54 sky130_fd_sc_hd__conb_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14226__357 clknet_1_1__leaf__08507_ VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__inv_2
X_12671_ _07488_ _07633_ VGND VGND VPWR VPWR _08028_ sky130_fd_sc_hd__nand2_4
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _08515_ _08640_ _08644_ _08653_ VGND VGND VPWR VPWR _08654_ sky130_fd_sc_hd__a31o_1
X_11622_ _07431_ VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15390_ CPU.registerFile\[10\]\[26\] CPU.registerFile\[11\]\[26\] _03183_ VGND VGND
+ VPWR VPWR _03446_ sky130_fd_sc_hd__mux2_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14341_ _08585_ _08586_ CPU.registerFile\[1\]\[0\] VGND VGND VPWR VPWR _08587_ sky130_fd_sc_hd__a21o_1
X_11553_ _07394_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17060_ CPU.registerFile\[19\]\[25\] CPU.registerFile\[18\]\[25\] _03745_ VGND VGND
+ VPWR VPWR _04762_ sky130_fd_sc_hd__mux2_1
X_10504_ net2057 _06106_ _06713_ VGND VGND VPWR VPWR _06716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14272_ CPU.registerFile\[16\]\[0\] _08412_ _08517_ _06037_ VGND VGND VPWR VPWR _08518_
+ sky130_fd_sc_hd__o211a_1
X_11484_ net1863 _07351_ _07333_ VGND VGND VPWR VPWR _07352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16011_ CPU.registerFile\[30\]\[0\] CPU.registerFile\[31\]\[0\] _03737_ VGND VGND
+ VPWR VPWR _03738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13223_ _08334_ _06517_ VGND VGND VPWR VPWR _08337_ sky130_fd_sc_hd__nand2_1
X_10435_ _06622_ net2404 _06676_ VGND VGND VPWR VPWR _06679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13154_ CPU.cycles\[13\] _08283_ net1553 VGND VGND VPWR VPWR _08286_ sky130_fd_sc_hd__a21oi_1
X_10366_ _06635_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__clkbuf_1
X_12105_ net1372 _07694_ _07696_ VGND VGND VPWR VPWR _07698_ sky130_fd_sc_hd__a21o_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ net1440 VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__clkbuf_1
X_17962_ net973 _01490_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_10297_ net1872 _06486_ _06580_ VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12036_ CPU.registerFile\[24\]\[16\] _07343_ _07646_ VGND VGND VPWR VPWR _07652_
+ sky130_fd_sc_hd__mux2_1
X_16913_ _04579_ _04580_ CPU.registerFile\[17\]\[21\] VGND VGND VPWR VPWR _04619_
+ sky130_fd_sc_hd__a21o_1
X_17893_ clknet_leaf_26_clk _01421_ VGND VGND VPWR VPWR CPU.mem_wmask\[3\] sky130_fd_sc_hd__dfxtp_1
X_16844_ CPU.registerFile\[15\]\[20\] CPU.registerFile\[14\]\[20\] _04550_ VGND VGND
+ VPWR VPWR _04551_ sky130_fd_sc_hd__mux2_1
X_16775_ _05689_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18514_ net335 _02038_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ _06361_ net2354 _08167_ VGND VGND VPWR VPWR _08171_ sky130_fd_sc_hd__mux2_1
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15860__606 clknet_1_0__leaf__03681_ VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__inv_2
X_18445_ net266 _01973_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _08134_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14608_ CPU.registerFile\[27\]\[7\] CPU.registerFile\[26\]\[7\] _06063_ VGND VGND
+ VPWR VPWR _08847_ sky130_fd_sc_hd__mux2_1
X_18376_ net197 _01904_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14539_ _08557_ _08774_ _08779_ _08423_ VGND VGND VPWR VPWR _08780_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17258_ _04952_ _04953_ _03769_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16209_ _03693_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__buf_4
X_17189_ CPU.registerFile\[0\]\[29\] _04637_ _03741_ _04886_ VGND VGND VPWR VPWR _04887_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__08454_ _08454_ VGND VGND VPWR VPWR clknet_0__08454_ sky130_fd_sc_hd__clkbuf_16
X_08962_ CPU.aluIn1\[11\] _05312_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__nor2_1
X_08893_ _05244_ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09514_ _05698_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__buf_4
X_09445_ _05793_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__clkbuf_4
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09376_ _05520_ _05697_ _05726_ _05727_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__a31o_2
XFILLER_0_75_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15956__692 clknet_1_1__leaf__03691_ VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__inv_2
X_10220_ _05413_ _05509_ _05511_ VGND VGND VPWR VPWR _06541_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10151_ _06288_ _06393_ _06473_ _06395_ _06474_ VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__a32o_1
X_15655__453 clknet_1_1__leaf__03644_ VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__inv_2
X_10082_ _05555_ _05298_ _05299_ _05526_ _05799_ VGND VGND VPWR VPWR _06409_ sky130_fd_sc_hd__a2111oi_1
X_14890_ _02751_ _02955_ _02957_ _02759_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_0__f__08443_ clknet_0__08443_ VGND VGND VPWR VPWR clknet_1_0__leaf__08443_
+ sky130_fd_sc_hd__clkbuf_16
X_16560_ _03943_ _04271_ _04273_ _04117_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__a211o_1
X_13377__871 clknet_1_1__leaf__08369_ VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__inv_2
X_10984_ _05612_ _07029_ VGND VGND VPWR VPWR _07030_ sky130_fd_sc_hd__xnor2_1
X_15511_ _03555_ _03563_ _03241_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12723_ _06647_ net2644 _08051_ VGND VGND VPWR VPWR _08056_ sky130_fd_sc_hd__mux2_1
X_16491_ CPU.registerFile\[24\]\[11\] _03915_ _04165_ _04206_ VGND VGND VPWR VPWR
+ _04207_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18230_ net1241 _01758_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_38_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12654_ _08019_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__clkbuf_1
X_15442_ CPU.registerFile\[19\]\[28\] CPU.registerFile\[18\]\[28\] _03157_ VGND VGND
+ VPWR VPWR _03496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11605_ _07422_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18161_ net1172 _01689_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[0\] sky130_fd_sc_hd__dfxtp_2
X_12585_ net2305 _07360_ _07979_ VGND VGND VPWR VPWR _07983_ sky130_fd_sc_hd__mux2_1
X_15373_ _03156_ _03426_ _03428_ _03163_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__a211o_1
XFILLER_0_154_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17112_ CPU.registerFile\[6\]\[27\] CPU.registerFile\[7\]\[27\] _03847_ VGND VGND
+ VPWR VPWR _04812_ sky130_fd_sc_hd__mux2_1
X_14324_ _08567_ _08569_ CPU.registerFile\[9\]\[0\] VGND VGND VPWR VPWR _08570_ sky130_fd_sc_hd__a21o_1
X_11536_ _07385_ VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18092_ net1103 _01620_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17043_ CPU.registerFile\[2\]\[25\] CPU.registerFile\[3\]\[25\] _04431_ VGND VGND
+ VPWR VPWR _04745_ sky130_fd_sc_hd__mux2_1
X_11467_ _07340_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__03681_ clknet_0__03681_ VGND VGND VPWR VPWR clknet_1_1__leaf__03681_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_151_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13206_ _05863_ _06275_ _08318_ _08319_ VGND VGND VPWR VPWR _08320_ sky130_fd_sc_hd__or4_1
X_10418_ _06605_ net2160 _06665_ VGND VGND VPWR VPWR _06670_ sky130_fd_sc_hd__mux2_1
X_14186_ clknet_1_1__leaf__08495_ VGND VGND VPWR VPWR _08503_ sky130_fd_sc_hd__buf_1
X_11398_ net1798 _06292_ _07296_ VGND VGND VPWR VPWR _07297_ sky130_fd_sc_hd__mux2_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _08275_ _08276_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__nor2_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _06123_ VGND VGND VPWR VPWR _06624_ sky130_fd_sc_hd__clkbuf_4
X_18994_ clknet_leaf_14_clk _02514_ VGND VGND VPWR VPWR CPU.aluIn1\[11\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13913__75 clknet_1_0__leaf__08476_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__inv_2
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ CPU.registerFile\[4\]\[11\] _06291_ _08239_ VGND VGND VPWR VPWR _08240_ sky130_fd_sc_hd__mux2_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ net956 _01473_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_12019_ net2466 _07326_ _07635_ VGND VGND VPWR VPWR _07643_ sky130_fd_sc_hd__mux2_1
X_17876_ clknet_leaf_23_clk _00025_ VGND VGND VPWR VPWR CPU.cycles\[19\] sky130_fd_sc_hd__dfxtp_1
X_16827_ CPU.registerFile\[20\]\[19\] CPU.registerFile\[21\]\[19\] _04287_ VGND VGND
+ VPWR VPWR _04535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16758_ _04419_ _04464_ _04466_ _04383_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__a211o_1
XFILLER_0_159_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16689_ _04080_ _04081_ CPU.registerFile\[25\]\[16\] VGND VGND VPWR VPWR _04400_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09230_ CPU.aluIn1\[2\] _05574_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__and2_1
X_18428_ net249 _01956_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09161_ _05420_ _05512_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__xnor2_1
X_18359_ net180 _01887_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09092_ _05433_ _05441_ _05443_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__a21o_1
X_13649__1028 clknet_1_1__leaf__08449_ VGND VGND VPWR VPWR net1084 sky130_fd_sc_hd__inv_2
XFILLER_0_44_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13770__1137 clknet_1_0__leaf__08461_ VGND VGND VPWR VPWR net1193 sky130_fd_sc_hd__inv_2
Xhold900 CPU.registerFile\[22\]\[6\] VGND VGND VPWR VPWR net2197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 CPU.registerFile\[3\]\[27\] VGND VGND VPWR VPWR net2208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 CPU.registerFile\[7\]\[28\] VGND VGND VPWR VPWR net2219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__08506_ _08506_ VGND VGND VPWR VPWR clknet_0__08506_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold933 CPU.registerFile\[29\]\[1\] VGND VGND VPWR VPWR net2230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 CPU.registerFile\[29\]\[28\] VGND VGND VPWR VPWR net2241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 CPU.registerFile\[26\]\[17\] VGND VGND VPWR VPWR net2252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 CPU.registerFile\[16\]\[1\] VGND VGND VPWR VPWR net2263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__08437_ _08437_ VGND VGND VPWR VPWR clknet_0__08437_ sky130_fd_sc_hd__clkbuf_16
Xhold977 CPU.registerFile\[23\]\[22\] VGND VGND VPWR VPWR net2274 sky130_fd_sc_hd__dlygate4sd3_1
X_14255__383 clknet_1_1__leaf__08510_ VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__inv_2
X_09994_ _05265_ _05522_ _05749_ VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__o21ai_1
Xhold988 CPU.registerFile\[19\]\[9\] VGND VGND VPWR VPWR net2285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 CPU.registerFile\[18\]\[2\] VGND VGND VPWR VPWR net2296 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__08368_ _08368_ VGND VGND VPWR VPWR clknet_0__08368_ sky130_fd_sc_hd__clkbuf_16
X_08945_ CPU.mem_wdata\[6\] CPU.Bimm\[6\] _05245_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13515__907 clknet_1_1__leaf__08436_ VGND VGND VPWR VPWR net963 sky130_fd_sc_hd__inv_2
X_17413__35 clknet_1_1__leaf__05014_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__inv_2
X_09428_ _05776_ _05777_ _05425_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_136_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09359_ _05582_ _05575_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__or2b_1
X_17716__47 clknet_1_0__leaf__05015_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__inv_2
XFILLER_0_35_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12370_ _07868_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17342__3 clknet_1_1__leaf__04984_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__inv_2
X_11321_ net2501 _06200_ _07249_ VGND VGND VPWR VPWR _07256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11252_ _06630_ net2123 _07212_ VGND VGND VPWR VPWR _07219_ sky130_fd_sc_hd__mux2_1
X_10203_ _06519_ _05523_ VGND VGND VPWR VPWR _06525_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11183_ net3 _07132_ _07174_ _07175_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10134_ _06456_ _06395_ _06457_ _06458_ VGND VGND VPWR VPWR _06459_ sky130_fd_sc_hd__o2bb2a_1
X_15991_ CPU.registerFile\[6\]\[0\] CPU.registerFile\[7\]\[0\] _03717_ VGND VGND VPWR
+ VPWR _03718_ sky130_fd_sc_hd__mux2_1
X_17730_ net815 _01296_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_14942_ CPU.registerFile\[24\]\[15\] _02928_ _03008_ _02771_ VGND VGND VPWR VPWR
+ _03009_ sky130_fd_sc_hd__o211a_1
X_10065_ _06390_ _06391_ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__and2_1
X_17661_ per_uart.uart0.rx_bitcount\[0\] _05194_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__or2_1
X_14873_ _08857_ _02939_ _02941_ _02903_ VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16612_ CPU.registerFile\[20\]\[14\] CPU.registerFile\[21\]\[14\] _04287_ VGND VGND
+ VPWR VPWR _04325_ sky130_fd_sc_hd__mux2_1
X_17592_ _05236_ _05134_ net2026 VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_159_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16543_ _04141_ _04238_ _04257_ _04096_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__a211o_1
X_10967_ net1499 _07007_ _07016_ _07014_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12706_ _06630_ net2550 _08040_ VGND VGND VPWR VPWR _08047_ sky130_fd_sc_hd__mux2_1
X_16474_ CPU.registerFile\[12\]\[11\] _04017_ _04018_ _04189_ VGND VGND VPWR VPWR
+ _04190_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10898_ _06963_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__clkbuf_1
X_18213_ net1224 _01741_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15425_ _03478_ _03479_ _08541_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19193_ net103 _02711_ VGND VGND VPWR VPWR mapped_spi_ram.div_counter\[0\] sky130_fd_sc_hd__dfxtp_1
X_12637_ _08010_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18144_ net1155 _01672_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15356_ CPU.registerFile\[8\]\[25\] _08545_ _03412_ _03268_ VGND VGND VPWR VPWR _03413_
+ sky130_fd_sc_hd__o211a_1
X_12568_ CPU.registerFile\[12\]\[16\] _07343_ _07968_ VGND VGND VPWR VPWR _07974_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11519_ _07375_ VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__clkbuf_1
X_14307_ _08543_ _08544_ _08551_ _08552_ VGND VGND VPWR VPWR _08553_ sky130_fd_sc_hd__a211o_1
XFILLER_0_40_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18075_ net1086 _01603_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_15287_ CPU.registerFile\[5\]\[23\] CPU.registerFile\[4\]\[23\] _03105_ VGND VGND
+ VPWR VPWR _03346_ sky130_fd_sc_hd__mux2_1
X_12499_ net2185 _07343_ _07931_ VGND VGND VPWR VPWR _07937_ sky130_fd_sc_hd__mux2_1
Xhold207 mapped_spi_flash.cmd_addr\[14\] VGND VGND VPWR VPWR net1504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold218 mapped_spi_flash.cmd_addr\[18\] VGND VGND VPWR VPWR net1515 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold229 per_uart.uart0.enable16_counter\[9\] VGND VGND VPWR VPWR net1526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17026_ CPU.registerFile\[16\]\[24\] _04656_ _04494_ _04728_ VGND VGND VPWR VPWR
+ _04729_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18977_ net751 _02497_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ net939 _01456_ VGND VGND VPWR VPWR CPU.aluShamt\[3\] sky130_fd_sc_hd__dfxtp_1
X_17859_ clknet_leaf_22_clk _00037_ VGND VGND VPWR VPWR CPU.cycles\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09213_ CPU.aluIn1\[18\] _05543_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09144_ _05374_ _05494_ _05495_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13252__772 clknet_1_0__leaf__08344_ VGND VGND VPWR VPWR net828 sky130_fd_sc_hd__inv_2
XFILLER_0_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09075_ _05424_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold730 CPU.registerFile\[31\]\[28\] VGND VGND VPWR VPWR net2027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 CPU.registerFile\[27\]\[5\] VGND VGND VPWR VPWR net2038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold752 CPU.registerFile\[17\]\[1\] VGND VGND VPWR VPWR net2049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold763 CPU.registerFile\[17\]\[16\] VGND VGND VPWR VPWR net2060 sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 CPU.registerFile\[28\]\[6\] VGND VGND VPWR VPWR net2071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 CPU.registerFile\[9\]\[30\] VGND VGND VPWR VPWR net2082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 CPU.registerFile\[9\]\[0\] VGND VGND VPWR VPWR net2093 sky130_fd_sc_hd__dlygate4sd3_1
X_09977_ _05886_ _06307_ VGND VGND VPWR VPWR _06308_ sky130_fd_sc_hd__or2_1
X_08928_ _05277_ _05245_ _05278_ _05279_ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__a211oi_1
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _06599_ net2169 _07562_ VGND VGND VPWR VPWR _07564_ sky130_fd_sc_hd__mux2_1
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15767__554 clknet_1_0__leaf__03655_ VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__inv_2
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03684_ clknet_0__03684_ VGND VGND VPWR VPWR clknet_1_0__leaf__03684_
+ sky130_fd_sc_hd__clkbuf_16
X_10821_ CPU.aluReg\[21\] _06904_ _06889_ VGND VGND VPWR VPWR _06905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13885__1241 clknet_1_1__leaf__08472_ VGND VGND VPWR VPWR net1297 sky130_fd_sc_hd__inv_2
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10752_ _06849_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13471_ CPU.Bimm\[5\] _05841_ _08416_ VGND VGND VPWR VPWR _08427_ sky130_fd_sc_hd__mux2_1
X_10683_ _06811_ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__clkbuf_1
X_15210_ _03133_ _03265_ _03270_ _03188_ VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__o211a_1
X_12422_ _07896_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__clkbuf_1
X_16190_ _03911_ _03912_ _03875_ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12353_ _06617_ net1918 _07859_ VGND VGND VPWR VPWR _07860_ sky130_fd_sc_hd__mux2_1
X_15141_ CPU.registerFile\[19\]\[20\] CPU.registerFile\[18\]\[20\] _03157_ VGND VGND
+ VPWR VPWR _03203_ sky130_fd_sc_hd__mux2_1
X_11304_ net2092 _06010_ _07238_ VGND VGND VPWR VPWR _07247_ sky130_fd_sc_hd__mux2_1
X_15072_ _03134_ _03135_ _02937_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12284_ mapped_spi_ram.rcv_data\[8\] _07813_ VGND VGND VPWR VPWR _07817_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18900_ net674 _02420_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_11235_ _06613_ net1775 _07201_ VGND VGND VPWR VPWR _07210_ sky130_fd_sc_hd__mux2_1
X_18831_ net620 _02355_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_11166_ net1409 _07160_ _07166_ _07164_ VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10117_ _05794_ _05445_ VGND VGND VPWR VPWR _06442_ sky130_fd_sc_hd__nand2_1
X_18762_ net551 net1507 VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[24\] sky130_fd_sc_hd__dfxtp_1
X_15974_ _08398_ _03695_ _03700_ _08401_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__a211o_1
X_11097_ mapped_spi_flash.snd_bitcount\[0\] _07114_ net1661 VGND VGND VPWR VPWR _07123_
+ sky130_fd_sc_hd__o21ai_1
X_17713_ CPU.mem_wdata\[7\] per_uart.d_in_uart\[7\] _05218_ VGND VGND VPWR VPWR _05233_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14925_ _07163_ VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__clkbuf_4
X_10048_ _05425_ _06375_ VGND VGND VPWR VPWR _06376_ sky130_fd_sc_hd__nand2_1
X_18693_ net482 _02217_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_bitcount\[0\] sky130_fd_sc_hd__dfxtp_1
X_13648__1027 clknet_1_0__leaf__08449_ VGND VGND VPWR VPWR net1083 sky130_fd_sc_hd__inv_2
XFILLER_0_117_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold90 CPU.aluReg\[13\] VGND VGND VPWR VPWR net1387 sky130_fd_sc_hd__dlygate4sd3_1
X_17644_ _08360_ _05183_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__nand2_1
X_14856_ CPU.registerFile\[28\]\[13\] CPU.registerFile\[29\]\[13\] _02808_ VGND VGND
+ VPWR VPWR _02925_ sky130_fd_sc_hd__mux2_1
X_17575_ _03659_ _05133_ _05137_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__a21o_1
X_14787_ _02798_ _02844_ _02848_ _02857_ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__a31o_1
X_11999_ _07631_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__clkbuf_1
X_16526_ _04239_ _04240_ _03875_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16457_ CPU.registerFile\[19\]\[10\] CPU.registerFile\[18\]\[10\] _03923_ VGND VGND
+ VPWR VPWR _04174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15408_ CPU.registerFile\[16\]\[27\] _03159_ _03462_ _03161_ VGND VGND VPWR VPWR
+ _03463_ sky130_fd_sc_hd__o211a_1
X_19176_ clknet_leaf_6_clk _02696_ VGND VGND VPWR VPWR per_uart.uart0.rx_bitcount\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16388_ _04099_ _04100_ _04104_ _04105_ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18127_ net1138 _01655_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15339_ CPU.registerFile\[21\]\[25\] _02752_ VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18058_ net1069 _01586_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_13544__933 clknet_1_0__leaf__08439_ VGND VGND VPWR VPWR net989 sky130_fd_sc_hd__inv_2
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17009_ CPU.registerFile\[0\]\[24\] _04637_ _04472_ _04711_ VGND VGND VPWR VPWR _04712_
+ sky130_fd_sc_hd__o211a_1
X_09900_ _05323_ _05769_ _05770_ net1387 _06233_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__a221o_1
Xclkbuf_1_1__f__03647_ clknet_0__03647_ VGND VGND VPWR VPWR clknet_1_1__leaf__03647_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09831_ _05764_ _06151_ _06154_ _06167_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__a211o_4
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__03678_ _03678_ VGND VGND VPWR VPWR clknet_0__03678_ sky130_fd_sc_hd__clkbuf_16
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ CPU.Jimm\[19\] _05550_ _05790_ CPU.cycles\[19\] _06101_ VGND VGND VPWR VPWR
+ _06102_ sky130_fd_sc_hd__a221o_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09693_ mapped_spi_flash.rcv_data\[13\] _05698_ _06034_ VGND VGND VPWR VPWR _06035_
+ sky130_fd_sc_hd__a21oi_4
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09127_ _05339_ CPU.aluIn1\[16\] VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09058_ _05258_ _05409_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__nand2_2
XFILLER_0_4_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold560 CPU.registerFile\[6\]\[24\] VGND VGND VPWR VPWR net1857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 CPU.registerFile\[2\]\[20\] VGND VGND VPWR VPWR net1868 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ mapped_spi_flash.cmd_addr\[10\] _07061_ _07039_ VGND VGND VPWR VPWR _07062_
+ sky130_fd_sc_hd__mux2_1
Xhold582 CPU.registerFile\[21\]\[9\] VGND VGND VPWR VPWR net1879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 CPU.registerFile\[7\]\[29\] VGND VGND VPWR VPWR net1890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12971_ _08188_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__clkbuf_1
Xhold1260 CPU.registerFile\[1\]\[28\] VGND VGND VPWR VPWR net2557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14710_ _08857_ _02780_ _02782_ _08661_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__a211o_1
Xhold1271 CPU.registerFile\[25\]\[9\] VGND VGND VPWR VPWR net2568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1282 CPU.registerFile\[25\]\[26\] VGND VGND VPWR VPWR net2579 sky130_fd_sc_hd__dlygate4sd3_1
X_11922_ _06651_ net2494 _07584_ VGND VGND VPWR VPWR _07591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1293 CPU.PC\[9\] VGND VGND VPWR VPWR net2590 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ CPU.registerFile\[22\]\[8\] CPU.registerFile\[23\]\[8\] _08756_ VGND VGND
+ VPWR VPWR _08879_ sky130_fd_sc_hd__mux2_1
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _07554_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ CPU.aluIn1\[25\] _06891_ _06881_ VGND VGND VPWR VPWR _06892_ sky130_fd_sc_hd__mux2_1
X_17360_ per_uart.uart0.rx_bitcount\[3\] per_uart.uart0.rx_bitcount\[2\] per_uart.uart0.rx_bitcount\[1\]
+ per_uart.uart0.rx_bitcount\[0\] VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__or4_1
X_14572_ _08764_ _08807_ _08811_ _08552_ VGND VGND VPWR VPWR _08812_ sky130_fd_sc_hd__a211o_1
X_11784_ _06649_ net2041 _07512_ VGND VGND VPWR VPWR _07518_ sky130_fd_sc_hd__mux2_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16311_ _03943_ _04028_ _04030_ _03730_ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__a211o_1
X_10735_ net2452 _06337_ _06838_ VGND VGND VPWR VPWR _06841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19030_ net772 _02550_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_16242_ CPU.registerFile\[19\]\[5\] CPU.registerFile\[18\]\[5\] _03923_ VGND VGND
+ VPWR VPWR _03964_ sky130_fd_sc_hd__mux2_1
X_10666_ CPU.registerFile\[1\]\[8\] _06361_ _06799_ VGND VGND VPWR VPWR _06803_ sky130_fd_sc_hd__mux2_1
X_13454_ _06418_ VGND VGND VPWR VPWR _08414_ sky130_fd_sc_hd__buf_4
XFILLER_0_137_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12405_ _07887_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__clkbuf_1
X_16173_ _08398_ _03893_ _03895_ _08401_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__a211o_1
X_10597_ _06765_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15124_ _03098_ _03184_ _03186_ _02903_ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__a211o_1
X_12336_ _06601_ net1776 _07848_ VGND VGND VPWR VPWR _07851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12267_ mapped_spi_ram.rcv_data\[15\] _07800_ VGND VGND VPWR VPWR _07807_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15055_ _02751_ _03116_ _03118_ _02759_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11218_ _07200_ VGND VGND VPWR VPWR _07201_ sky130_fd_sc_hd__buf_4
X_12198_ mapped_spi_ram.snd_bitcount\[5\] _07704_ _07759_ _07671_ _07672_ VGND VGND
+ VPWR VPWR _07760_ sky130_fd_sc_hd__o32a_1
XFILLER_0_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11149_ net1962 _07147_ _07156_ _07151_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__o211a_1
X_18814_ net603 _02338_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_18745_ net534 _02269_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[7\] sky130_fd_sc_hd__dfxtp_1
X_14089__234 clknet_1_1__leaf__08493_ VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__inv_2
X_14908_ _02974_ _02975_ _02937_ VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__mux2_1
X_18676_ net465 _02200_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15888_ clknet_1_1__leaf__03654_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__buf_1
X_17627_ net1671 VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__clkbuf_1
X_14839_ CPU.registerFile\[2\]\[12\] CPU.registerFile\[3\]\[12\] _02871_ VGND VGND
+ VPWR VPWR _02909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17558_ net1451 _05123_ _05124_ _05125_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16509_ _04099_ _04221_ _04223_ _04105_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__a211o_1
X_17489_ _05016_ net2641 _05067_ _05068_ _05053_ VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__o221a_1
XFILLER_0_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19159_ clknet_leaf_5_clk net1479 VGND VGND VPWR VPWR per_uart.uart0.txd_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13884__1240 clknet_1_1__leaf__08472_ VGND VGND VPWR VPWR net1296 sky130_fd_sc_hd__inv_2
X_13325__824 clknet_1_0__leaf__08364_ VGND VGND VPWR VPWR net880 sky130_fd_sc_hd__inv_2
X_15950__687 clknet_1_1__leaf__03690_ VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__inv_2
X_09814_ _05855_ _06150_ VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__nand2_1
X_09745_ mapped_spi_ram.rcv_data\[11\] _05858_ _05860_ net1327 VGND VGND VPWR VPWR
+ _06085_ sky130_fd_sc_hd__a22oi_4
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _05379_ _05902_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__xnor2_2
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10520_ _06701_ VGND VGND VPWR VPWR _06724_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10451_ _06664_ VGND VGND VPWR VPWR _06687_ sky130_fd_sc_hd__buf_4
X_13647__1026 clknet_1_0__leaf__08449_ VGND VGND VPWR VPWR net1082 sky130_fd_sc_hd__inv_2
X_13170_ CPU.cycles\[21\] _08293_ VGND VGND VPWR VPWR _08295_ sky130_fd_sc_hd__and2_1
X_10382_ _06646_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12121_ _07696_ _07707_ VGND VGND VPWR VPWR _07708_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12052_ _07660_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold390 CPU.registerFile\[6\]\[6\] VGND VGND VPWR VPWR net1687 sky130_fd_sc_hd__dlygate4sd3_1
X_14038__188 clknet_1_1__leaf__08488_ VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__inv_2
X_11003_ _07008_ _07046_ VGND VGND VPWR VPWR _07047_ sky130_fd_sc_hd__or2_1
X_16860_ _04565_ _04566_ _04279_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__mux2_1
X_15811_ net1541 _08356_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__nand2_1
X_16791_ _08596_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18530_ net351 _02054_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_12954_ _06555_ CPU.registerFile\[31\]\[0\] _08144_ VGND VGND VPWR VPWR _08179_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1090 CPU.registerFile\[17\]\[7\] VGND VGND VPWR VPWR net2387 sky130_fd_sc_hd__dlygate4sd3_1
X_18461_ net282 _01989_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_11905_ _06634_ net1919 _07573_ VGND VGND VPWR VPWR _07582_ sky130_fd_sc_hd__mux2_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _08142_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__clkbuf_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ CPU.registerFile\[6\]\[7\] CPU.registerFile\[7\]\[7\] _08740_ VGND VGND VPWR
+ VPWR _08863_ sky130_fd_sc_hd__mux2_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _07545_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__clkbuf_1
X_18392_ net213 _01920_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15626__428 clknet_1_0__leaf__03640_ VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__inv_2
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14555_ _08794_ VGND VGND VPWR VPWR _08795_ sky130_fd_sc_hd__buf_2
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _06632_ net2275 _07501_ VGND VGND VPWR VPWR _07509_ sky130_fd_sc_hd__mux2_1
X_18571__28 VGND VGND VPWR VPWR _18571__28/HI net28 sky130_fd_sc_hd__conb_1
X_17274_ CPU.registerFile\[20\]\[31\] CPU.registerFile\[21\]\[31\] _03737_ VGND VGND
+ VPWR VPWR _04970_ sky130_fd_sc_hd__mux2_1
X_10718_ net1976 _06145_ _06827_ VGND VGND VPWR VPWR _06832_ sky130_fd_sc_hd__mux2_1
X_14486_ CPU.registerFile\[24\]\[4\] _08686_ _08727_ _08550_ VGND VGND VPWR VPWR _08728_
+ sky130_fd_sc_hd__o211a_1
X_11698_ net2261 _07347_ _07464_ VGND VGND VPWR VPWR _07472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19013_ clknet_leaf_12_clk _02533_ VGND VGND VPWR VPWR CPU.aluIn1\[30\] sky130_fd_sc_hd__dfxtp_1
X_16225_ _03943_ _03944_ _03946_ _03730_ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__a211o_1
XFILLER_0_125_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13437_ _08400_ VGND VGND VPWR VPWR _08401_ sky130_fd_sc_hd__buf_4
XFILLER_0_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10649_ net2629 _06169_ _06788_ VGND VGND VPWR VPWR _06794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__08470_ _08470_ VGND VGND VPWR VPWR clknet_0__08470_ sky130_fd_sc_hd__clkbuf_16
X_16156_ _03702_ _03877_ _03879_ _03803_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_1__f__08370_ clknet_0__08370_ VGND VGND VPWR VPWR clknet_1_1__leaf__08370_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15107_ CPU.registerFile\[28\]\[19\] CPU.registerFile\[29\]\[19\] _02808_ VGND VGND
+ VPWR VPWR _03170_ sky130_fd_sc_hd__mux2_1
X_12319_ net1310 _07780_ VGND VGND VPWR VPWR _07840_ sky130_fd_sc_hd__nand2_1
X_16087_ _03758_ _03808_ _03812_ _03775_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15038_ _02728_ _03097_ _03102_ _02784_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16989_ _04579_ _04580_ CPU.registerFile\[17\]\[23\] VGND VGND VPWR VPWR _04693_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09530_ _05874_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__clkbuf_1
X_18728_ net517 _02252_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[28\] sky130_fd_sc_hd__dfxtp_1
X_09461_ _05400_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__inv_2
X_18659_ clknet_leaf_19_clk _02183_ VGND VGND VPWR VPWR CPU.rs2\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09392_ _05743_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13919__81 clknet_1_1__leaf__08476_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__inv_2
XFILLER_0_6_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__08499_ clknet_0__08499_ VGND VGND VPWR VPWR clknet_1_1__leaf__08499_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09728_ _05366_ _05359_ _05361_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09659_ CPU.PC\[21\] _05919_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__and2_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13295__797 clknet_1_1__leaf__08361_ VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__inv_2
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _08027_ VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__clkbuf_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ net1884 _07339_ _07427_ VGND VGND VPWR VPWR _07431_ sky130_fd_sc_hd__mux2_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14340_ _08568_ VGND VGND VPWR VPWR _08586_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11552_ net1723 _07339_ _07390_ VGND VGND VPWR VPWR _07394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10503_ _06715_ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__clkbuf_1
X_11483_ _06266_ VGND VGND VPWR VPWR _07351_ sky130_fd_sc_hd__buf_4
X_14271_ CPU.registerFile\[17\]\[0\] _06456_ VGND VGND VPWR VPWR _08517_ sky130_fd_sc_hd__or2_1
X_16010_ _03736_ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__buf_4
X_10434_ _06678_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__clkbuf_1
X_13222_ _08311_ _08331_ VGND VGND VPWR VPWR _08336_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10365_ _06634_ net1770 _06618_ VGND VGND VPWR VPWR _06635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13153_ CPU.cycles\[13\] CPU.cycles\[14\] _08283_ VGND VGND VPWR VPWR _08285_ sky130_fd_sc_hd__and3_1
X_12104_ net12 _07693_ _07697_ _07175_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__o211a_1
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17961_ net972 _01489_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_13084_ CPU.registerFile\[4\]\[3\] _06485_ _08239_ VGND VGND VPWR VPWR _08248_ sky130_fd_sc_hd__mux2_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605__988 clknet_1_0__leaf__08445_ VGND VGND VPWR VPWR net1044 sky130_fd_sc_hd__inv_2
X_10296_ _06588_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__clkbuf_1
X_12035_ _07651_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__clkbuf_1
X_16912_ CPU.registerFile\[19\]\[21\] CPU.registerFile\[18\]\[21\] _04327_ VGND VGND
+ VPWR VPWR _04618_ sky130_fd_sc_hd__mux2_1
X_17892_ clknet_leaf_26_clk _01420_ VGND VGND VPWR VPWR CPU.mem_wmask\[2\] sky130_fd_sc_hd__dfxtp_1
X_17419__41 clknet_1_0__leaf__05014_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__inv_2
X_16843_ _03704_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__buf_4
X_16774_ CPU.registerFile\[27\]\[18\] CPU.registerFile\[26\]\[18\] _04242_ VGND VGND
+ VPWR VPWR _04483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13986_ clknet_1_1__leaf__08473_ VGND VGND VPWR VPWR _08483_ sky130_fd_sc_hd__buf_1
X_18513_ net334 _02037_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12937_ _08170_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__clkbuf_1
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18444_ net265 _01972_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _06337_ net2468 _08131_ VGND VGND VPWR VPWR _08134_ sky130_fd_sc_hd__mux2_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13354__850 clknet_1_0__leaf__08367_ VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__inv_2
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14607_ _08844_ _08845_ _08609_ VGND VGND VPWR VPWR _08846_ sky130_fd_sc_hd__mux2_1
X_11819_ _07536_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__clkbuf_1
X_18375_ net196 _01903_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15587_ net2451 _03566_ _03637_ _03390_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _06655_ net2561 _08087_ VGND VGND VPWR VPWR _08096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14538_ _08520_ _08775_ _08778_ _08661_ VGND VGND VPWR VPWR _08779_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17257_ CPU.registerFile\[5\]\[31\] CPU.registerFile\[4\]\[31\] _03697_ VGND VGND
+ VPWR VPWR _04953_ sky130_fd_sc_hd__mux2_1
X_14469_ _08425_ _08691_ _08711_ _08597_ VGND VGND VPWR VPWR _08712_ sky130_fd_sc_hd__a211o_1
X_17320__733 clknet_1_0__leaf__04982_ VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__inv_2
XFILLER_0_70_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16208_ net2658 _03566_ _03930_ _03855_ VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17188_ _03748_ _03750_ CPU.registerFile\[1\]\[29\] VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__a21o_1
XFILLER_0_141_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__08453_ _08453_ VGND VGND VPWR VPWR clknet_0__08453_ sky130_fd_sc_hd__clkbuf_16
X_16139_ _03703_ _03860_ _03862_ _03714_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08961_ CPU.aluIn1\[11\] _05312_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__and2_1
X_08892_ _05240_ _05241_ _05243_ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__a21o_2
X_09513_ _05857_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13646__1025 clknet_1_0__leaf__08449_ VGND VGND VPWR VPWR net1081 sky130_fd_sc_hd__inv_2
XFILLER_0_91_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09444_ CPU.Bimm\[10\] _05422_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15609__412 clknet_1_1__leaf__03639_ VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__inv_2
XFILLER_0_94_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09375_ _05515_ _05692_ _05694_ _05514_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10150_ mapped_spi_ram.rcv_data\[11\] _05857_ _05762_ net1327 VGND VGND VPWR VPWR
+ _06474_ sky130_fd_sc_hd__a22o_4
XFILLER_0_112_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10081_ _06126_ _06405_ _06407_ _05818_ VGND VGND VPWR VPWR _06408_ sky130_fd_sc_hd__o211a_1
X_14232__362 clknet_1_0__leaf__08508_ VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__08511_ clknet_0__08511_ VGND VGND VPWR VPWR clknet_1_0__leaf__08511_
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f__08442_ clknet_0__08442_ VGND VGND VPWR VPWR clknet_1_0__leaf__08442_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10983_ _05614_ _07028_ _05613_ VGND VGND VPWR VPWR _07029_ sky130_fd_sc_hd__a21bo_1
X_15510_ _03230_ _03558_ _03562_ _05876_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__o211a_1
X_12722_ _08055_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16490_ _04080_ _04081_ CPU.registerFile\[25\]\[11\] VGND VGND VPWR VPWR _04206_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15441_ net1581 _03201_ _03495_ _03390_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__o211a_1
X_12653_ _06645_ net2103 _08015_ VGND VGND VPWR VPWR _08019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11604_ net2459 _07322_ _07416_ VGND VGND VPWR VPWR _07422_ sky130_fd_sc_hd__mux2_1
X_18160_ net1171 _01688_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dfxtp_1
X_15372_ CPU.registerFile\[16\]\[26\] _03159_ _03427_ _03161_ VGND VGND VPWR VPWR
+ _03428_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12584_ _07982_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17111_ _03766_ _04808_ _04810_ _03716_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__a211o_1
XFILLER_0_52_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14323_ _08568_ VGND VGND VPWR VPWR _08569_ sky130_fd_sc_hd__buf_4
X_18091_ net1102 _01619_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_11535_ net1815 _07322_ _07379_ VGND VGND VPWR VPWR _07385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17042_ _04742_ _04743_ _04557_ VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11466_ net1794 _07339_ _07333_ VGND VGND VPWR VPWR _07340_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__03680_ clknet_0__03680_ VGND VGND VPWR VPWR clknet_1_1__leaf__03680_
+ sky130_fd_sc_hd__clkbuf_16
X_15738__529 clknet_1_1__leaf__03651_ VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__inv_2
X_13205_ _06184_ _06213_ _06130_ VGND VGND VPWR VPWR _08319_ sky130_fd_sc_hd__a21o_1
X_10417_ _06669_ VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__clkbuf_1
X_11397_ _07273_ VGND VGND VPWR VPWR _07296_ sky130_fd_sc_hd__buf_4
XFILLER_0_110_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13136_ net1568 _08273_ VGND VGND VPWR VPWR _08276_ sky130_fd_sc_hd__nor2_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _06623_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__clkbuf_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18993_ clknet_leaf_14_clk _02513_ VGND VGND VPWR VPWR CPU.aluIn1\[10\] sky130_fd_sc_hd__dfxtp_2
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _08216_ VGND VGND VPWR VPWR _08239_ sky130_fd_sc_hd__buf_4
X_17944_ net955 _01472_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_10279_ _06579_ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__clkbuf_1
X_13706__1079 clknet_1_0__leaf__08455_ VGND VGND VPWR VPWR net1135 sky130_fd_sc_hd__inv_2
X_12018_ _07642_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__clkbuf_1
X_17875_ clknet_leaf_24_clk _00024_ VGND VGND VPWR VPWR CPU.cycles\[18\] sky130_fd_sc_hd__dfxtp_1
X_16826_ CPU.registerFile\[22\]\[19\] CPU.registerFile\[23\]\[19\] _04362_ VGND VGND
+ VPWR VPWR _04534_ sky130_fd_sc_hd__mux2_1
X_16757_ CPU.registerFile\[12\]\[18\] _04421_ _04422_ _04465_ VGND VGND VPWR VPWR
+ _04466_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15708_ clknet_1_1__leaf__03643_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__buf_1
X_14209__342 clknet_1_0__leaf__08505_ VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__inv_2
X_16688_ CPU.registerFile\[27\]\[16\] CPU.registerFile\[26\]\[16\] _04242_ VGND VGND
+ VPWR VPWR _04399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18427_ net248 _01955_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_09160_ _05413_ _05510_ _05511_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18358_ net179 _01886_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09091_ _05442_ _05269_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__nor2_2
X_18289_ net110 _01817_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold901 CPU.registerFile\[7\]\[31\] VGND VGND VPWR VPWR net2198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__08505_ _08505_ VGND VGND VPWR VPWR clknet_0__08505_ sky130_fd_sc_hd__clkbuf_16
Xhold912 CPU.registerFile\[22\]\[28\] VGND VGND VPWR VPWR net2209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 CPU.registerFile\[16\]\[16\] VGND VGND VPWR VPWR net2220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold934 CPU.registerFile\[30\]\[11\] VGND VGND VPWR VPWR net2231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 CPU.registerFile\[16\]\[5\] VGND VGND VPWR VPWR net2242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__08436_ _08436_ VGND VGND VPWR VPWR clknet_0__08436_ sky130_fd_sc_hd__clkbuf_16
Xhold956 CPU.registerFile\[31\]\[15\] VGND VGND VPWR VPWR net2253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 CPU.registerFile\[29\]\[3\] VGND VGND VPWR VPWR net2264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 CPU.registerFile\[21\]\[14\] VGND VGND VPWR VPWR net2275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 CPU.registerFile\[12\]\[7\] VGND VGND VPWR VPWR net2286 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ _06126_ _06322_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08367_ _08367_ VGND VGND VPWR VPWR clknet_0__08367_ sky130_fd_sc_hd__clkbuf_16
X_08944_ _05294_ _05295_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__or2_2
XFILLER_0_149_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09427_ _05255_ _05256_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09358_ CPU.PC\[1\] _05709_ _05643_ VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13941__101 clknet_1_0__leaf__08478_ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__inv_2
XFILLER_0_151_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09289_ _05558_ _05639_ _05640_ _05235_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__o211a_1
X_11320_ _07255_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11251_ _07218_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10202_ _06126_ _06520_ _06523_ _05818_ VGND VGND VPWR VPWR _06524_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11182_ _07163_ VGND VGND VPWR VPWR _07175_ sky130_fd_sc_hd__clkbuf_4
X_10133_ _06393_ VGND VGND VPWR VPWR _06458_ sky130_fd_sc_hd__inv_2
X_15990_ _06171_ VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__clkbuf_8
X_14941_ _08808_ _08809_ CPU.registerFile\[25\]\[15\] VGND VGND VPWR VPWR _03008_
+ sky130_fd_sc_hd__a21o_1
X_10064_ _05520_ _05709_ VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__nand2_2
X_17660_ per_uart.uart0.rx_bitcount\[0\] _05194_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__and2_1
X_14872_ CPU.registerFile\[8\]\[13\] _08776_ _02940_ _02864_ VGND VGND VPWR VPWR _02941_
+ sky130_fd_sc_hd__o211a_1
X_16611_ CPU.registerFile\[22\]\[14\] CPU.registerFile\[23\]\[14\] _03958_ VGND VGND
+ VPWR VPWR _04324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17591_ _05122_ per_uart.uart0.tx_bitcount\[0\] _05147_ _05150_ VGND VGND VPWR VPWR
+ _02670_ sky130_fd_sc_hd__a31o_1
X_16542_ _04247_ _04256_ _04138_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14083__229 clknet_1_0__leaf__08492_ VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__inv_2
XFILLER_0_97_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10966_ _07008_ _07015_ VGND VGND VPWR VPWR _07016_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12705_ _08046_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__clkbuf_1
X_16473_ CPU.registerFile\[13\]\[11\] _03976_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10897_ net2647 _06962_ _06868_ VGND VGND VPWR VPWR _06963_ sky130_fd_sc_hd__mux2_1
X_18212_ net1223 _01740_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[13\] sky130_fd_sc_hd__dfxtp_1
X_15424_ CPU.registerFile\[13\]\[27\] CPU.registerFile\[12\]\[27\] _08794_ VGND VGND
+ VPWR VPWR _03479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12636_ _06628_ net2235 _08004_ VGND VGND VPWR VPWR _08010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19192_ clknet_leaf_3_clk _02710_ VGND VGND VPWR VPWR per_uart.d_in_uart\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18143_ net1154 _01671_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15355_ _03138_ _03139_ CPU.registerFile\[9\]\[25\] VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12567_ _07973_ VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14306_ _08418_ VGND VGND VPWR VPWR _08552_ sky130_fd_sc_hd__clkbuf_4
X_18074_ net1085 _01602_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_11518_ net1745 _07374_ _07311_ VGND VGND VPWR VPWR _07375_ sky130_fd_sc_hd__mux2_1
X_15286_ CPU.registerFile\[6\]\[23\] CPU.registerFile\[7\]\[23\] _02982_ VGND VGND
+ VPWR VPWR _03345_ sky130_fd_sc_hd__mux2_1
X_12498_ _07936_ VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold208 mapped_spi_flash.cmd_addr\[7\] VGND VGND VPWR VPWR net1505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 mapped_spi_ram.rcv_data\[21\] VGND VGND VPWR VPWR net1516 sky130_fd_sc_hd__dlygate4sd3_1
X_17025_ _04579_ _04580_ CPU.registerFile\[17\]\[24\] VGND VGND VPWR VPWR _04728_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11449_ _06009_ VGND VGND VPWR VPWR _07328_ sky130_fd_sc_hd__buf_4
X_13645__1024 clknet_1_0__leaf__08449_ VGND VGND VPWR VPWR net1080 sky130_fd_sc_hd__inv_2
XFILLER_0_22_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _05237_ _07023_ _08266_ VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__nor3_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18976_ net750 _02496_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ net938 _01455_ VGND VGND VPWR VPWR CPU.aluShamt\[2\] sky130_fd_sc_hd__dfxtp_1
X_17858_ clknet_leaf_22_clk _00026_ VGND VGND VPWR VPWR CPU.cycles\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16809_ _04515_ _04516_ _04153_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__mux2_1
X_17789_ net869 _01351_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15684__480 clknet_1_1__leaf__03646_ VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__inv_2
XFILLER_0_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09212_ CPU.aluIn1\[18\] _05543_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09143_ _05371_ CPU.aluIn1\[23\] VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04979_ clknet_0__04979_ VGND VGND VPWR VPWR clknet_1_1__leaf__04979_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09074_ _05420_ _05253_ _05415_ _05425_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__o31a_1
XFILLER_0_31_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold720 CPU.registerFile\[17\]\[12\] VGND VGND VPWR VPWR net2017 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 CPU.registerFile\[7\]\[4\] VGND VGND VPWR VPWR net2028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 CPU.registerFile\[30\]\[0\] VGND VGND VPWR VPWR net2039 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold753 CPU.registerFile\[28\]\[16\] VGND VGND VPWR VPWR net2050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 CPU.registerFile\[5\]\[28\] VGND VGND VPWR VPWR net2061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 CPU.registerFile\[16\]\[23\] VGND VGND VPWR VPWR net2072 sky130_fd_sc_hd__dlygate4sd3_1
X_13889__53 clknet_1_0__leaf__08474_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__inv_2
X_13521__912 clknet_1_1__leaf__08437_ VGND VGND VPWR VPWR net968 sky130_fd_sc_hd__inv_2
Xhold786 CPU.registerFile\[16\]\[25\] VGND VGND VPWR VPWR net2083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 CPU.registerFile\[7\]\[23\] VGND VGND VPWR VPWR net2094 sky130_fd_sc_hd__dlygate4sd3_1
X_09976_ CPU.PC\[9\] _05885_ CPU.PC\[10\] VGND VGND VPWR VPWR _06307_ sky130_fd_sc_hd__a21oi_1
X_08927_ CPU.aluIn1\[1\] VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__inv_2
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03683_ clknet_0__03683_ VGND VGND VPWR VPWR clknet_1_0__leaf__03683_
+ sky130_fd_sc_hd__clkbuf_16
X_10820_ CPU.aluIn1\[21\] _06903_ _06881_ VGND VGND VPWR VPWR _06904_ sky130_fd_sc_hd__mux2_1
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10751_ net2537 _06530_ _06815_ VGND VGND VPWR VPWR _06849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13470_ _08426_ VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__clkbuf_1
X_10682_ net2572 _06555_ _06776_ VGND VGND VPWR VPWR _06811_ sky130_fd_sc_hd__mux2_1
X_13705__1078 clknet_1_0__leaf__08455_ VGND VGND VPWR VPWR net1134 sky130_fd_sc_hd__inv_2
X_12421_ net1874 _07332_ _07895_ VGND VGND VPWR VPWR _07896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15140_ _05876_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__clkbuf_4
X_12352_ _07847_ VGND VGND VPWR VPWR _07859_ sky130_fd_sc_hd__buf_4
XFILLER_0_90_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11303_ _07246_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__clkbuf_1
X_15071_ CPU.registerFile\[13\]\[18\] CPU.registerFile\[12\]\[18\] _02935_ VGND VGND
+ VPWR VPWR _03135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12283_ net1465 _07812_ _07816_ _07809_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11234_ _07209_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__clkbuf_1
X_18830_ net619 _02354_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_11165_ mapped_spi_flash.rcv_data\[8\] _07134_ VGND VGND VPWR VPWR _07166_ sky130_fd_sc_hd__or2_1
X_10116_ _06441_ VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__clkbuf_1
X_15973_ CPU.registerFile\[8\]\[0\] _08394_ _06150_ _03699_ VGND VGND VPWR VPWR _03700_
+ sky130_fd_sc_hd__o211a_1
X_11096_ _07119_ _07122_ _07120_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__o21ba_1
X_18761_ net550 _02285_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[23\] sky130_fd_sc_hd__dfxtp_1
X_14924_ _02750_ _02973_ _02991_ _02839_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__a211o_1
X_17712_ _05232_ VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__clkbuf_1
X_10047_ _05296_ _06374_ VGND VGND VPWR VPWR _06375_ sky130_fd_sc_hd__xnor2_2
X_18692_ net481 _02216_ VGND VGND VPWR VPWR mapped_spi_flash.clk_div sky130_fd_sc_hd__dfxtp_1
Xhold80 _06412_ VGND VGND VPWR VPWR net1377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 _06244_ VGND VGND VPWR VPWR net1388 sky130_fd_sc_hd__dlygate4sd3_1
X_14855_ CPU.registerFile\[30\]\[13\] CPU.registerFile\[31\]\[13\] _02887_ VGND VGND
+ VPWR VPWR _02924_ sky130_fd_sc_hd__mux2_1
X_17643_ _04989_ _04990_ _05182_ per_uart.uart0.uart_rxd2 VGND VGND VPWR VPWR _05183_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_86_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13948__107 clknet_1_0__leaf__08479_ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__inv_2
X_17574_ _03659_ _05136_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__nor2_1
X_14786_ _08722_ _02852_ _02856_ _08851_ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__o211a_1
X_11998_ _06659_ net2432 _07597_ VGND VGND VPWR VPWR _07631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16525_ CPU.registerFile\[28\]\[12\] CPU.registerFile\[29\]\[12\] _04122_ VGND VGND
+ VPWR VPWR _04240_ sky130_fd_sc_hd__mux2_1
X_10949_ mapped_spi_flash.cmd_addr\[23\] _06983_ _06985_ mapped_spi_flash.cmd_addr\[22\]
+ VGND VGND VPWR VPWR _07003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__08339_ clknet_0__08339_ VGND VGND VPWR VPWR clknet_1_0__leaf__08339_
+ sky130_fd_sc_hd__clkbuf_16
X_16456_ _04171_ _04172_ _03961_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15407_ CPU.registerFile\[17\]\[27\] _08528_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__or2_1
X_19175_ clknet_leaf_6_clk _02695_ VGND VGND VPWR VPWR per_uart.uart0.rx_bitcount\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12619_ _06611_ net2251 _07993_ VGND VGND VPWR VPWR _08001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16387_ _08400_ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_109_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15896__639 clknet_1_0__leaf__03684_ VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__inv_2
XFILLER_0_42_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18126_ net1137 _01654_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15338_ CPU.registerFile\[22\]\[25\] CPU.registerFile\[23\]\[25\] _08584_ VGND VGND
+ VPWR VPWR _03395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18057_ net1068 _01585_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_15269_ CPU.registerFile\[30\]\[23\] CPU.registerFile\[31\]\[23\] _03291_ VGND VGND
+ VPWR VPWR _03328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17008_ _04389_ _04390_ CPU.registerFile\[1\]\[24\] VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03646_ clknet_0__03646_ VGND VGND VPWR VPWR clknet_1_1__leaf__03646_
+ sky130_fd_sc_hd__clkbuf_16
X_13994__149 clknet_1_1__leaf__08483_ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__inv_2
XFILLER_0_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09830_ CPU.Jimm\[16\] _05758_ _05790_ CPU.cycles\[16\] _06166_ VGND VGND VPWR VPWR
+ _06167_ sky130_fd_sc_hd__a221o_1
XFILLER_0_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _05881_ _06088_ _06100_ _05540_ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__a2bb2o_1
X_18959_ net733 _02479_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ mapped_spi_ram.rcv_data\[13\] _05685_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18577__34 VGND VGND VPWR VPWR _18577__34/HI net34 sky130_fd_sc_hd__conb_1
X_14066__213 clknet_1_0__leaf__08491_ VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__inv_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09126_ _05351_ _05343_ _05477_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09057_ CPU.aluIn1\[28\] _05257_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold550 CPU.registerFile\[15\]\[20\] VGND VGND VPWR VPWR net1847 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold561 CPU.registerFile\[15\]\[15\] VGND VGND VPWR VPWR net1858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 CPU.registerFile\[11\]\[28\] VGND VGND VPWR VPWR net1869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 CPU.registerFile\[18\]\[3\] VGND VGND VPWR VPWR net1880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 CPU.registerFile\[3\]\[28\] VGND VGND VPWR VPWR net1891 sky130_fd_sc_hd__dlygate4sd3_1
X_09959_ _05745_ _06280_ _06286_ _06290_ VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__a211o_2
X_13302__803 clknet_1_0__leaf__08362_ VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__inv_2
X_12970_ net2207 _07324_ _08181_ VGND VGND VPWR VPWR _08188_ sky130_fd_sc_hd__mux2_1
Xhold1250 CPU.registerFile\[8\]\[31\] VGND VGND VPWR VPWR net2547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 CPU.registerFile\[25\]\[30\] VGND VGND VPWR VPWR net2558 sky130_fd_sc_hd__dlygate4sd3_1
X_11921_ _07590_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__clkbuf_1
Xhold1272 CPU.registerFile\[23\]\[11\] VGND VGND VPWR VPWR net2569 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1283 CPU.registerFile\[1\]\[26\] VGND VGND VPWR VPWR net2580 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1294 CPU.aluIn1\[25\] VGND VGND VPWR VPWR net2591 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _08415_ _08875_ _08877_ _08420_ VGND VGND VPWR VPWR _08878_ sky130_fd_sc_hd__a211o_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ net1852 _07364_ _07548_ VGND VGND VPWR VPWR _07554_ sky130_fd_sc_hd__mux2_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13259__779 clknet_1_0__leaf__08344_ VGND VGND VPWR VPWR net835 sky130_fd_sc_hd__inv_2
X_13644__1023 clknet_1_0__leaf__08449_ VGND VGND VPWR VPWR net1079 sky130_fd_sc_hd__inv_2
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10803_ CPU.aluReg\[26\] CPU.aluReg\[24\] _06872_ VGND VGND VPWR VPWR _06891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ CPU.registerFile\[24\]\[6\] _08686_ _08810_ _08550_ VGND VGND VPWR VPWR _08811_
+ sky130_fd_sc_hd__o211a_1
X_13491__885 clknet_1_0__leaf__08434_ VGND VGND VPWR VPWR net941 sky130_fd_sc_hd__inv_2
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _07517_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__clkbuf_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16310_ CPU.registerFile\[0\]\[7\] _03828_ _03725_ _04029_ VGND VGND VPWR VPWR _04030_
+ sky130_fd_sc_hd__o211a_1
X_10734_ _06840_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16241_ _03765_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13453_ _08413_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__clkbuf_1
X_10665_ _06802_ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15821__571 clknet_1_0__leaf__03656_ VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__inv_2
X_12404_ net1715 _07316_ _07884_ VGND VGND VPWR VPWR _07887_ sky130_fd_sc_hd__mux2_1
X_16172_ CPU.registerFile\[8\]\[4\] _08394_ _06150_ _03894_ VGND VGND VPWR VPWR _03895_
+ sky130_fd_sc_hd__o211a_1
X_10596_ net1977 _06361_ _06761_ VGND VGND VPWR VPWR _06765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15123_ CPU.registerFile\[8\]\[19\] _03018_ _03185_ _02864_ VGND VGND VPWR VPWR _03186_
+ sky130_fd_sc_hd__o211a_1
X_12335_ _07850_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15054_ CPU.registerFile\[16\]\[18\] _02755_ _03117_ _02757_ VGND VGND VPWR VPWR
+ _03118_ sky130_fd_sc_hd__o211a_1
X_12266_ net1536 _07799_ _07806_ _07796_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__o211a_1
X_11217_ _06663_ _07199_ VGND VGND VPWR VPWR _07200_ sky130_fd_sc_hd__nand2_4
X_12197_ mapped_spi_ram.snd_bitcount\[4\] _07758_ VGND VGND VPWR VPWR _07759_ sky130_fd_sc_hd__or2_1
X_18813_ net602 _02337_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_11148_ _05721_ _07132_ VGND VGND VPWR VPWR _07156_ sky130_fd_sc_hd__nand2_1
X_18744_ net533 _02268_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[6\] sky130_fd_sc_hd__dfxtp_1
X_14015__167 clknet_1_0__leaf__08486_ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__inv_2
X_11079_ _07108_ _07109_ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__nor2_1
X_14907_ CPU.registerFile\[13\]\[14\] CPU.registerFile\[12\]\[14\] _02935_ VGND VGND
+ VPWR VPWR _02975_ sky130_fd_sc_hd__mux2_1
X_18675_ net464 _02199_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17626_ per_uart.rx_data\[2\] net1670 _05170_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__mux2_1
X_14838_ _02906_ _02907_ _08783_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14769_ net1577 _02797_ _02840_ _08751_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__o211a_1
X_17557_ _05121_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15904__646 clknet_1_0__leaf__03685_ VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__inv_2
X_16508_ CPU.registerFile\[8\]\[12\] _04101_ _04102_ _04222_ VGND VGND VPWR VPWR _04223_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17488_ _05022_ _06255_ _08256_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16439_ _03985_ _03986_ CPU.registerFile\[1\]\[10\] VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15603__407 clknet_1_0__leaf__03638_ VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__inv_2
XFILLER_0_42_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19158_ clknet_leaf_5_clk net1511 VGND VGND VPWR VPWR per_uart.uart0.txd_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18109_ net1120 _01637_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19089_ net72 _02609_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09813_ _06149_ VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__buf_4
X_13704__1077 clknet_1_0__leaf__08455_ VGND VGND VPWR VPWR net1133 sky130_fd_sc_hd__inv_2
X_09744_ _06084_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__clkbuf_1
X_09675_ _05379_ _05899_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15879__623 clknet_1_1__leaf__03683_ VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__inv_2
XFILLER_0_80_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10450_ _06686_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09109_ _05264_ CPU.aluIn1\[9\] VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__or2b_1
X_10381_ _06645_ net2091 _06639_ VGND VGND VPWR VPWR _06646_ sky130_fd_sc_hd__mux2_1
X_12120_ mapped_spi_ram.cmd_addr\[23\] _07704_ _07706_ VGND VGND VPWR VPWR _07707_
+ sky130_fd_sc_hd__o21ba_1
X_13977__133 clknet_1_0__leaf__08482_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__inv_2
XFILLER_0_32_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12051_ CPU.registerFile\[24\]\[9\] _07358_ _07657_ VGND VGND VPWR VPWR _07660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold380 CPU.registerFile\[3\]\[1\] VGND VGND VPWR VPWR net1677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 CPU.registerFile\[19\]\[4\] VGND VGND VPWR VPWR net1688 sky130_fd_sc_hd__dlygate4sd3_1
X_11002_ mapped_spi_flash.cmd_addr\[12\] _07045_ _07039_ VGND VGND VPWR VPWR _07046_
+ sky130_fd_sc_hd__mux2_1
X_15810_ _08356_ _03673_ _03661_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__a21oi_1
X_16790_ _04489_ _04498_ _04138_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__o21a_1
X_15741_ clknet_1_1__leaf__03643_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__buf_1
X_12953_ _08178_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__clkbuf_1
Xhold1080 CPU.registerFile\[31\]\[30\] VGND VGND VPWR VPWR net2377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 CPU.PC\[5\] VGND VGND VPWR VPWR net2388 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ _07581_ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18460_ net281 _01988_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_12884_ _06530_ net2230 _08108_ VGND VGND VPWR VPWR _08142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _08557_ _08856_ _08861_ _08423_ VGND VGND VPWR VPWR _08862_ sky130_fd_sc_hd__o211a_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11835_ net2476 _07347_ _07537_ VGND VGND VPWR VPWR _07545_ sky130_fd_sc_hd__mux2_1
X_18391_ net212 _01919_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_25_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03649_ clknet_0__03649_ VGND VGND VPWR VPWR clknet_1_0__leaf__03649_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _06061_ VGND VGND VPWR VPWR _08794_ sky130_fd_sc_hd__clkbuf_8
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _07508_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14203__337 clknet_1_0__leaf__08504_ VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__inv_2
X_17273_ CPU.registerFile\[22\]\[31\] CPU.registerFile\[23\]\[31\] _03761_ VGND VGND
+ VPWR VPWR _04969_ sky130_fd_sc_hd__mux2_1
X_10717_ _06831_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__clkbuf_1
X_14485_ _08546_ _08547_ CPU.registerFile\[25\]\[4\] VGND VGND VPWR VPWR _08727_ sky130_fd_sc_hd__a21o_1
X_11697_ _07471_ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16224_ CPU.registerFile\[0\]\[5\] _03828_ _03725_ _03945_ VGND VGND VPWR VPWR _03946_
+ sky130_fd_sc_hd__o211a_1
X_19012_ clknet_leaf_12_clk _02532_ VGND VGND VPWR VPWR CPU.aluIn1\[29\] sky130_fd_sc_hd__dfxtp_1
X_13436_ _06141_ VGND VGND VPWR VPWR _08400_ sky130_fd_sc_hd__clkbuf_8
X_10648_ _06793_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16155_ CPU.registerFile\[24\]\[3\] _08393_ _03747_ _03878_ VGND VGND VPWR VPWR _03879_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13367_ clknet_1_1__leaf__08366_ VGND VGND VPWR VPWR _08369_ sky130_fd_sc_hd__buf_1
XFILLER_0_106_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10579_ net1870 _06169_ _06750_ VGND VGND VPWR VPWR _06756_ sky130_fd_sc_hd__mux2_1
X_15106_ CPU.registerFile\[30\]\[19\] CPU.registerFile\[31\]\[19\] _02887_ VGND VGND
+ VPWR VPWR _03169_ sky130_fd_sc_hd__mux2_1
X_12318_ net1306 _07837_ _07838_ _07839_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__a22o_1
X_16086_ _03766_ _03809_ _03811_ _06142_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15037_ _03098_ _03099_ _03101_ _02903_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__a211o_1
X_12249_ mapped_spi_ram.rcv_data\[23\] _07787_ VGND VGND VPWR VPWR _07797_ sky130_fd_sc_hd__or2_1
X_16988_ CPU.registerFile\[19\]\[23\] CPU.registerFile\[18\]\[23\] _04327_ VGND VGND
+ VPWR VPWR _04692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18727_ net516 _02251_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[27\] sky130_fd_sc_hd__dfxtp_1
Xwire14 _07690_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__05015_ clknet_0__05015_ VGND VGND VPWR VPWR clknet_1_1__leaf__05015_
+ sky130_fd_sc_hd__clkbuf_16
X_09460_ _05381_ _05382_ _05391_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_64_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18658_ clknet_leaf_18_clk _02182_ VGND VGND VPWR VPWR CPU.rs2\[30\] sky130_fd_sc_hd__dfxtp_1
X_15828__577 clknet_1_0__leaf__03678_ VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__inv_2
X_17609_ net1474 _05159_ _05162_ _07108_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__o22a_1
X_09391_ net2276 _05734_ _05742_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18589_ net410 net46 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[25\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_16_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14178__314 clknet_1_0__leaf__08502_ VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__inv_2
XFILLER_0_117_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08498_ clknet_0__08498_ VGND VGND VPWR VPWR clknet_1_1__leaf__08498_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_112_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13643__1022 clknet_1_0__leaf__08449_ VGND VGND VPWR VPWR net1078 sky130_fd_sc_hd__inv_2
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09727_ _05366_ _05486_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__xor2_1
X_13557__944 clknet_1_1__leaf__08441_ VGND VGND VPWR VPWR net1000 sky130_fd_sc_hd__inv_2
XFILLER_0_69_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09658_ _05925_ _05995_ _05999_ _06001_ _05998_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__a32o_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _05931_ _05932_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _07430_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__clkbuf_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11551_ _07393_ VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10502_ net1873 _06083_ _06713_ VGND VGND VPWR VPWR _06715_ sky130_fd_sc_hd__mux2_1
X_14044__193 clknet_1_1__leaf__08489_ VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__inv_2
X_14270_ CPU.registerFile\[19\]\[0\] CPU.registerFile\[18\]\[0\] _06064_ VGND VGND
+ VPWR VPWR _08516_ sky130_fd_sc_hd__mux2_1
X_11482_ _07350_ VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13221_ _08334_ VGND VGND VPWR VPWR _08335_ sky130_fd_sc_hd__clkbuf_4
X_10433_ _06620_ net2523 _06676_ VGND VGND VPWR VPWR _06678_ sky130_fd_sc_hd__mux2_1
X_13819__1181 clknet_1_0__leaf__08466_ VGND VGND VPWR VPWR net1237 sky130_fd_sc_hd__inv_2
XFILLER_0_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13152_ net1621 _08283_ VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__xor2_1
X_10364_ _06244_ VGND VGND VPWR VPWR _06634_ sky130_fd_sc_hd__buf_4
XFILLER_0_103_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12103_ net1365 _07694_ _07696_ VGND VGND VPWR VPWR _07697_ sky130_fd_sc_hd__a21o_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ net1392 VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__clkbuf_1
X_17960_ net971 _01488_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_10295_ net1688 _06465_ _06580_ VGND VGND VPWR VPWR _06588_ sky130_fd_sc_hd__mux2_1
X_12034_ CPU.registerFile\[24\]\[17\] _07341_ _07646_ VGND VGND VPWR VPWR _07651_
+ sky130_fd_sc_hd__mux2_1
X_16911_ _04615_ _04616_ _04365_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__mux2_1
X_17891_ clknet_leaf_26_clk _01419_ VGND VGND VPWR VPWR CPU.mem_wmask\[1\] sky130_fd_sc_hd__dfxtp_1
X_16842_ _04503_ _04546_ _04548_ _04509_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__a211o_1
X_15632__433 clknet_1_0__leaf__03641_ VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__inv_2
X_13497__891 clknet_1_0__leaf__08434_ VGND VGND VPWR VPWR net947 sky130_fd_sc_hd__inv_2
X_16773_ _04480_ _04481_ _04279_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__mux2_1
X_18512_ net333 _02036_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12936_ _06337_ net1612 _08167_ VGND VGND VPWR VPWR _08170_ sky130_fd_sc_hd__mux2_1
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18443_ net264 _01971_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ _08133_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ net2260 _07330_ _07526_ VGND VGND VPWR VPWR _07536_ sky130_fd_sc_hd__mux2_1
X_14606_ CPU.registerFile\[28\]\[7\] CPU.registerFile\[29\]\[7\] _08538_ VGND VGND
+ VPWR VPWR _08845_ sky130_fd_sc_hd__mux2_1
X_14127__268 clknet_1_0__leaf__08497_ VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__inv_2
X_15586_ _06339_ _03619_ _03636_ _03601_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__a211o_1
X_18374_ net195 _01902_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ _08095_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ CPU.registerFile\[8\]\[5\] _08776_ _08777_ _08622_ VGND VGND VPWR VPWR _08778_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11749_ _07499_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_839 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17256_ CPU.registerFile\[6\]\[31\] CPU.registerFile\[7\]\[31\] _03847_ VGND VGND
+ VPWR VPWR _04952_ sky130_fd_sc_hd__mux2_1
X_13703__1076 clknet_1_1__leaf__08455_ VGND VGND VPWR VPWR net1132 sky130_fd_sc_hd__inv_2
X_14468_ _08701_ _08710_ _08594_ VGND VGND VPWR VPWR _08711_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13419_ _05739_ _06287_ _08388_ VGND VGND VPWR VPWR _08389_ sky130_fd_sc_hd__mux2_1
X_16207_ _03692_ _03910_ _03929_ _03601_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__a211o_1
X_17187_ CPU.registerFile\[2\]\[29\] CPU.registerFile\[3\]\[29\] _03759_ VGND VGND
+ VPWR VPWR _04885_ sky130_fd_sc_hd__mux2_1
X_14399_ CPU.registerFile\[20\]\[2\] _08527_ _08642_ _08530_ VGND VGND VPWR VPWR _08643_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16138_ CPU.registerFile\[12\]\[3\] _03707_ _03708_ _03861_ VGND VGND VPWR VPWR _03862_
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_0__08452_ _08452_ VGND VGND VPWR VPWR clknet_0__08452_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16069_ _08404_ _03782_ _03786_ _03794_ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__a31o_2
X_08960_ CPU.rs2\[11\] _05245_ _05249_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_5_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_16
X_15715__508 clknet_1_1__leaf__03649_ VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__inv_2
X_08891_ _05242_ VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09512_ _05761_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__clkbuf_4
X_09443_ _05409_ _05528_ _05535_ CPU.aluReg\[28\] _05791_ VGND VGND VPWR VPWR _05792_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09374_ _05693_ _05699_ _05720_ _05725_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__a31o_1
XFILLER_0_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17295__711 clknet_1_0__leaf__04979_ VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__inv_2
XFILLER_0_43_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10080_ _06126_ _06406_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__nand2_1
Xclkbuf_1_0__f__08510_ clknet_0__08510_ VGND VGND VPWR VPWR clknet_1_0__leaf__08510_
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f__08441_ clknet_0__08441_ VGND VGND VPWR VPWR clknet_1_0__leaf__08441_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10982_ _07024_ _05609_ _07026_ _07027_ VGND VGND VPWR VPWR _07028_ sky130_fd_sc_hd__a31o_1
X_12721_ _06645_ net2639 _08051_ VGND VGND VPWR VPWR _08055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15440_ _03155_ _03477_ _03494_ _03243_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__a211o_2
X_12652_ _08018_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11603_ _07421_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__clkbuf_1
X_15371_ CPU.registerFile\[17\]\[26\] _08528_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12583_ net2106 _07358_ _07979_ VGND VGND VPWR VPWR _07982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13611__993 clknet_1_0__leaf__08446_ VGND VGND VPWR VPWR net1049 sky130_fd_sc_hd__inv_2
X_17110_ CPU.registerFile\[12\]\[27\] _03694_ _03763_ _04809_ VGND VGND VPWR VPWR
+ _04810_ sky130_fd_sc_hd__o211a_1
X_14322_ _06059_ VGND VGND VPWR VPWR _08568_ sky130_fd_sc_hd__clkbuf_4
X_11534_ _07384_ VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__clkbuf_1
X_18090_ net1101 _01618_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17041_ CPU.registerFile\[5\]\[25\] CPU.registerFile\[4\]\[25\] _04428_ VGND VGND
+ VPWR VPWR _04743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14253_ clknet_1_1__leaf__08506_ VGND VGND VPWR VPWR _08510_ sky130_fd_sc_hd__buf_1
XFILLER_0_162_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11465_ _06123_ VGND VGND VPWR VPWR _07339_ sky130_fd_sc_hd__buf_4
XFILLER_0_150_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13204_ _06068_ _06227_ _06296_ _08317_ VGND VGND VPWR VPWR _08318_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10416_ _06603_ net2119 _06665_ VGND VGND VPWR VPWR _06669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11396_ _07295_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__clkbuf_1
X_13384__877 clknet_1_1__leaf__08370_ VGND VGND VPWR VPWR net933 sky130_fd_sc_hd__inv_2
X_13135_ CPU.cycles\[6\] _08273_ VGND VGND VPWR VPWR _08275_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10347_ _06622_ net2172 _06618_ VGND VGND VPWR VPWR _06623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18992_ clknet_leaf_13_clk _02512_ VGND VGND VPWR VPWR CPU.aluIn1\[9\] sky130_fd_sc_hd__dfxtp_2
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ net1407 VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__clkbuf_1
X_17943_ net954 _01471_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_10278_ net1749 _06267_ _06569_ VGND VGND VPWR VPWR _06579_ sky130_fd_sc_hd__mux2_1
X_12017_ net2592 _07324_ _07635_ VGND VGND VPWR VPWR _07642_ sky130_fd_sc_hd__mux2_1
X_17874_ clknet_leaf_23_clk _00023_ VGND VGND VPWR VPWR CPU.cycles\[17\] sky130_fd_sc_hd__dfxtp_1
X_16825_ _04479_ _04528_ _04532_ _04446_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__o211a_1
X_16756_ CPU.registerFile\[13\]\[18\] _04380_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__or2_1
XFILLER_0_159_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12919_ _06145_ net1628 _08156_ VGND VGND VPWR VPWR _08161_ sky130_fd_sc_hd__mux2_1
X_16687_ _04396_ _04397_ _04279_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__mux2_1
X_18426_ net247 _01954_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14060__208 clknet_1_1__leaf__08490_ VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__inv_2
XFILLER_0_29_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18357_ net178 _01885_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15569_ CPU.registerFile\[15\]\[31\] CPU.registerFile\[14\]\[31\] _08560_ VGND VGND
+ VPWR VPWR _03620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09090_ CPU.aluIn1\[3\] _05268_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__nor2_1
X_18288_ net109 _01816_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17239_ _04934_ _04935_ _03742_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__08504_ _08504_ VGND VGND VPWR VPWR clknet_0__08504_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold902 per_uart.uart0.tx_bitcount\[1\] VGND VGND VPWR VPWR net2199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold913 CPU.registerFile\[26\]\[14\] VGND VGND VPWR VPWR net2210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold924 CPU.registerFile\[23\]\[24\] VGND VGND VPWR VPWR net2221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 CPU.registerFile\[29\]\[2\] VGND VGND VPWR VPWR net2232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 CPU.registerFile\[23\]\[8\] VGND VGND VPWR VPWR net2243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 CPU.registerFile\[26\]\[18\] VGND VGND VPWR VPWR net2254 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__08435_ _08435_ VGND VGND VPWR VPWR clknet_0__08435_ sky130_fd_sc_hd__clkbuf_16
Xhold968 CPU.registerFile\[31\]\[12\] VGND VGND VPWR VPWR net2265 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ _05451_ _06321_ VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__xnor2_2
Xhold979 CPU.registerFile\[16\]\[31\] VGND VGND VPWR VPWR net2276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__08366_ _08366_ VGND VGND VPWR VPWR clknet_0__08366_ sky130_fd_sc_hd__clkbuf_16
X_08943_ CPU.aluIn1\[7\] _05293_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13818__1180 clknet_1_0__leaf__08466_ VGND VGND VPWR VPWR net1236 sky130_fd_sc_hd__inv_2
XFILLER_0_94_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09426_ CPU.aluIn1\[28\] _05257_ _05775_ VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09357_ _05696_ _05693_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09288_ CPU.PC\[20\] _05636_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11250_ _06628_ net2267 _07212_ VGND VGND VPWR VPWR _07218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10201_ _05427_ _06522_ VGND VGND VPWR VPWR _06523_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11181_ net2664 _07134_ VGND VGND VPWR VPWR _07174_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14156__294 clknet_1_0__leaf__08500_ VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__inv_2
X_10132_ _05788_ _06247_ _06203_ VGND VGND VPWR VPWR _06457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14940_ CPU.registerFile\[27\]\[15\] CPU.registerFile\[26\]\[15\] _02768_ VGND VGND
+ VPWR VPWR _03007_ sky130_fd_sc_hd__mux2_1
X_10063_ _05534_ _05691_ VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__nand2_1
X_14871_ _02733_ _02734_ CPU.registerFile\[9\]\[13\] VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__a21o_1
X_13702__1075 clknet_1_1__leaf__08455_ VGND VGND VPWR VPWR net1131 sky130_fd_sc_hd__inv_2
X_16610_ _04075_ _04317_ _04322_ _04042_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__o211a_1
X_17590_ _05122_ _05149_ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13753_ clknet_1_0__leaf__08451_ VGND VGND VPWR VPWR _08460_ sky130_fd_sc_hd__buf_1
X_16541_ _04170_ _04250_ _04255_ _04180_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10965_ mapped_spi_flash.cmd_addr\[18\] _05677_ _07009_ VGND VGND VPWR VPWR _07015_
+ sky130_fd_sc_hd__mux2_1
X_12704_ _06628_ net2577 _08040_ VGND VGND VPWR VPWR _08046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16472_ CPU.registerFile\[15\]\[11\] CPU.registerFile\[14\]\[11\] _04146_ VGND VGND
+ VPWR VPWR _04188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15744__534 clknet_1_0__leaf__03652_ VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__inv_2
XFILLER_0_39_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10896_ CPU.aluIn1\[3\] _06961_ _06880_ VGND VGND VPWR VPWR _06962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18211_ net1222 _01739_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15423_ CPU.registerFile\[15\]\[27\] CPU.registerFile\[14\]\[27\] _08560_ VGND VGND
+ VPWR VPWR _03478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12635_ _08009_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19191_ clknet_leaf_3_clk _02709_ VGND VGND VPWR VPWR per_uart.d_in_uart\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18142_ net1153 _01670_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_15354_ CPU.registerFile\[10\]\[25\] CPU.registerFile\[11\]\[25\] _03183_ VGND VGND
+ VPWR VPWR _03411_ sky130_fd_sc_hd__mux2_1
X_12566_ net2601 _07341_ _07968_ VGND VGND VPWR VPWR _07973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11517_ net1362 VGND VGND VPWR VPWR _07374_ sky130_fd_sc_hd__clkbuf_4
X_14305_ CPU.registerFile\[24\]\[0\] _08545_ _08548_ _08550_ VGND VGND VPWR VPWR _08551_
+ sky130_fd_sc_hd__o211a_1
X_15285_ _03133_ _03339_ _03343_ _03188_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__o211a_1
X_18073_ net1084 _01601_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_12497_ net2065 _07341_ _07931_ VGND VGND VPWR VPWR _07936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_831 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17024_ CPU.registerFile\[19\]\[24\] CPU.registerFile\[18\]\[24\] _03745_ VGND VGND
+ VPWR VPWR _04727_ sky130_fd_sc_hd__mux2_1
Xhold209 mapped_spi_flash.cmd_addr\[23\] VGND VGND VPWR VPWR net1506 sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ _07327_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__clkbuf_1
X_14239__369 clknet_1_1__leaf__08508_ VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__inv_2
XFILLER_0_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11379_ net1768 _06083_ _07285_ VGND VGND VPWR VPWR _07287_ sky130_fd_sc_hd__mux2_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ CPU.state\[1\] CPU.state\[0\] VGND VGND VPWR VPWR _08266_ sky130_fd_sc_hd__or2_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18975_ net749 _02495_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ net2211 _06082_ _08228_ VGND VGND VPWR VPWR _08230_ sky130_fd_sc_hd__mux2_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ net937 _01454_ VGND VGND VPWR VPWR CPU.aluShamt\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17857_ clknet_leaf_22_clk _00015_ VGND VGND VPWR VPWR CPU.cycles\[0\] sky130_fd_sc_hd__dfxtp_1
X_16808_ CPU.registerFile\[5\]\[19\] CPU.registerFile\[4\]\[19\] _04428_ VGND VGND
+ VPWR VPWR _04516_ sky130_fd_sc_hd__mux2_1
X_17788_ net868 _01350_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16739_ CPU.registerFile\[20\]\[17\] CPU.registerFile\[21\]\[17\] _04287_ VGND VGND
+ VPWR VPWR _04449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09211_ _05561_ _05562_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__nand2_1
X_18409_ net230 _01937_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09142_ _05379_ _05492_ _05493_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09073_ _05424_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15873__618 clknet_1_1__leaf__03682_ VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__inv_2
XFILLER_0_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold710 CPU.registerFile\[27\]\[6\] VGND VGND VPWR VPWR net2007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 CPU.registerFile\[20\]\[31\] VGND VGND VPWR VPWR net2018 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold732 CPU.registerFile\[18\]\[17\] VGND VGND VPWR VPWR net2029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold743 CPU.registerFile\[11\]\[1\] VGND VGND VPWR VPWR net2040 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold754 CPU.rs2\[9\] VGND VGND VPWR VPWR net2051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 CPU.registerFile\[3\]\[5\] VGND VGND VPWR VPWR net2062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 CPU.registerFile\[5\]\[13\] VGND VGND VPWR VPWR net2073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 CPU.registerFile\[3\]\[8\] VGND VGND VPWR VPWR net2084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold798 CPU.registerFile\[6\]\[21\] VGND VGND VPWR VPWR net2095 sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ _06305_ _05973_ VGND VGND VPWR VPWR _06306_ sky130_fd_sc_hd__xnor2_1
X_13971__128 clknet_1_1__leaf__08481_ VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__inv_2
X_08926_ _05240_ _05241_ CPU.mem_wdata\[1\] _05243_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__a211oi_2
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03682_ clknet_0__03682_ VGND VGND VPWR VPWR clknet_1_0__leaf__03682_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10750_ _06848_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09409_ CPU.Bimm\[10\] _05758_ _05759_ CPU.cycles\[30\] VGND VGND VPWR VPWR _05760_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10681_ _06810_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12420_ _07883_ VGND VGND VPWR VPWR _07895_ sky130_fd_sc_hd__buf_4
XFILLER_0_106_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12351_ _07858_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11302_ net2382 _05873_ _07238_ VGND VGND VPWR VPWR _07246_ sky130_fd_sc_hd__mux2_1
X_15070_ CPU.registerFile\[15\]\[18\] CPU.registerFile\[14\]\[18\] _03013_ VGND VGND
+ VPWR VPWR _03134_ sky130_fd_sc_hd__mux2_1
X_12282_ mapped_spi_ram.rcv_data\[9\] _07813_ VGND VGND VPWR VPWR _07816_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11233_ _06611_ net2108 _07201_ VGND VGND VPWR VPWR _07209_ sky130_fd_sc_hd__mux2_1
X_11164_ net1605 _07160_ _07165_ _07164_ VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__o211a_1
X_10115_ net2242 _06440_ _06293_ VGND VGND VPWR VPWR _06441_ sky130_fd_sc_hd__mux2_1
X_18760_ net549 _02284_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[22\] sky130_fd_sc_hd__dfxtp_1
X_15972_ CPU.registerFile\[9\]\[0\] _03698_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__or2_1
X_11095_ net2651 _07118_ VGND VGND VPWR VPWR _07122_ sky130_fd_sc_hd__and2_1
X_17711_ _05207_ _05231_ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__and2_1
X_14923_ _02981_ _02990_ _02837_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__o21a_2
X_10046_ _05300_ _06373_ _05298_ VGND VGND VPWR VPWR _06374_ sky130_fd_sc_hd__a21oi_1
X_18691_ net480 _02215_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[31\] sky130_fd_sc_hd__dfxtp_1
Xhold70 _06420_ VGND VGND VPWR VPWR net1367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 _08245_ VGND VGND VPWR VPWR net1378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 _08237_ VGND VGND VPWR VPWR net1389 sky130_fd_sc_hd__dlygate4sd3_1
X_17642_ _04988_ _04991_ per_uart.uart0.rx_busy VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__o21ai_1
X_14854_ _08837_ _02920_ _02922_ _08802_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__a211o_1
X_17573_ per_uart.uart0.tx_count16\[2\] per_uart.uart0.tx_count16\[1\] per_uart.uart0.tx_count16\[0\]
+ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__and3_1
X_14785_ _08764_ _02853_ _02855_ _02814_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__a211o_1
X_15668__465 clknet_1_1__leaf__03645_ VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__inv_2
X_11997_ _07630_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__clkbuf_1
X_16524_ CPU.registerFile\[30\]\[12\] CPU.registerFile\[31\]\[12\] _04201_ VGND VGND
+ VPWR VPWR _04239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_914 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10948_ mapped_spi_flash.cmd_addr\[24\] _06999_ _07000_ net1506 _07002_ VGND VGND
+ VPWR VPWR _02286_ sky130_fd_sc_hd__o221a_1
XFILLER_0_39_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13236__758 clknet_1_1__leaf__08342_ VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__inv_2
X_16455_ CPU.registerFile\[20\]\[10\] CPU.registerFile\[21\]\[10\] _03883_ VGND VGND
+ VPWR VPWR _04172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_923 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10879_ CPU.aluReg\[8\] CPU.aluReg\[6\] _06939_ VGND VGND VPWR VPWR _06949_ sky130_fd_sc_hd__mux2_1
X_13784__1149 clknet_1_0__leaf__08463_ VGND VGND VPWR VPWR net1205 sky130_fd_sc_hd__inv_2
XFILLER_0_144_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15406_ CPU.registerFile\[19\]\[27\] CPU.registerFile\[18\]\[27\] _03157_ VGND VGND
+ VPWR VPWR _03461_ sky130_fd_sc_hd__mux2_1
X_12618_ _08000_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__clkbuf_1
X_19174_ clknet_leaf_6_clk _02694_ VGND VGND VPWR VPWR per_uart.uart0.rx_count16\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13598_ clknet_1_0__leaf__08440_ VGND VGND VPWR VPWR _08445_ sky130_fd_sc_hd__buf_1
X_16386_ CPU.registerFile\[8\]\[9\] _04101_ _04102_ _04103_ VGND VGND VPWR VPWR _04104_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18125_ net1136 _01653_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12549_ net2048 _07324_ _07957_ VGND VGND VPWR VPWR _07964_ sky130_fd_sc_hd__mux2_1
X_15337_ _03156_ _03391_ _03393_ _03163_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__a211o_1
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18056_ net1067 _01584_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1 CPU.mem_wbusy VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15268_ _03078_ _03324_ _03326_ _03043_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__a211o_1
X_17007_ CPU.registerFile\[2\]\[24\] CPU.registerFile\[3\]\[24\] _04431_ VGND VGND
+ VPWR VPWR _04710_ sky130_fd_sc_hd__mux2_1
X_14172__309 clknet_1_1__leaf__08501_ VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__inv_2
X_14219_ clknet_1_1__leaf__08339_ VGND VGND VPWR VPWR _08506_ sky130_fd_sc_hd__buf_1
X_15199_ _03006_ _03257_ _03259_ _03218_ VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_1__f__03645_ clknet_0__03645_ VGND VGND VPWR VPWR clknet_1_1__leaf__03645_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_834 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _05349_ _05532_ _05535_ CPU.aluReg\[19\] _06099_ VGND VGND VPWR VPWR _06100_
+ sky130_fd_sc_hd__a221o_1
X_18958_ net732 _02478_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17909_ clknet_leaf_22_clk _01437_ VGND VGND VPWR VPWR CPU.Jimm\[16\] sky130_fd_sc_hd__dfxtp_1
X_09691_ _06033_ VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__clkbuf_1
X_18889_ net663 _02409_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18592__49 VGND VGND VPWR VPWR _18592__49/HI net49 sky130_fd_sc_hd__conb_1
XFILLER_0_119_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09125_ _05476_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_162_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13701__1074 clknet_1_1__leaf__08455_ VGND VGND VPWR VPWR net1130 sky130_fd_sc_hd__inv_2
X_09056_ _05255_ _05256_ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__or2_2
Xhold540 CPU.registerFile\[27\]\[25\] VGND VGND VPWR VPWR net1837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 CPU.registerFile\[15\]\[27\] VGND VGND VPWR VPWR net1848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 CPU.registerFile\[13\]\[5\] VGND VGND VPWR VPWR net1859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15773__560 clknet_1_1__leaf__03655_ VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__inv_2
Xhold573 CPU.registerFile\[18\]\[16\] VGND VGND VPWR VPWR net1870 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold584 CPU.registerFile\[29\]\[10\] VGND VGND VPWR VPWR net1881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 CPU.registerFile\[30\]\[17\] VGND VGND VPWR VPWR net1892 sky130_fd_sc_hd__dlygate4sd3_1
X_09958_ _06202_ _06289_ _06177_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__o21a_1
X_08909_ CPU.aluIn1\[10\] _05260_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__and2_1
X_09889_ _06223_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__buf_4
Xhold1240 CPU.registerFile\[20\]\[1\] VGND VGND VPWR VPWR net2537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1251 CPU.PC\[17\] VGND VGND VPWR VPWR net2548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1262 CPU.registerFile\[1\]\[15\] VGND VGND VPWR VPWR net2559 sky130_fd_sc_hd__dlygate4sd3_1
X_11920_ _06649_ net2197 _07584_ VGND VGND VPWR VPWR _07590_ sky130_fd_sc_hd__mux2_1
Xhold1273 CPU.registerFile\[25\]\[14\] VGND VGND VPWR VPWR net2570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1284 CPU.registerFile\[9\]\[17\] VGND VGND VPWR VPWR net2581 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1295 CPU.registerFile\[24\]\[25\] VGND VGND VPWR VPWR net2592 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _07553_ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__clkbuf_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _06890_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__clkbuf_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _08808_ _08809_ CPU.registerFile\[25\]\[6\] VGND VGND VPWR VPWR _08810_ sky130_fd_sc_hd__a21o_1
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ _06647_ net1883 _07512_ VGND VGND VPWR VPWR _07517_ sky130_fd_sc_hd__mux2_1
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10733_ net2415 _06316_ _06838_ VGND VGND VPWR VPWR _06840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13452_ CPU.Iimm\[0\] _08412_ _08388_ VGND VGND VPWR VPWR _08413_ sky130_fd_sc_hd__mux2_1
X_16240_ _03959_ _03960_ _03961_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__mux2_1
X_10664_ net2533 _06337_ _06799_ VGND VGND VPWR VPWR _06802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12403_ _07886_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16171_ CPU.registerFile\[9\]\[4\] _03698_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10595_ _06764_ VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__clkbuf_1
X_13528__919 clknet_1_0__leaf__08437_ VGND VGND VPWR VPWR net975 sky130_fd_sc_hd__inv_2
X_15856__602 clknet_1_0__leaf__03681_ VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__inv_2
XFILLER_0_134_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12334_ _06599_ net1635 _07848_ VGND VGND VPWR VPWR _07850_ sky130_fd_sc_hd__mux2_1
X_15122_ _03138_ _03139_ CPU.registerFile\[9\]\[19\] VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__a21o_1
X_15053_ CPU.registerFile\[17\]\[18\] _03036_ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__or2_1
X_12265_ mapped_spi_ram.rcv_data\[16\] _07800_ VGND VGND VPWR VPWR _07806_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11216_ _05739_ _05737_ _05738_ VGND VGND VPWR VPWR _07199_ sky130_fd_sc_hd__and3_4
X_12196_ mapped_spi_ram.snd_bitcount\[3\] mapped_spi_ram.snd_bitcount\[2\] mapped_spi_ram.snd_bitcount\[1\]
+ mapped_spi_ram.snd_bitcount\[0\] VGND VGND VPWR VPWR _07758_ sky130_fd_sc_hd__or4_1
X_13954__112 clknet_1_0__leaf__08480_ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__inv_2
X_18812_ net601 _02336_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_11147_ net1611 _07147_ _07155_ _07151_ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18743_ net532 _02267_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[5\] sky130_fd_sc_hd__dfxtp_1
X_15955_ clknet_1_0__leaf__03686_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__buf_1
X_11078_ net1563 _07008_ _06985_ VGND VGND VPWR VPWR _07109_ sky130_fd_sc_hd__a21oi_1
X_14906_ CPU.registerFile\[15\]\[14\] CPU.registerFile\[14\]\[14\] _08771_ VGND VGND
+ VPWR VPWR _02974_ sky130_fd_sc_hd__mux2_1
X_10029_ CPU.cycles\[8\] _05552_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__nand2_1
X_18674_ net463 _02198_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17625_ net1894 VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__clkbuf_1
X_14837_ CPU.registerFile\[5\]\[12\] CPU.registerFile\[4\]\[12\] _08864_ VGND VGND
+ VPWR VPWR _02907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17556_ per_uart.uart0.tx_bitcount\[1\] per_uart.uart0.tx_bitcount\[0\] per_uart.uart0.tx_bitcount\[2\]
+ per_uart.uart0.tx_bitcount\[3\] VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__or4_1
XFILLER_0_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14768_ _02750_ _02817_ _02838_ _02839_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__a211o_1
X_16507_ CPU.registerFile\[9\]\[12\] _04056_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17487_ _05065_ _05066_ _05020_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14699_ CPU.registerFile\[24\]\[9\] _08686_ _02770_ _02771_ VGND VGND VPWR VPWR _02772_
+ sky130_fd_sc_hd__o211a_1
X_16438_ CPU.registerFile\[2\]\[10\] CPU.registerFile\[3\]\[10\] _04027_ VGND VGND
+ VPWR VPWR _04155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19157_ clknet_leaf_5_clk net1477 VGND VGND VPWR VPWR per_uart.uart0.txd_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16369_ _04086_ _04087_ _03961_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18108_ net1119 _01636_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19088_ net71 _02608_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_18039_ net1050 _01567_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09812_ _06148_ VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__buf_4
X_09743_ net2256 _06083_ _06055_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__mux2_1
X_09674_ _05423_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__buf_2
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09108_ _05262_ CPU.aluIn1\[8\] VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10380_ _06360_ VGND VGND VPWR VPWR _06645_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_131_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09039_ _05390_ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__buf_2
X_12050_ _07659_ VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold370 per_uart.rx_data\[0\] VGND VGND VPWR VPWR net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 CPU.registerFile\[19\]\[24\] VGND VGND VPWR VPWR net1678 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ CPU.PC\[13\] _07031_ _07043_ _07044_ _06853_ VGND VGND VPWR VPWR _07045_
+ sky130_fd_sc_hd__o221a_1
Xhold392 CPU.registerFile\[19\]\[16\] VGND VGND VPWR VPWR net1689 sky130_fd_sc_hd__dlygate4sd3_1
X_13783__1148 clknet_1_0__leaf__08463_ VGND VGND VPWR VPWR net1204 sky130_fd_sc_hd__inv_2
X_15851__598 clknet_1_1__leaf__03680_ VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__inv_2
XFILLER_0_99_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12952_ _06530_ net1655 _08144_ VGND VGND VPWR VPWR _08178_ sky130_fd_sc_hd__mux2_1
Xhold1070 CPU.registerFile\[11\]\[0\] VGND VGND VPWR VPWR net2367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 CPU.registerFile\[14\]\[21\] VGND VGND VPWR VPWR net2378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1092 CPU.registerFile\[8\]\[7\] VGND VGND VPWR VPWR net2389 sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ _06632_ net2016 _07573_ VGND VGND VPWR VPWR _07581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _08141_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__clkbuf_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _08857_ _08858_ _08860_ _08661_ VGND VGND VPWR VPWR _08861_ sky130_fd_sc_hd__a211o_1
XFILLER_0_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _07544_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__clkbuf_1
X_18390_ net211 _01918_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03648_ clknet_0__03648_ VGND VGND VPWR VPWR clknet_1_0__leaf__03648_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11765_ _06630_ net2205 _07501_ VGND VGND VPWR VPWR _07508_ sky130_fd_sc_hd__mux2_1
X_14553_ CPU.registerFile\[19\]\[6\] CPU.registerFile\[18\]\[6\] _06064_ VGND VGND
+ VPWR VPWR _08793_ sky130_fd_sc_hd__mux2_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10716_ net1816 _06124_ _06827_ VGND VGND VPWR VPWR _06831_ sky130_fd_sc_hd__mux2_1
X_17272_ _03714_ _04963_ _04967_ _08403_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11696_ net2535 _07345_ _07464_ VGND VGND VPWR VPWR _07471_ sky130_fd_sc_hd__mux2_1
X_14484_ CPU.registerFile\[27\]\[4\] CPU.registerFile\[26\]\[4\] _06063_ VGND VGND
+ VPWR VPWR _08726_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19011_ clknet_leaf_12_clk _02531_ VGND VGND VPWR VPWR CPU.aluIn1\[28\] sky130_fd_sc_hd__dfxtp_2
X_16223_ _03726_ _03727_ CPU.registerFile\[1\]\[5\] VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__a21o_1
X_10647_ net2496 _06145_ _06788_ VGND VGND VPWR VPWR _06793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13435_ _08399_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16154_ _03749_ _03751_ CPU.registerFile\[25\]\[3\] VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10578_ _06755_ VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14021__172 clknet_1_0__leaf__08487_ VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__inv_2
X_15105_ _03078_ _03165_ _03167_ _03043_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__a211o_1
X_12317_ net1306 _07781_ VGND VGND VPWR VPWR _07839_ sky130_fd_sc_hd__nor2_1
X_14095__240 clknet_1_0__leaf__08493_ VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__inv_2
X_16085_ CPU.registerFile\[16\]\[1\] _06173_ _03769_ _03810_ VGND VGND VPWR VPWR _03811_
+ sky130_fd_sc_hd__o211a_1
X_13580__965 clknet_1_0__leaf__08443_ VGND VGND VPWR VPWR net1021 sky130_fd_sc_hd__inv_2
X_15036_ CPU.registerFile\[8\]\[17\] _03018_ _03100_ _02864_ VGND VGND VPWR VPWR _03101_
+ sky130_fd_sc_hd__o211a_1
X_12248_ net1535 _07785_ _07795_ _07796_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12179_ net1341 _07738_ _07748_ _07737_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16987_ _04689_ _04690_ _04365_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18726_ net515 net1579 VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13700__1073 clknet_1_1__leaf__08455_ VGND VGND VPWR VPWR net1129 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__05014_ clknet_0__05014_ VGND VGND VPWR VPWR clknet_1_1__leaf__05014_
+ sky130_fd_sc_hd__clkbuf_16
X_18657_ clknet_leaf_12_clk _02181_ VGND VGND VPWR VPWR CPU.rs2\[29\] sky130_fd_sc_hd__dfxtp_1
X_17608_ per_uart.d_in_uart\[3\] _05134_ _05157_ per_uart.uart0.txd_reg\[4\] VGND
+ VGND VPWR VPWR _05162_ sky130_fd_sc_hd__o22a_1
X_09390_ _05741_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18588_ net409 net45 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17539_ _08310_ _06016_ net13 VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__or3_1
XFILLER_0_74_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13331__830 clknet_1_1__leaf__08364_ VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__inv_2
XFILLER_0_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__08497_ clknet_0__08497_ VGND VGND VPWR VPWR clknet_1_1__leaf__08497_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14150__289 clknet_1_1__leaf__08499_ VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__inv_2
X_09726_ _05893_ _06066_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09657_ _05997_ _06000_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__nand2_1
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ CPU.PC\[17\] _05930_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__nor2_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11550_ net1838 _07337_ _07390_ VGND VGND VPWR VPWR _07393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10501_ _06714_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11481_ net2073 _07349_ _07333_ VGND VGND VPWR VPWR _07350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13220_ _08333_ VGND VGND VPWR VPWR _08334_ sky130_fd_sc_hd__clkbuf_2
X_10432_ _06677_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13151_ _08283_ _08284_ VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__nor2_1
X_10363_ _06633_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__clkbuf_1
X_12102_ _07695_ VGND VGND VPWR VPWR _07696_ sky130_fd_sc_hd__clkbuf_4
X_13925__86 clknet_1_0__leaf__08477_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__inv_2
X_13082_ CPU.registerFile\[4\]\[4\] net1391 _08239_ VGND VGND VPWR VPWR _08247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10294_ _06587_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12033_ _07650_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__clkbuf_1
X_16910_ CPU.registerFile\[20\]\[21\] CPU.registerFile\[21\]\[21\] _04287_ VGND VGND
+ VPWR VPWR _04616_ sky130_fd_sc_hd__mux2_1
X_17890_ clknet_leaf_26_clk _01418_ VGND VGND VPWR VPWR CPU.mem_wmask\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16841_ CPU.registerFile\[8\]\[20\] _04505_ _04506_ _04547_ VGND VGND VPWR VPWR _04548_
+ sky130_fd_sc_hd__o211a_1
X_16772_ CPU.registerFile\[28\]\[18\] CPU.registerFile\[29\]\[18\] _04122_ VGND VGND
+ VPWR VPWR _04481_ sky130_fd_sc_hd__mux2_1
X_18511_ net332 _02035_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ _08169_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ net263 _01970_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _06316_ net1881 _08131_ VGND VGND VPWR VPWR _08133_ sky130_fd_sc_hd__mux2_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ CPU.registerFile\[30\]\[7\] CPU.registerFile\[31\]\[7\] _08645_ VGND VGND
+ VPWR VPWR _08844_ sky130_fd_sc_hd__mux2_1
X_11817_ _07535_ VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__clkbuf_1
X_18373_ net194 _01901_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _03627_ _03635_ _05861_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__o21a_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _06653_ net2515 _08087_ VGND VGND VPWR VPWR _08095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14536_ _08567_ _08569_ CPU.registerFile\[9\]\[5\] VGND VGND VPWR VPWR _08777_ sky130_fd_sc_hd__a21o_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11748_ _06613_ net2408 _07490_ VGND VGND VPWR VPWR _07499_ sky130_fd_sc_hd__mux2_1
X_17255_ _03766_ _04948_ _04950_ _03716_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__a211o_1
X_14467_ _08574_ _08704_ _08709_ _08592_ VGND VGND VPWR VPWR _08710_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11679_ net2582 _07328_ _07453_ VGND VGND VPWR VPWR _07462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16206_ _03919_ _03928_ _08406_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__o21a_1
X_13418_ _08265_ VGND VGND VPWR VPWR _08388_ sky130_fd_sc_hd__buf_4
X_17186_ _04882_ _04883_ _04557_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__mux2_1
X_14398_ CPU.registerFile\[21\]\[2\] _08528_ VGND VGND VPWR VPWR _08642_ sky130_fd_sc_hd__or2_1
Xclkbuf_0__08451_ _08451_ VGND VGND VPWR VPWR clknet_0__08451_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16137_ CPU.registerFile\[13\]\[3\] _03709_ VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16068_ _03716_ _03789_ _03793_ _03732_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__o211a_1
X_15019_ _03078_ _03079_ _03083_ _03043_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__a211o_1
X_08890_ CPU.instr\[3\] CPU.instr\[2\] VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__or2_1
X_13506__899 clknet_1_1__leaf__08435_ VGND VGND VPWR VPWR net955 sky130_fd_sc_hd__inv_2
X_15834__582 clknet_1_0__leaf__03679_ VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__inv_2
X_13361__856 clknet_1_1__leaf__08368_ VGND VGND VPWR VPWR net912 sky130_fd_sc_hd__inv_2
X_17425__46 clknet_1_1__leaf__05015_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__inv_2
X_09511_ _05855_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18709_ net498 _02233_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[9\] sky130_fd_sc_hd__dfxtp_1
X_09442_ CPU.aluIn1\[28\] _05257_ _05532_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__and3_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09373_ _05691_ _05722_ _05723_ _05724_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__a31o_1
XFILLER_0_137_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13782__1147 clknet_1_1__leaf__08463_ VGND VGND VPWR VPWR net1203 sky130_fd_sc_hd__inv_2
XFILLER_0_74_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15917__657 clknet_1_0__leaf__03687_ VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__inv_2
XFILLER_0_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__08440_ clknet_0__08440_ VGND VGND VPWR VPWR clknet_1_0__leaf__08440_
+ sky130_fd_sc_hd__clkbuf_16
X_09709_ _06050_ _06002_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__xnor2_1
X_10981_ CPU.aluIn1\[13\] CPU.aluIn1\[12\] _05545_ VGND VGND VPWR VPWR _07027_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12720_ _08054_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__clkbuf_1
X_13338__836 clknet_1_1__leaf__08365_ VGND VGND VPWR VPWR net892 sky130_fd_sc_hd__inv_2
XFILLER_0_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15963__699 clknet_1_0__leaf__03691_ VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__inv_2
XFILLER_0_38_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12651_ _06643_ net1748 _08015_ VGND VGND VPWR VPWR _08018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11602_ net2166 _07320_ _07416_ VGND VGND VPWR VPWR _07421_ sky130_fd_sc_hd__mux2_1
X_12582_ _07981_ VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__clkbuf_1
X_15370_ CPU.registerFile\[19\]\[26\] CPU.registerFile\[18\]\[26\] _03157_ VGND VGND
+ VPWR VPWR _03426_ sky130_fd_sc_hd__mux2_1
X_17304__719 clknet_1_1__leaf__04980_ VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__inv_2
XFILLER_0_154_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14321_ _08566_ VGND VGND VPWR VPWR _08567_ sky130_fd_sc_hd__buf_4
XFILLER_0_80_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11533_ net2479 _07320_ _07379_ VGND VGND VPWR VPWR _07384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17040_ CPU.registerFile\[6\]\[25\] CPU.registerFile\[7\]\[25\] _04426_ VGND VGND
+ VPWR VPWR _04742_ sky130_fd_sc_hd__mux2_1
X_11464_ _07338_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17352__12 clknet_1_0__leaf__04985_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__inv_2
XFILLER_0_162_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10415_ _06668_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__clkbuf_1
X_13203_ _06157_ _06252_ _06319_ _08316_ VGND VGND VPWR VPWR _08317_ sky130_fd_sc_hd__or4_1
XFILLER_0_150_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11395_ net1713 _06267_ _07285_ VGND VGND VPWR VPWR _07295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10346_ _06105_ VGND VGND VPWR VPWR _06622_ sky130_fd_sc_hd__buf_4
X_13134_ _08273_ net1576 VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18991_ clknet_leaf_13_clk _02511_ VGND VGND VPWR VPWR CPU.aluIn1\[8\] sky130_fd_sc_hd__dfxtp_4
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ CPU.registerFile\[4\]\[12\] net1406 _08228_ VGND VGND VPWR VPWR _08238_ sky130_fd_sc_hd__mux2_1
X_17942_ net953 _01470_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_10277_ _06578_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12016_ _07641_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__clkbuf_1
X_17873_ clknet_leaf_23_clk _00022_ VGND VGND VPWR VPWR CPU.cycles\[16\] sky130_fd_sc_hd__dfxtp_1
X_14133__273 clknet_1_0__leaf__08498_ VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__inv_2
X_16824_ _04441_ _04529_ _04531_ _04208_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__a211o_1
XFILLER_0_136_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16755_ CPU.registerFile\[15\]\[18\] CPU.registerFile\[14\]\[18\] _04146_ VGND VGND
+ VPWR VPWR _04464_ sky130_fd_sc_hd__mux2_1
X_12918_ _08160_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16686_ CPU.registerFile\[28\]\[16\] CPU.registerFile\[29\]\[16\] _04122_ VGND VGND
+ VPWR VPWR _04397_ sky130_fd_sc_hd__mux2_1
X_13898_ clknet_1_1__leaf__08473_ VGND VGND VPWR VPWR _08475_ sky130_fd_sc_hd__buf_1
X_18425_ net246 _01953_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _06124_ net2222 _08120_ VGND VGND VPWR VPWR _08124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18356_ net177 _01884_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ _08592_ _03606_ _03610_ _03618_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15721__513 clknet_1_0__leaf__03650_ VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__inv_2
XFILLER_0_28_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17307_ clknet_1_0__leaf__03686_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__buf_1
X_14519_ _08521_ _08757_ _08759_ _08533_ VGND VGND VPWR VPWR _08760_ sky130_fd_sc_hd__a211o_1
X_18287_ net108 _01815_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_15499_ _08546_ _08547_ CPU.registerFile\[9\]\[29\] VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13586__971 clknet_1_1__leaf__08443_ VGND VGND VPWR VPWR net1027 sky130_fd_sc_hd__inv_2
X_17238_ CPU.registerFile\[20\]\[30\] CPU.registerFile\[21\]\[30\] _03737_ VGND VGND
+ VPWR VPWR _04935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_834 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08503_ _08503_ VGND VGND VPWR VPWR clknet_0__08503_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold903 _02670_ VGND VGND VPWR VPWR net2200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold914 CPU.registerFile\[4\]\[20\] VGND VGND VPWR VPWR net2211 sky130_fd_sc_hd__dlygate4sd3_1
X_17169_ _04579_ _04580_ CPU.registerFile\[17\]\[28\] VGND VGND VPWR VPWR _04868_
+ sky130_fd_sc_hd__a21o_1
Xhold925 CPU.registerFile\[29\]\[18\] VGND VGND VPWR VPWR net2222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 CPU.registerFile\[31\]\[3\] VGND VGND VPWR VPWR net2233 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__08434_ _08434_ VGND VGND VPWR VPWR clknet_0__08434_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold947 CPU.registerFile\[20\]\[3\] VGND VGND VPWR VPWR net2244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold958 CPU.registerFile\[17\]\[29\] VGND VGND VPWR VPWR net2255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 CPU.registerFile\[26\]\[23\] VGND VGND VPWR VPWR net2266 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ _05263_ _05307_ VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13904__67 clknet_1_0__leaf__08475_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__inv_2
Xclkbuf_0__08365_ _08365_ VGND VGND VPWR VPWR clknet_0__08365_ sky130_fd_sc_hd__clkbuf_16
X_08942_ CPU.aluIn1\[7\] _05293_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09425_ _05402_ _05407_ _05410_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09356_ CPU.PC\[4\] _05643_ _05707_ _05703_ VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__o211a_2
XFILLER_0_47_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09287_ _05629_ _05632_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__xor2_1
XFILLER_0_90_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10200_ _06519_ _06521_ VGND VGND VPWR VPWR _06522_ sky130_fd_sc_hd__xnor2_2
X_11180_ net1379 _07132_ _07173_ _07164_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__o211a_1
X_10131_ _06061_ VGND VGND VPWR VPWR _06456_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10062_ net1375 _05860_ _05719_ per_uart.rx_data\[6\] _06388_ VGND VGND VPWR VPWR
+ _06389_ sky130_fd_sc_hd__a221o_1
X_14870_ CPU.registerFile\[10\]\[13\] CPU.registerFile\[11\]\[13\] _02779_ VGND VGND
+ VPWR VPWR _02939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17404__27 clknet_1_1__leaf__05013_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__inv_2
XFILLER_0_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16540_ _03963_ _04251_ _04254_ _04006_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__a211o_1
X_10964_ net1520 _07007_ _07013_ _07014_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__o211a_1
X_12703_ _08045_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__clkbuf_1
X_16471_ _04099_ _04184_ _04186_ _04105_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__a211o_1
XFILLER_0_155_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10895_ CPU.aluReg\[4\] CPU.aluReg\[2\] _06939_ VGND VGND VPWR VPWR _06961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18210_ net1221 _01738_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[11\] sky130_fd_sc_hd__dfxtp_1
X_15422_ _03202_ _03464_ _03468_ _03476_ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__a31o_1
X_12634_ _06626_ net1968 _08004_ VGND VGND VPWR VPWR _08009_ sky130_fd_sc_hd__mux2_1
X_19190_ clknet_leaf_3_clk _02708_ VGND VGND VPWR VPWR per_uart.d_in_uart\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18141_ net1152 _01669_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15353_ _03408_ _03409_ _08541_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12565_ _07972_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__clkbuf_1
X_14304_ _08549_ VGND VGND VPWR VPWR _08550_ sky130_fd_sc_hd__clkbuf_4
X_18072_ net1083 _01600_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11516_ _07373_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15284_ _03098_ _03340_ _03342_ _03307_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__a211o_1
XFILLER_0_123_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12496_ _07935_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17023_ _04724_ _04725_ _04365_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__mux2_1
X_11447_ net1985 _07326_ _07312_ VGND VGND VPWR VPWR _07327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11378_ _07286_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__clkbuf_1
X_10329_ _06610_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__clkbuf_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _08265_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__clkbuf_4
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ clknet_1_1__leaf__08484_ VGND VGND VPWR VPWR _08494_ sky130_fd_sc_hd__buf_1
X_18974_ net748 _02494_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ net2498 VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__clkbuf_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925_ net936 _01453_ VGND VGND VPWR VPWR CPU.aluShamt\[0\] sky130_fd_sc_hd__dfxtp_1
X_17856_ _00013_ _00014_ VGND VGND VPWR VPWR CPU.writeBack sky130_fd_sc_hd__dlxtn_4
X_13781__1146 clknet_1_1__leaf__08463_ VGND VGND VPWR VPWR net1202 sky130_fd_sc_hd__inv_2
XFILLER_0_89_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16807_ CPU.registerFile\[6\]\[19\] CPU.registerFile\[7\]\[19\] _04426_ VGND VGND
+ VPWR VPWR _04515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17787_ net867 _01349_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_14999_ CPU.registerFile\[5\]\[16\] CPU.registerFile\[4\]\[16\] _08864_ VGND VGND
+ VPWR VPWR _03065_ sky130_fd_sc_hd__mux2_1
X_16738_ CPU.registerFile\[22\]\[17\] CPU.registerFile\[23\]\[17\] _04362_ VGND VGND
+ VPWR VPWR _04448_ sky130_fd_sc_hd__mux2_1
X_15946__683 clknet_1_0__leaf__03690_ VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__inv_2
XFILLER_0_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16669_ _03744_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__buf_2
XFILLER_0_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09210_ CPU.aluIn1\[19\] _05543_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__or2_1
X_18408_ net229 _01936_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09141_ _05375_ CPU.aluIn1\[22\] VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__and2b_1
X_18339_ net160 _01867_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09072_ _05423_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold700 CPU.registerFile\[20\]\[29\] VGND VGND VPWR VPWR net1997 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold711 CPU.registerFile\[22\]\[31\] VGND VGND VPWR VPWR net2008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 CPU.registerFile\[9\]\[24\] VGND VGND VPWR VPWR net2019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 CPU.registerFile\[9\]\[26\] VGND VGND VPWR VPWR net2030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold744 CPU.registerFile\[21\]\[6\] VGND VGND VPWR VPWR net2041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold755 CPU.registerFile\[21\]\[26\] VGND VGND VPWR VPWR net2052 sky130_fd_sc_hd__dlygate4sd3_1
Xhold766 CPU.registerFile\[11\]\[4\] VGND VGND VPWR VPWR net2063 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 CPU.registerFile\[6\]\[9\] VGND VGND VPWR VPWR net2074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 CPU.registerFile\[6\]\[13\] VGND VGND VPWR VPWR net2085 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ _05974_ _05944_ VGND VGND VPWR VPWR _06305_ sky130_fd_sc_hd__and2b_1
Xhold799 CPU.registerFile\[30\]\[18\] VGND VGND VPWR VPWR net2096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08925_ CPU.Iimm\[1\] VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__inv_2
X_17333__745 clknet_1_0__leaf__04983_ VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__inv_2
X_15691__486 clknet_1_0__leaf__03647_ VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__inv_2
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03681_ clknet_0__03681_ VGND VGND VPWR VPWR clknet_1_0__leaf__03681_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09408_ _05552_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__buf_4
X_10680_ net2593 _06530_ _06776_ VGND VGND VPWR VPWR _06810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09339_ _05577_ _05579_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__xor2_4
XFILLER_0_8_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12350_ _06615_ net2107 _07848_ VGND VGND VPWR VPWR _07858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11301_ _07245_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__clkbuf_1
X_12281_ mapped_spi_ram.rcv_data\[9\] _07812_ _07815_ _07809_ VGND VGND VPWR VPWR
+ _01699_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_889 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14020_ clknet_1_0__leaf__08484_ VGND VGND VPWR VPWR _08487_ sky130_fd_sc_hd__buf_1
X_11232_ _07208_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__clkbuf_1
X_11163_ mapped_spi_flash.rcv_data\[9\] _07149_ VGND VGND VPWR VPWR _07165_ sky130_fd_sc_hd__or2_1
X_13641__1021 clknet_1_0__leaf__08448_ VGND VGND VPWR VPWR net1077 sky130_fd_sc_hd__inv_2
X_10114_ _06439_ VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__buf_4
X_15971_ _03697_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__buf_4
X_11094_ net1456 _07119_ _07121_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__a21boi_1
X_17710_ CPU.mem_wdata\[6\] per_uart.d_in_uart\[6\] _05218_ VGND VGND VPWR VPWR _05231_
+ sky130_fd_sc_hd__mux2_1
X_14922_ _02826_ _02985_ _02989_ _02746_ VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__o211a_1
X_10045_ _05292_ _05303_ VGND VGND VPWR VPWR _06373_ sky130_fd_sc_hd__or2b_1
X_18690_ net479 _02214_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold60 _06540_ VGND VGND VPWR VPWR net1357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold71 _06439_ VGND VGND VPWR VPWR net1368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 mapped_spi_flash.rcv_data\[0\] VGND VGND VPWR VPWR net1379 sky130_fd_sc_hd__clkbuf_2
X_17641_ _07108_ net1660 VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__nor2_1
X_14853_ CPU.registerFile\[20\]\[13\] _08839_ _02921_ _08841_ VGND VGND VPWR VPWR
+ _02922_ sky130_fd_sc_hd__o211a_1
Xhold93 mapped_spi_flash.rcv_data\[28\] VGND VGND VPWR VPWR net1390 sky130_fd_sc_hd__dlygate4sd3_1
X_17572_ _05132_ _05135_ _06856_ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__o21a_1
X_14784_ CPU.registerFile\[24\]\[11\] _08686_ _02854_ _02771_ VGND VGND VPWR VPWR
+ _02855_ sky130_fd_sc_hd__o211a_1
X_11996_ _06657_ net2314 _07620_ VGND VGND VPWR VPWR _07630_ sky130_fd_sc_hd__mux2_1
X_16523_ _04098_ _04224_ _04228_ _04237_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__a31o_4
XFILLER_0_156_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10947_ mapped_spi_flash.cmd_addr\[25\] _06999_ _07000_ net1530 _07002_ VGND VGND
+ VPWR VPWR _02287_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_926 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14245__374 clknet_1_0__leaf__08509_ VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__inv_2
X_16454_ CPU.registerFile\[22\]\[10\] CPU.registerFile\[23\]\[10\] _03958_ VGND VGND
+ VPWR VPWR _04171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10878_ _06948_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15405_ net1595 _03201_ _03460_ _03390_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__o211a_1
X_12617_ _06609_ net1837 _07993_ VGND VGND VPWR VPWR _08000_ sky130_fd_sc_hd__mux2_1
X_19173_ clknet_leaf_5_clk _02693_ VGND VGND VPWR VPWR per_uart.uart0.rx_count16\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16385_ CPU.registerFile\[9\]\[9\] _04056_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18124_ net1135 _01652_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_15336_ CPU.registerFile\[16\]\[25\] _03159_ _03392_ _03161_ VGND VGND VPWR VPWR
+ _03393_ sky130_fd_sc_hd__o211a_1
X_12548_ _07963_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18055_ net1066 _01583_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_15267_ CPU.registerFile\[20\]\[23\] _03080_ _03325_ _03082_ VGND VGND VPWR VPWR
+ _03326_ sky130_fd_sc_hd__o211a_1
X_12479_ _07926_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_2 CPU.mem_wdata\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17006_ _04707_ _04708_ _04557_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03644_ clknet_0__03644_ VGND VGND VPWR VPWR clknet_1_1__leaf__03644_
+ sky130_fd_sc_hd__clkbuf_16
X_15198_ CPU.registerFile\[24\]\[21\] _02928_ _03258_ _03175_ VGND VGND VPWR VPWR
+ _03259_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18957_ net731 _02477_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17908_ clknet_leaf_22_clk _01436_ VGND VGND VPWR VPWR CPU.Jimm\[15\] sky130_fd_sc_hd__dfxtp_1
X_09690_ net2283 _06032_ _05742_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__mux2_1
X_18888_ net662 _02408_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_17839_ net919 _01401_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09124_ _05475_ _05346_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09055_ _05394_ _05398_ _05405_ _05406_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__o31a_1
XFILLER_0_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold530 CPU.registerFile\[13\]\[4\] VGND VGND VPWR VPWR net1827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold541 CPU.registerFile\[6\]\[19\] VGND VGND VPWR VPWR net1838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 CPU.registerFile\[15\]\[7\] VGND VGND VPWR VPWR net1849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 CPU.registerFile\[28\]\[24\] VGND VGND VPWR VPWR net1860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 CPU.registerFile\[12\]\[24\] VGND VGND VPWR VPWR net1871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 CPU.registerFile\[3\]\[31\] VGND VGND VPWR VPWR net1882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 per_uart.rx_data\[1\] VGND VGND VPWR VPWR net1893 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09957_ _06204_ _06287_ _06288_ _05855_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__o22a_1
X_08908_ CPU.rs2\[10\] CPU.Bimm\[10\] _05245_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__mux2_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _06208_ _06209_ _06217_ _06222_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__or4b_4
Xhold1230 CPU.registerFile\[17\]\[5\] VGND VGND VPWR VPWR net2527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 CPU.registerFile\[26\]\[30\] VGND VGND VPWR VPWR net2538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 CPU.registerFile\[12\]\[28\] VGND VGND VPWR VPWR net2549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1263 CPU.registerFile\[8\]\[5\] VGND VGND VPWR VPWR net2560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 CPU.registerFile\[26\]\[2\] VGND VGND VPWR VPWR net2571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1285 CPU.registerFile\[8\]\[23\] VGND VGND VPWR VPWR net2582 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1296 CPU.registerFile\[1\]\[1\] VGND VGND VPWR VPWR net2593 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ net2588 _07362_ _07548_ VGND VGND VPWR VPWR _07553_ sky130_fd_sc_hd__mux2_1
X_18568__25 VGND VGND VPWR VPWR _18568__25/HI net25 sky130_fd_sc_hd__conb_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10801_ net2667 _06888_ _06889_ VGND VGND VPWR VPWR _06890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _07516_ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__clkbuf_1
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13520_ clknet_1_0__leaf__08366_ VGND VGND VPWR VPWR _08437_ sky130_fd_sc_hd__buf_1
X_10732_ _06839_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13451_ _08411_ VGND VGND VPWR VPWR _08412_ sky130_fd_sc_hd__buf_4
XFILLER_0_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10663_ _06801_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__clkbuf_1
X_12402_ net1672 _07314_ _07884_ VGND VGND VPWR VPWR _07886_ sky130_fd_sc_hd__mux2_1
X_16170_ CPU.registerFile\[10\]\[4\] CPU.registerFile\[11\]\[4\] _03694_ VGND VGND
+ VPWR VPWR _03893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10594_ net2175 _06337_ _06761_ VGND VGND VPWR VPWR _06764_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13780__1145 clknet_1_1__leaf__08463_ VGND VGND VPWR VPWR net1201 sky130_fd_sc_hd__inv_2
X_15121_ CPU.registerFile\[10\]\[19\] CPU.registerFile\[11\]\[19\] _03183_ VGND VGND
+ VPWR VPWR _03184_ sky130_fd_sc_hd__mux2_1
X_12333_ _07849_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15052_ CPU.registerFile\[19\]\[18\] CPU.registerFile\[18\]\[18\] _02753_ VGND VGND
+ VPWR VPWR _03116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12264_ net1566 _07799_ _07805_ _07796_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__o211a_1
X_11215_ _07108_ _07198_ VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__nor2_1
X_12195_ net1318 _07692_ _07757_ _07755_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__o211a_1
X_18811_ net600 _02335_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11146_ net1384 _07149_ VGND VGND VPWR VPWR _07155_ sky130_fd_sc_hd__or2_1
X_11077_ _05237_ VGND VGND VPWR VPWR _07108_ sky130_fd_sc_hd__buf_4
X_18742_ net531 _02266_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[4\] sky130_fd_sc_hd__dfxtp_1
X_13242__763 clknet_1_0__leaf__08343_ VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__inv_2
X_10028_ _05885_ _06356_ VGND VGND VPWR VPWR _06357_ sky130_fd_sc_hd__or2_1
X_14905_ _02798_ _02958_ _02963_ _02972_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__a31o_1
X_18673_ net462 _02197_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_14836_ CPU.registerFile\[6\]\[12\] CPU.registerFile\[7\]\[12\] _08740_ VGND VGND
+ VPWR VPWR _02906_ sky130_fd_sc_hd__mux2_1
X_17624_ net1893 per_uart.uart0.rxd_reg\[2\] _05170_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17555_ _05122_ per_uart.uart0.tx_bitcount\[0\] _05116_ VGND VGND VPWR VPWR _05123_
+ sky130_fd_sc_hd__and3_1
X_14767_ _08596_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__clkbuf_4
X_11979_ _07621_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__clkbuf_1
X_16506_ CPU.registerFile\[10\]\[12\] CPU.registerFile\[11\]\[12\] _03931_ VGND VGND
+ VPWR VPWR _04221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17486_ _05055_ _06264_ _05061_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__or3_1
X_14698_ _06035_ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16437_ _04151_ _04152_ _04153_ VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13861__1219 clknet_1_1__leaf__08470_ VGND VGND VPWR VPWR net1275 sky130_fd_sc_hd__inv_2
XFILLER_0_128_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19156_ clknet_leaf_3_clk net1475 VGND VGND VPWR VPWR per_uart.uart0.txd_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16368_ CPU.registerFile\[20\]\[8\] CPU.registerFile\[21\]\[8\] _03883_ VGND VGND
+ VPWR VPWR _04087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18107_ net1118 _01635_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15319_ CPU.registerFile\[8\]\[24\] _03018_ _03376_ _03268_ VGND VGND VPWR VPWR _03377_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19087_ clknet_leaf_0_clk _02607_ VGND VGND VPWR VPWR per_uart.uart0.rxd_reg\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16299_ CPU.registerFile\[13\]\[7\] _03976_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18038_ net1049 _01566_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09811_ mapped_spi_flash.rcv_data\[8\] _05698_ _06147_ VGND VGND VPWR VPWR _06148_
+ sky130_fd_sc_hd__a21oi_4
X_09742_ _06082_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__buf_4
XFILLER_0_118_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09673_ _05894_ _06015_ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__or2_1
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13640__1020 clknet_1_0__leaf__08448_ VGND VGND VPWR VPWR net1076 sky130_fd_sc_hd__inv_2
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09107_ CPU.aluIn1\[11\] VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__inv_2
XFILLER_0_162_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09038_ _05388_ _05389_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17339__751 clknet_1_1__leaf__04983_ VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__inv_2
Xhold360 CPU.rs2\[21\] VGND VGND VPWR VPWR net1657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 _05171_ VGND VGND VPWR VPWR net1668 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold382 CPU.registerFile\[5\]\[7\] VGND VGND VPWR VPWR net1679 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ _05606_ _05609_ _07042_ _07023_ VGND VGND VPWR VPWR _07044_ sky130_fd_sc_hd__a31o_1
Xhold393 CPU.registerFile\[19\]\[17\] VGND VGND VPWR VPWR net1690 sky130_fd_sc_hd__dlygate4sd3_1
X_12951_ _08177_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1060 CPU.registerFile\[26\]\[7\] VGND VGND VPWR VPWR net2357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 CPU.registerFile\[12\]\[29\] VGND VGND VPWR VPWR net2368 sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ _07580_ VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__clkbuf_1
Xhold1082 CPU.registerFile\[29\]\[21\] VGND VGND VPWR VPWR net2379 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1093 CPU.registerFile\[7\]\[16\] VGND VGND VPWR VPWR net2390 sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ _06508_ net2232 _08131_ VGND VGND VPWR VPWR _08141_ sky130_fd_sc_hd__mux2_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ CPU.registerFile\[8\]\[7\] _08776_ _08859_ _08622_ VGND VGND VPWR VPWR _08860_
+ sky130_fd_sc_hd__o211a_1
X_13534__924 clknet_1_0__leaf__08438_ VGND VGND VPWR VPWR net980 sky130_fd_sc_hd__inv_2
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11833_ net2154 _07345_ _07537_ VGND VGND VPWR VPWR _07544_ sky130_fd_sc_hd__mux2_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03647_ clknet_0__03647_ VGND VGND VPWR VPWR clknet_1_0__leaf__03647_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ clknet_1_1__leaf__08340_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__buf_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ CPU.mem_wdata\[5\] _08514_ _08792_ _08751_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__o211a_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _07507_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__clkbuf_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _03722_ _04964_ _04966_ _03730_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__a211o_1
XFILLER_0_83_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _06830_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__clkbuf_1
X_14483_ _08723_ _08724_ _08609_ VGND VGND VPWR VPWR _08725_ sky130_fd_sc_hd__mux2_1
X_11695_ _07470_ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19010_ clknet_leaf_11_clk _02530_ VGND VGND VPWR VPWR CPU.aluIn1\[27\] sky130_fd_sc_hd__dfxtp_1
X_16222_ CPU.registerFile\[2\]\[5\] CPU.registerFile\[3\]\[5\] _03693_ VGND VGND VPWR
+ VPWR _03944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13434_ CPU.Jimm\[16\] _08398_ _08388_ VGND VGND VPWR VPWR _08399_ sky130_fd_sc_hd__mux2_1
X_10646_ _06792_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16153_ CPU.registerFile\[27\]\[3\] CPU.registerFile\[26\]\[3\] _03837_ VGND VGND
+ VPWR VPWR _03877_ sky130_fd_sc_hd__mux2_1
X_10577_ net2029 _06145_ _06750_ VGND VGND VPWR VPWR _06755_ sky130_fd_sc_hd__mux2_1
X_15104_ CPU.registerFile\[20\]\[19\] _03080_ _03166_ _03082_ VGND VGND VPWR VPWR
+ _03167_ sky130_fd_sc_hd__o211a_1
X_12316_ _07779_ net1303 VGND VGND VPWR VPWR _07838_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16084_ _03770_ _03771_ CPU.registerFile\[17\]\[1\] VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__a21o_1
X_15035_ _02733_ _02734_ CPU.registerFile\[9\]\[17\] VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__a21o_1
X_12247_ _07163_ VGND VGND VPWR VPWR _07796_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12178_ mapped_spi_ram.cmd_addr\[6\] _07694_ _07706_ CPU.mem_wdata\[7\] _07739_ VGND
+ VGND VPWR VPWR _07748_ sky130_fd_sc_hd__a221o_1
X_11129_ _05688_ _07132_ VGND VGND VPWR VPWR _07145_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16986_ CPU.registerFile\[20\]\[23\] CPU.registerFile\[21\]\[23\] _03737_ VGND VGND
+ VPWR VPWR _04690_ sky130_fd_sc_hd__mux2_1
X_18725_ net514 _02249_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__05013_ clknet_0__05013_ VGND VGND VPWR VPWR clknet_1_1__leaf__05013_
+ sky130_fd_sc_hd__clkbuf_16
X_18656_ clknet_leaf_11_clk _02180_ VGND VGND VPWR VPWR CPU.rs2\[28\] sky130_fd_sc_hd__dfxtp_1
X_17607_ net1532 _05159_ _05161_ _07108_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__o22a_1
X_14819_ CPU.registerFile\[28\]\[12\] CPU.registerFile\[29\]\[12\] _02808_ VGND VGND
+ VPWR VPWR _02889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15799_ net1508 _08350_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__nand2_1
X_18587_ net408 net44 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17538_ _05075_ _05025_ _06029_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17469_ _05022_ _06322_ _08256_ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_157_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14104__248 clknet_1_1__leaf__08494_ VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__inv_2
XFILLER_0_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19139_ clknet_leaf_15_clk _02659_ VGND VGND VPWR VPWR CPU.PC\[21\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_14_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08496_ clknet_0__08496_ VGND VGND VPWR VPWR clknet_1_1__leaf__08496_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09725_ CPU.PC\[20\] _05892_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__nor2_1
X_09656_ CPU.PC\[19\] _05924_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__nand2_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ CPU.PC\[17\] _05930_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__and2_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345__6 clknet_1_1__leaf__04984_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__inv_2
XFILLER_0_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10500_ net2418 _06054_ _06713_ VGND VGND VPWR VPWR _06714_ sky130_fd_sc_hd__mux2_1
X_11480_ _06244_ VGND VGND VPWR VPWR _07349_ sky130_fd_sc_hd__buf_4
XFILLER_0_46_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14079__225 clknet_1_1__leaf__08492_ VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__inv_2
X_10431_ _06617_ net2378 _06676_ VGND VGND VPWR VPWR _06677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13150_ net1583 _08281_ VGND VGND VPWR VPWR _08284_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10362_ _06632_ net1967 _06618_ VGND VGND VPWR VPWR _06633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12101_ _07670_ net1312 _07688_ _07691_ VGND VGND VPWR VPWR _07695_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_20_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13081_ net1369 VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__clkbuf_1
X_10293_ net1755 _06440_ _06580_ VGND VGND VPWR VPWR _06587_ sky130_fd_sc_hd__mux2_1
X_12032_ CPU.registerFile\[24\]\[18\] _07339_ _07646_ VGND VGND VPWR VPWR _07650_
+ sky130_fd_sc_hd__mux2_1
Xhold190 mapped_spi_flash.rcv_bitcount\[5\] VGND VGND VPWR VPWR net1487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16840_ CPU.registerFile\[9\]\[20\] _04460_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__or2_1
X_13739__1109 clknet_1_0__leaf__08458_ VGND VGND VPWR VPWR net1165 sky130_fd_sc_hd__inv_2
X_13860__1218 clknet_1_1__leaf__08470_ VGND VGND VPWR VPWR net1274 sky130_fd_sc_hd__inv_2
X_16771_ CPU.registerFile\[30\]\[18\] CPU.registerFile\[31\]\[18\] _04201_ VGND VGND
+ VPWR VPWR _04480_ sky130_fd_sc_hd__mux2_1
X_18510_ net331 _02034_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12934_ _06316_ net1774 _08167_ VGND VGND VPWR VPWR _08169_ sky130_fd_sc_hd__mux2_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18441_ net262 _01969_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_15653_ clknet_1_0__leaf__03643_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__buf_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ _08132_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__clkbuf_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14604_ _08837_ _08838_ _08842_ _08802_ VGND VGND VPWR VPWR _08843_ sky130_fd_sc_hd__a211o_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ net2246 _07328_ _07526_ VGND VGND VPWR VPWR _07535_ sky130_fd_sc_hd__mux2_1
X_18372_ net193 _01900_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15584_ _08557_ _03630_ _03634_ _05876_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__o211a_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12796_ _08094_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13315__815 clknet_1_0__leaf__08363_ VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__inv_2
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _08410_ VGND VGND VPWR VPWR _08776_ sky130_fd_sc_hd__clkbuf_4
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _07498_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__clkbuf_1
X_15940__678 clknet_1_0__leaf__03689_ VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__inv_2
XFILLER_0_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17254_ CPU.registerFile\[12\]\[31\] _03694_ _03763_ _04949_ VGND VGND VPWR VPWR
+ _04950_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14466_ _08581_ _08705_ _08708_ _08590_ VGND VGND VPWR VPWR _08709_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11678_ _07461_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16205_ _03758_ _03922_ _03927_ _03775_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__o211a_1
X_13417_ _08387_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__clkbuf_1
X_17185_ CPU.registerFile\[5\]\[29\] CPU.registerFile\[4\]\[29\] _03697_ VGND VGND
+ VPWR VPWR _04883_ sky130_fd_sc_hd__mux2_1
X_10629_ _06783_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14397_ CPU.registerFile\[22\]\[2\] CPU.registerFile\[23\]\[2\] _08523_ VGND VGND
+ VPWR VPWR _08641_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__08450_ _08450_ VGND VGND VPWR VPWR clknet_0__08450_ sky130_fd_sc_hd__clkbuf_16
X_16136_ CPU.registerFile\[15\]\[3\] CPU.registerFile\[14\]\[3\] _03705_ VGND VGND
+ VPWR VPWR _03860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16067_ _03722_ _03790_ _03792_ _03730_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__a211o_1
X_13279_ per_uart.uart0.enable16_counter\[15\] _08359_ VGND VGND VPWR VPWR _08360_
+ sky130_fd_sc_hd__nor2_2
XFILLER_0_110_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15018_ CPU.registerFile\[20\]\[17\] _03080_ _03081_ _03082_ VGND VGND VPWR VPWR
+ _03083_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16969_ CPU.registerFile\[5\]\[23\] CPU.registerFile\[4\]\[23\] _04428_ VGND VGND
+ VPWR VPWR _04673_ sky130_fd_sc_hd__mux2_1
X_09510_ CPU.Jimm\[13\] VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__clkbuf_4
X_18708_ net497 _02232_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[8\] sky130_fd_sc_hd__dfxtp_1
X_14110__252 clknet_1_0__leaf__08496_ VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__inv_2
X_14184__320 clknet_1_1__leaf__08502_ VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__inv_2
X_09441_ _05552_ VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18639_ clknet_leaf_15_clk _02163_ VGND VGND VPWR VPWR CPU.rs2\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09372_ _05577_ _05695_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14028__179 clknet_1_1__leaf__08487_ VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__inv_2
XFILLER_0_90_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13563__950 clknet_1_0__leaf__08441_ VGND VGND VPWR VPWR net1006 sky130_fd_sc_hd__inv_2
XFILLER_0_112_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__08479_ clknet_0__08479_ VGND VGND VPWR VPWR clknet_1_1__leaf__08479_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15616__419 clknet_1_0__leaf__03639_ VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__inv_2
X_09708_ _06003_ _05920_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__and2b_1
X_10980_ _07025_ _05605_ _05621_ VGND VGND VPWR VPWR _07026_ sky130_fd_sc_hd__o21ai_2
Xclkbuf_1_0__f__08370_ clknet_0__08370_ VGND VGND VPWR VPWR clknet_1_0__leaf__08370_
+ sky130_fd_sc_hd__clkbuf_16
X_09639_ _05981_ _05982_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__and2_1
X_12650_ _08017_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__clkbuf_1
X_11601_ _07420_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12581_ net2542 _07356_ _07979_ VGND VGND VPWR VPWR _07981_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14320_ _06058_ VGND VGND VPWR VPWR _08566_ sky130_fd_sc_hd__clkbuf_4
X_11532_ _07383_ VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11463_ net1682 _07337_ _07333_ VGND VGND VPWR VPWR _07338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13202_ _06345_ _08315_ VGND VGND VPWR VPWR _08316_ sky130_fd_sc_hd__or2_1
X_10414_ _06601_ net2373 _06665_ VGND VGND VPWR VPWR _06668_ sky130_fd_sc_hd__mux2_1
X_11394_ _07294_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13133_ CPU.cycles\[4\] _08271_ net1575 VGND VGND VPWR VPWR _08274_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10345_ _06621_ VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__clkbuf_1
X_18990_ clknet_leaf_19_clk _02510_ VGND VGND VPWR VPWR CPU.aluIn1\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ net1389 VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__clkbuf_1
X_17941_ net952 _01469_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_10276_ net1946 _06245_ _06569_ VGND VGND VPWR VPWR _06578_ sky130_fd_sc_hd__mux2_1
X_12015_ net2587 _07322_ _07635_ VGND VGND VPWR VPWR _07641_ sky130_fd_sc_hd__mux2_1
X_17872_ clknet_leaf_23_clk _00021_ VGND VGND VPWR VPWR CPU.cycles\[15\] sky130_fd_sc_hd__dfxtp_1
X_16823_ CPU.registerFile\[24\]\[19\] _04319_ _04165_ _04530_ VGND VGND VPWR VPWR
+ _04531_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16754_ _04099_ _04459_ _04462_ _04105_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__a211o_1
X_12917_ _06124_ net2487 _08156_ VGND VGND VPWR VPWR _08160_ sky130_fd_sc_hd__mux2_1
X_16685_ CPU.registerFile\[30\]\[16\] CPU.registerFile\[31\]\[16\] _04201_ VGND VGND
+ VPWR VPWR _04396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__08499_ clknet_0__08499_ VGND VGND VPWR VPWR clknet_1_0__leaf__08499_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_158_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18424_ net245 _01952_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12848_ _08123_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18355_ net176 _01883_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_15567_ _06013_ _03613_ _03617_ _08422_ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__o211a_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _08085_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__clkbuf_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14518_ CPU.registerFile\[20\]\[5\] _08527_ _08758_ _08530_ VGND VGND VPWR VPWR _08759_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15498_ CPU.registerFile\[10\]\[29\] CPU.registerFile\[11\]\[29\] _08522_ VGND VGND
+ VPWR VPWR _03551_ sky130_fd_sc_hd__mux2_1
X_18286_ net1297 _01814_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14449_ CPU.registerFile\[15\]\[3\] CPU.registerFile\[14\]\[3\] _08558_ VGND VGND
+ VPWR VPWR _08692_ sky130_fd_sc_hd__mux2_1
X_17237_ CPU.registerFile\[22\]\[30\] CPU.registerFile\[23\]\[30\] _03761_ VGND VGND
+ VPWR VPWR _04934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__08502_ _08502_ VGND VGND VPWR VPWR clknet_0__08502_ sky130_fd_sc_hd__clkbuf_16
X_17168_ CPU.registerFile\[19\]\[28\] CPU.registerFile\[18\]\[28\] _03745_ VGND VGND
+ VPWR VPWR _04867_ sky130_fd_sc_hd__mux2_1
Xhold904 CPU.registerFile\[23\]\[17\] VGND VGND VPWR VPWR net2201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 CPU.registerFile\[29\]\[12\] VGND VGND VPWR VPWR net2212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 CPU.registerFile\[26\]\[24\] VGND VGND VPWR VPWR net2223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 CPU.registerFile\[27\]\[1\] VGND VGND VPWR VPWR net2234 sky130_fd_sc_hd__dlygate4sd3_1
X_16119_ CPU.registerFile\[20\]\[2\] CPU.registerFile\[21\]\[2\] _03761_ VGND VGND
+ VPWR VPWR _03844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold948 CPU.registerFile\[23\]\[29\] VGND VGND VPWR VPWR net2245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17099_ _08397_ _04797_ _04799_ _08400_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__a211o_1
Xhold959 CPU.registerFile\[16\]\[20\] VGND VGND VPWR VPWR net2256 sky130_fd_sc_hd__dlygate4sd3_1
X_09990_ _05425_ _06319_ VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__or2_1
X_14216__349 clknet_1_1__leaf__08505_ VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__inv_2
X_13285__788 clknet_1_0__leaf__08345_ VGND VGND VPWR VPWR net844 sky130_fd_sc_hd__inv_2
XFILLER_0_110_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08941_ CPU.mem_wdata\[7\] CPU.Bimm\[7\] _05244_ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__08364_ _08364_ VGND VGND VPWR VPWR clknet_0__08364_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09424_ _05425_ _05773_ _05517_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09355_ _05705_ _05706_ _05558_ VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__a21o_1
X_15923__662 clknet_1_1__leaf__03688_ VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__inv_2
XFILLER_0_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09286_ _05558_ _05634_ _05635_ _05637_ _05235_ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__o311a_1
XFILLER_0_118_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13738__1108 clknet_1_0__leaf__08458_ VGND VGND VPWR VPWR net1164 sky130_fd_sc_hd__inv_2
XFILLER_0_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10130_ _05911_ _06451_ _06454_ VGND VGND VPWR VPWR _06455_ sky130_fd_sc_hd__o21ai_1
X_10061_ mapped_spi_ram.rcv_data\[30\] _05858_ VGND VGND VPWR VPWR _06388_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17310__724 clknet_1_0__leaf__04981_ VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__inv_2
X_13820_ clknet_1_0__leaf__08462_ VGND VGND VPWR VPWR _08467_ sky130_fd_sc_hd__buf_1
XFILLER_0_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10963_ _07001_ VGND VGND VPWR VPWR _07014_ sky130_fd_sc_hd__buf_2
XFILLER_0_97_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12702_ _06626_ net2552 _08040_ VGND VGND VPWR VPWR _08045_ sky130_fd_sc_hd__mux2_1
X_16470_ CPU.registerFile\[8\]\[11\] _04101_ _04102_ _04185_ VGND VGND VPWR VPWR _04186_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10894_ _06960_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15421_ _06013_ _03471_ _03475_ _08422_ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__o211a_1
X_12633_ _08008_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15352_ CPU.registerFile\[13\]\[25\] CPU.registerFile\[12\]\[25\] _08794_ VGND VGND
+ VPWR VPWR _03409_ sky130_fd_sc_hd__mux2_1
X_18140_ net1151 _01668_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12564_ net2492 _07339_ _07968_ VGND VGND VPWR VPWR _07972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14303_ _06035_ VGND VGND VPWR VPWR _08549_ sky130_fd_sc_hd__buf_8
X_18071_ net1082 _01599_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_11515_ net1761 _07372_ _07354_ VGND VGND VPWR VPWR _07373_ sky130_fd_sc_hd__mux2_1
X_15283_ CPU.registerFile\[8\]\[23\] _03018_ _03341_ _03268_ VGND VGND VPWR VPWR _03342_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12495_ net1741 _07339_ _07931_ VGND VGND VPWR VPWR _07935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17022_ CPU.registerFile\[20\]\[24\] CPU.registerFile\[21\]\[24\] _03737_ VGND VGND
+ VPWR VPWR _04725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11446_ _05872_ VGND VGND VPWR VPWR _07326_ sky130_fd_sc_hd__buf_4
XFILLER_0_150_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__03691_ _03691_ VGND VGND VPWR VPWR clknet_0__03691_ sky130_fd_sc_hd__clkbuf_16
X_11377_ net1826 _06054_ _07285_ VGND VGND VPWR VPWR _07286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13116_ _05236_ _08264_ VGND VGND VPWR VPWR _08265_ sky130_fd_sc_hd__nor2_1
X_10328_ _06609_ net1929 _06597_ VGND VGND VPWR VPWR _06610_ sky130_fd_sc_hd__mux2_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18973_ net747 _02493_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ net2497 _06053_ _08228_ VGND VGND VPWR VPWR _08229_ sky130_fd_sc_hd__mux2_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ clknet_leaf_2_clk _01452_ VGND VGND VPWR VPWR CPU.Bimm\[12\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_56_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10259_ _06557_ VGND VGND VPWR VPWR _06569_ sky130_fd_sc_hd__buf_4
X_17855_ net935 _01417_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_16806_ _04419_ _04511_ _04513_ _04383_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__a211o_1
X_17786_ net866 _01348_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14998_ CPU.registerFile\[6\]\[16\] CPU.registerFile\[7\]\[16\] _02982_ VGND VGND
+ VPWR VPWR _03064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16737_ _04075_ _04440_ _04445_ _04446_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16668_ CPU.registerFile\[15\]\[16\] CPU.registerFile\[14\]\[16\] _04146_ VGND VGND
+ VPWR VPWR _04379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18407_ net228 _01935_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_15619_ clknet_1_0__leaf__08506_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__buf_1
X_15645__445 clknet_1_0__leaf__03642_ VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__inv_2
X_16599_ _03943_ _04309_ _04311_ _04117_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09140_ _05488_ _05490_ _05491_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18338_ net159 _01866_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14222__353 clknet_1_1__leaf__08507_ VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__inv_2
XFILLER_0_84_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09071_ CPU.Bimm\[10\] _05422_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__nand2_1
X_18269_ net1280 _01797_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold701 CPU.registerFile\[7\]\[25\] VGND VGND VPWR VPWR net1998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold712 CPU.registerFile\[28\]\[17\] VGND VGND VPWR VPWR net2009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 CPU.registerFile\[15\]\[5\] VGND VGND VPWR VPWR net2020 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold734 CPU.registerFile\[16\]\[24\] VGND VGND VPWR VPWR net2031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 CPU.registerFile\[29\]\[23\] VGND VGND VPWR VPWR net2042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 CPU.registerFile\[11\]\[21\] VGND VGND VPWR VPWR net2053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 CPU.registerFile\[30\]\[22\] VGND VGND VPWR VPWR net2064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold778 CPU.registerFile\[17\]\[25\] VGND VGND VPWR VPWR net2075 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ _05514_ _05310_ _06202_ _06301_ _06303_ VGND VGND VPWR VPWR _06304_ sky130_fd_sc_hd__a311o_4
Xhold789 CPU.registerFile\[30\]\[30\] VGND VGND VPWR VPWR net2086 sky130_fd_sc_hd__dlygate4sd3_1
X_08924_ CPU.Iimm\[0\] _05248_ _05275_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__o21a_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03680_ clknet_0__03680_ VGND VGND VPWR VPWR clknet_1_0__leaf__03680_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09407_ _05549_ VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09338_ mapped_spi_ram.rcv_data\[23\] _05683_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__nand2_8
XFILLER_0_8_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09269_ _05618_ _05602_ _05619_ _05620_ _05595_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__a311oi_2
XFILLER_0_133_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11300_ net1752 _05853_ _07238_ VGND VGND VPWR VPWR _07245_ sky130_fd_sc_hd__mux2_1
X_12280_ mapped_spi_ram.rcv_data\[10\] _07813_ VGND VGND VPWR VPWR _07815_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11231_ _06609_ net1757 _07201_ VGND VGND VPWR VPWR _07208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11162_ net1926 _07160_ _07162_ _07164_ VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__o211a_1
X_10113_ _06176_ net1367 _06426_ _06438_ VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__a211o_2
X_15970_ _03696_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__buf_4
X_11093_ mapped_spi_flash.snd_bitcount\[3\] _07119_ _07120_ VGND VGND VPWR VPWR _07121_
+ sky130_fd_sc_hd__o21ba_1
X_15750__540 clknet_1_1__leaf__03652_ VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__inv_2
X_13895__59 clknet_1_1__leaf__08474_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__inv_2
X_14921_ _08785_ _02986_ _02988_ _08870_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__a211o_1
X_10044_ _05448_ _06371_ _05424_ VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__a21o_1
Xhold50 _05766_ VGND VGND VPWR VPWR net1347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold61 mapped_spi_ram.state\[3\] VGND VGND VPWR VPWR net1358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 _08246_ VGND VGND VPWR VPWR net1369 sky130_fd_sc_hd__dlygate4sd3_1
X_17640_ _05179_ net1659 _05180_ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__a21oi_1
Xhold83 _08225_ VGND VGND VPWR VPWR net1380 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14852_ CPU.registerFile\[21\]\[13\] _08718_ VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__or2_1
Xhold94 _06464_ VGND VGND VPWR VPWR net1391 sky130_fd_sc_hd__dlygate4sd3_1
X_14783_ _08808_ _08809_ CPU.registerFile\[25\]\[11\] VGND VGND VPWR VPWR _02854_
+ sky130_fd_sc_hd__a21o_1
X_17571_ per_uart.uart0.tx_count16\[1\] _03659_ _05134_ VGND VGND VPWR VPWR _05135_
+ sky130_fd_sc_hd__and3_1
X_11995_ _07629_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__clkbuf_1
X_16522_ _03901_ _04231_ _04236_ _04072_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__o211a_1
X_10946_ _07001_ VGND VGND VPWR VPWR _07002_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13665_ clknet_1_0__leaf__08451_ VGND VGND VPWR VPWR _08452_ sky130_fd_sc_hd__buf_1
X_16453_ _03757_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__clkbuf_4
X_10877_ CPU.aluReg\[8\] _06947_ _06922_ VGND VGND VPWR VPWR _06948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12616_ _07999_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__clkbuf_1
X_15404_ _03155_ _03442_ _03459_ _03243_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__a211o_2
XFILLER_0_27_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16384_ _06149_ VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__clkbuf_4
X_19172_ clknet_leaf_5_clk _02692_ VGND VGND VPWR VPWR per_uart.uart0.rx_count16\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18123_ net1134 _01651_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_15335_ CPU.registerFile\[17\]\[25\] _03036_ VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__or2_1
X_12547_ net2362 _07322_ _07957_ VGND VGND VPWR VPWR _07963_ sky130_fd_sc_hd__mux2_1
X_18054_ net1065 _01582_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_15266_ CPU.registerFile\[21\]\[23\] _02960_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__or2_1
X_12478_ net2291 _07322_ _07920_ VGND VGND VPWR VPWR _07926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_3 CPU.mem_wdata\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17005_ CPU.registerFile\[5\]\[24\] CPU.registerFile\[4\]\[24\] _04428_ VGND VGND
+ VPWR VPWR _04708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11429_ net1751 _07314_ _07312_ VGND VGND VPWR VPWR _07315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15197_ _03049_ _03050_ CPU.registerFile\[25\]\[21\] VGND VGND VPWR VPWR _03258_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03643_ clknet_0__03643_ VGND VGND VPWR VPWR clknet_1_1__leaf__03643_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_22_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18956_ net730 _02476_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17907_ clknet_leaf_22_clk _01435_ VGND VGND VPWR VPWR CPU.Jimm\[14\] sky130_fd_sc_hd__dfxtp_2
X_18887_ net661 _02407_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_13737__1107 clknet_1_1__leaf__08458_ VGND VGND VPWR VPWR net1163 sky130_fd_sc_hd__inv_2
X_17838_ net918 _01400_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17769_ net849 _01331_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[9\] sky130_fd_sc_hd__dfxtp_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17395__19 clknet_1_1__leaf__04985_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__inv_2
XFILLER_0_119_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09123_ CPU.aluIn1\[17\] _05345_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09054_ _05393_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold520 CPU.registerFile\[6\]\[15\] VGND VGND VPWR VPWR net1817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 CPU.registerFile\[28\]\[28\] VGND VGND VPWR VPWR net1828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold542 CPU.registerFile\[13\]\[10\] VGND VGND VPWR VPWR net1839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold553 CPU.registerFile\[19\]\[20\] VGND VGND VPWR VPWR net1850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 CPU.registerFile\[15\]\[3\] VGND VGND VPWR VPWR net1861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold575 CPU.registerFile\[19\]\[3\] VGND VGND VPWR VPWR net1872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 CPU.registerFile\[21\]\[7\] VGND VGND VPWR VPWR net1883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 _05172_ VGND VGND VPWR VPWR net1894 sky130_fd_sc_hd__dlygate4sd3_1
X_09956_ _05693_ _05822_ VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__or2_1
X_13599__982 clknet_1_1__leaf__08445_ VGND VGND VPWR VPWR net1038 sky130_fd_sc_hd__inv_2
X_08907_ _05256_ _05258_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__nor2_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _05911_ _06219_ _06221_ _06197_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__o22a_1
Xhold1220 CPU.registerFile\[26\]\[15\] VGND VGND VPWR VPWR net2517 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1231 CPU.registerFile\[7\]\[30\] VGND VGND VPWR VPWR net2528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1242 CPU.registerFile\[21\]\[18\] VGND VGND VPWR VPWR net2539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1253 CPU.registerFile\[25\]\[15\] VGND VGND VPWR VPWR net2550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1264 CPU.registerFile\[26\]\[3\] VGND VGND VPWR VPWR net2561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 CPU.registerFile\[1\]\[0\] VGND VGND VPWR VPWR net2572 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1286 CPU.registerFile\[9\]\[13\] VGND VGND VPWR VPWR net2583 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1297 CPU.registerFile\[9\]\[4\] VGND VGND VPWR VPWR net2594 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _06868_ VGND VGND VPWR VPWR _06889_ sky130_fd_sc_hd__clkbuf_4
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _06645_ net2134 _07512_ VGND VGND VPWR VPWR _07516_ sky130_fd_sc_hd__mux2_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10731_ net2269 _06292_ _06838_ VGND VGND VPWR VPWR _06839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15780__566 clknet_1_1__leaf__03656_ VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__inv_2
X_13450_ _08410_ VGND VGND VPWR VPWR _08411_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10662_ net2436 _06316_ _06799_ VGND VGND VPWR VPWR _06801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12401_ _07885_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10593_ _06763_ VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__clkbuf_1
X_13659__1037 clknet_1_0__leaf__08450_ VGND VGND VPWR VPWR net1093 sky130_fd_sc_hd__inv_2
X_15120_ _08525_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__buf_4
XFILLER_0_91_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12332_ _06593_ net1843 _07848_ VGND VGND VPWR VPWR _07849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15051_ net1656 _02797_ _03115_ _02993_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__o211a_1
X_12263_ mapped_spi_ram.rcv_data\[17\] _07800_ VGND VGND VPWR VPWR _07805_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11214_ mapped_spi_flash.div_counter\[1\] _07176_ VGND VGND VPWR VPWR _07198_ sky130_fd_sc_hd__nor2_1
Xoutput5 net5 VGND VGND VPWR VPWR LEDS sky130_fd_sc_hd__clkbuf_4
X_12194_ CPU.mem_wdata\[0\] _07680_ _07696_ _07694_ VGND VGND VPWR VPWR _07757_ sky130_fd_sc_hd__a211o_1
X_18810_ net599 _02334_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_17316__730 clknet_1_1__leaf__04981_ VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__inv_2
X_11145_ net1384 _07147_ _07154_ _07151_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__o211a_1
X_15674__471 clknet_1_1__leaf__03645_ VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__inv_2
X_18741_ net530 _02265_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[3\] sky130_fd_sc_hd__dfxtp_1
X_11076_ _07107_ VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__04979_ clknet_0__04979_ VGND VGND VPWR VPWR clknet_1_0__leaf__04979_
+ sky130_fd_sc_hd__clkbuf_16
X_10027_ CPU.PC\[8\] _05884_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__nor2_1
X_14904_ _02964_ _02967_ _02971_ _08851_ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__o211a_1
X_18672_ net461 _02196_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_17623_ net1668 VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__clkbuf_1
X_14835_ _02728_ _02899_ _02904_ _02784_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17554_ net2199 VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__inv_2
X_14766_ _02825_ _02836_ _02837_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__o21a_2
X_11978_ _06638_ net2569 _07620_ VGND VGND VPWR VPWR _07621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16505_ CPU.aluIn1\[11\] _04054_ _04220_ _03855_ VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__o211a_1
X_10929_ _06989_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__clkbuf_1
X_14697_ _08808_ _08809_ CPU.registerFile\[25\]\[9\] VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__a21o_1
X_17485_ _08379_ _05017_ _06263_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_160_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13511__903 clknet_1_0__leaf__08436_ VGND VGND VPWR VPWR net959 sky130_fd_sc_hd__inv_2
XFILLER_0_129_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16436_ _06534_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19155_ clknet_leaf_3_clk net1533 VGND VGND VPWR VPWR per_uart.uart0.txd_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16367_ CPU.registerFile\[22\]\[8\] CPU.registerFile\[23\]\[8\] _03958_ VGND VGND
+ VPWR VPWR _04086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18106_ net1117 _01634_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_15318_ _03138_ _03139_ CPU.registerFile\[9\]\[24\] VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__a21o_1
X_16298_ _06149_ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__clkbuf_4
X_19086_ clknet_leaf_0_clk _02606_ VGND VGND VPWR VPWR per_uart.uart0.rxd_reg\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18037_ net1048 _01565_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15249_ _03133_ _03303_ _03308_ _03188_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__o211a_1
X_15757__546 clknet_1_0__leaf__03653_ VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__inv_2
XFILLER_0_140_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09810_ mapped_spi_ram.rcv_data\[8\] _05685_ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09741_ _05764_ _06065_ _06078_ _06081_ VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__a211o_4
X_18939_ net713 _02459_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_09672_ CPU.PC\[21\] _05893_ CPU.PC\[22\] VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_19_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09106_ _05328_ _05333_ _05319_ _05457_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__and4_1
XFILLER_0_21_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09037_ CPU.aluIn1\[24\] _05387_ VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold350 CPU.rs2\[15\] VGND VGND VPWR VPWR net1647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold361 CPU.registerFile\[31\]\[24\] VGND VGND VPWR VPWR net1658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 mapped_spi_flash.state\[1\] VGND VGND VPWR VPWR net1669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 CPU.registerFile\[5\]\[31\] VGND VGND VPWR VPWR net1680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 CPU.registerFile\[5\]\[0\] VGND VGND VPWR VPWR net1691 sky130_fd_sc_hd__dlygate4sd3_1
X_09939_ _05428_ _05448_ _05449_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__a21o_1
X_12950_ _06508_ net2507 _08167_ VGND VGND VPWR VPWR _08177_ sky130_fd_sc_hd__mux2_1
Xhold1050 CPU.registerFile\[16\]\[26\] VGND VGND VPWR VPWR net2347 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ _06630_ net1854 _07573_ VGND VGND VPWR VPWR _07580_ sky130_fd_sc_hd__mux2_1
Xhold1061 CPU.registerFile\[29\]\[20\] VGND VGND VPWR VPWR net2358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 CPU.registerFile\[23\]\[27\] VGND VGND VPWR VPWR net2369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 CPU.registerFile\[5\]\[8\] VGND VGND VPWR VPWR net2380 sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ _08140_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__clkbuf_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1094 CPU.registerFile\[22\]\[1\] VGND VGND VPWR VPWR net2391 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _08567_ _08569_ CPU.registerFile\[9\]\[7\] VGND VGND VPWR VPWR _08859_ sky130_fd_sc_hd__a21o_1
X_11832_ _07543_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__clkbuf_1
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03646_ clknet_0__03646_ VGND VGND VPWR VPWR clknet_1_0__leaf__03646_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14551_ _08425_ _08770_ _08791_ _08597_ VGND VGND VPWR VPWR _08792_ sky130_fd_sc_hd__a211o_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _06628_ net1966 _07501_ VGND VGND VPWR VPWR _07507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ net1831 _06106_ _06827_ VGND VGND VPWR VPWR _06830_ sky130_fd_sc_hd__mux2_1
X_17270_ CPU.registerFile\[24\]\[31\] _03724_ _03725_ _04965_ VGND VGND VPWR VPWR
+ _04966_ sky130_fd_sc_hd__o211a_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ CPU.registerFile\[28\]\[4\] CPU.registerFile\[29\]\[4\] _08538_ VGND VGND
+ VPWR VPWR _08724_ sky130_fd_sc_hd__mux2_1
X_11694_ net2140 _07343_ _07464_ VGND VGND VPWR VPWR _07470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13433_ _08397_ VGND VGND VPWR VPWR _08398_ sky130_fd_sc_hd__buf_4
X_16221_ _08396_ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10645_ net2611 _06124_ _06788_ VGND VGND VPWR VPWR _06792_ sky130_fd_sc_hd__mux2_1
X_16152_ _03873_ _03874_ _03875_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__mux2_1
X_13736__1106 clknet_1_1__leaf__08458_ VGND VGND VPWR VPWR net1162 sky130_fd_sc_hd__inv_2
XFILLER_0_122_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10576_ _06754_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__clkbuf_1
X_12315_ net1298 _07781_ net1303 VGND VGND VPWR VPWR _07837_ sky130_fd_sc_hd__a21o_1
X_15103_ CPU.registerFile\[21\]\[19\] _02960_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__or2_1
X_16083_ CPU.registerFile\[19\]\[1\] CPU.registerFile\[18\]\[1\] _03767_ VGND VGND
+ VPWR VPWR _03809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14056__204 clknet_1_0__leaf__08490_ VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__inv_2
X_15034_ CPU.registerFile\[10\]\[17\] CPU.registerFile\[11\]\[17\] _02779_ VGND VGND
+ VPWR VPWR _03099_ sky130_fd_sc_hd__mux2_1
X_12246_ net1523 _07787_ VGND VGND VPWR VPWR _07795_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12177_ net1467 _07738_ _07747_ _07737_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__o211a_1
X_11128_ net1540 _07133_ _07144_ _07138_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__o211a_1
X_16985_ CPU.registerFile\[22\]\[23\] CPU.registerFile\[23\]\[23\] _04362_ VGND VGND
+ VPWR VPWR _04689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18724_ net513 _02248_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[24\] sky130_fd_sc_hd__dfxtp_1
X_11059_ _05591_ _07094_ _05590_ VGND VGND VPWR VPWR _07095_ sky130_fd_sc_hd__a21oi_1
X_18655_ clknet_leaf_12_clk _02179_ VGND VGND VPWR VPWR CPU.rs2\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17606_ per_uart.d_in_uart\[2\] _05134_ _05157_ net1474 VGND VGND VPWR VPWR _05161_
+ sky130_fd_sc_hd__o22a_1
X_14818_ CPU.registerFile\[30\]\[12\] CPU.registerFile\[31\]\[12\] _02887_ VGND VGND
+ VPWR VPWR _02888_ sky130_fd_sc_hd__mux2_1
X_18586_ net407 net43 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_15798_ _08350_ _03667_ _03661_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__a21oi_1
X_17537_ _05069_ CPU.PC\[21\] _05106_ _05107_ _06858_ VGND VGND VPWR VPWR _02659_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_157_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14749_ CPU.registerFile\[10\]\[10\] CPU.registerFile\[11\]\[10\] _02779_ VGND VGND
+ VPWR VPWR _02821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17468_ _05049_ _05050_ _05020_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16419_ _03758_ _04132_ _04136_ _03775_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19138_ clknet_leaf_15_clk _02658_ VGND VGND VPWR VPWR CPU.PC\[20\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19069_ net61 _02589_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[22\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_8_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__08495_ clknet_0__08495_ VGND VGND VPWR VPWR clknet_1_1__leaf__08495_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09724_ _05856_ _06064_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__nand2_1
X_13658__1036 clknet_1_0__leaf__08450_ VGND VGND VPWR VPWR net1092 sky130_fd_sc_hd__inv_2
X_09655_ _05997_ _05998_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09586_ CPU.Jimm\[17\] _05921_ _05923_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__a21o_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10430_ _06664_ VGND VGND VPWR VPWR _06676_ sky130_fd_sc_hd__buf_4
XFILLER_0_73_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14005__158 clknet_1_0__leaf__08485_ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__inv_2
XFILLER_0_162_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10361_ _06223_ VGND VGND VPWR VPWR _06632_ sky130_fd_sc_hd__buf_4
XFILLER_0_115_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12100_ net1312 VGND VGND VPWR VPWR _07694_ sky130_fd_sc_hd__clkbuf_4
X_13080_ CPU.registerFile\[4\]\[5\] net1368 _08239_ VGND VGND VPWR VPWR _08246_ sky130_fd_sc_hd__mux2_1
X_10292_ _06586_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__clkbuf_1
X_12031_ _07649_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__clkbuf_1
Xhold180 _02677_ VGND VGND VPWR VPWR net1477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 _07129_ VGND VGND VPWR VPWR net1488 sky130_fd_sc_hd__dlygate4sd3_1
X_16770_ _03713_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__clkbuf_4
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ _08168_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__clkbuf_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ net261 _01968_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ clknet_1_1__leaf__08339_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__buf_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _06292_ net2145 _08131_ VGND VGND VPWR VPWR _08132_ sky130_fd_sc_hd__mux2_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ CPU.registerFile\[20\]\[7\] _08839_ _08840_ _08841_ VGND VGND VPWR VPWR _08842_
+ sky130_fd_sc_hd__o211a_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _07534_ VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__clkbuf_1
X_18371_ net192 _01899_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15583_ _08414_ _03631_ _03633_ _08419_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__a211o_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _06651_ net2504 _08087_ VGND VGND VPWR VPWR _08094_ sky130_fd_sc_hd__mux2_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14534_ CPU.registerFile\[10\]\[5\] CPU.registerFile\[11\]\[5\] _08564_ VGND VGND
+ VPWR VPWR _08775_ sky130_fd_sc_hd__mux2_1
X_11746_ _06611_ net2394 _07490_ VGND VGND VPWR VPWR _07498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17253_ CPU.registerFile\[13\]\[31\] _03767_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11677_ net2509 _07326_ _07453_ VGND VGND VPWR VPWR _07461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14465_ CPU.registerFile\[0\]\[3\] _08706_ _08707_ _08588_ VGND VGND VPWR VPWR _08708_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16204_ _03766_ _03924_ _03926_ _06142_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__a211o_1
X_10628_ net2580 _05839_ _06777_ VGND VGND VPWR VPWR _06783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13416_ _05737_ _06311_ _00000_ VGND VGND VPWR VPWR _08387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17184_ CPU.registerFile\[6\]\[29\] CPU.registerFile\[7\]\[29\] _03847_ VGND VGND
+ VPWR VPWR _04882_ sky130_fd_sc_hd__mux2_1
X_14396_ _08415_ _08637_ _08639_ _08420_ VGND VGND VPWR VPWR _08640_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16135_ _08398_ _03856_ _03858_ _08401_ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10559_ _06745_ VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16066_ CPU.registerFile\[0\]\[1\] _03724_ _03725_ _03791_ VGND VGND VPWR VPWR _03792_
+ sky130_fd_sc_hd__o211a_1
X_13278_ per_uart.uart0.enable16_counter\[14\] _08358_ VGND VGND VPWR VPWR _08359_
+ sky130_fd_sc_hd__or2_1
X_12229_ _07784_ VGND VGND VPWR VPWR _07785_ sky130_fd_sc_hd__buf_2
X_15017_ _06036_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__clkbuf_4
X_15869__614 clknet_1_0__leaf__03682_ VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__inv_2
X_16968_ CPU.registerFile\[6\]\[23\] CPU.registerFile\[7\]\[23\] _04426_ VGND VGND
+ VPWR VPWR _04672_ sky130_fd_sc_hd__mux2_1
X_18707_ net496 _02231_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[7\] sky130_fd_sc_hd__dfxtp_1
X_16899_ _03736_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__buf_4
X_09440_ _05556_ _05788_ _05731_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__o21a_1
XFILLER_0_91_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18638_ clknet_leaf_15_clk _02162_ VGND VGND VPWR VPWR CPU.rs2\[10\] sky130_fd_sc_hd__dfxtp_1
X_13967__124 clknet_1_1__leaf__08481_ VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__inv_2
XFILLER_0_59_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09371_ mapped_spi_ram.rcv_data\[15\] _05683_ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__nand2_2
XFILLER_0_93_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18569_ net390 net26 VGND VGND VPWR VPWR CPU.registerFile\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__08478_ clknet_0__08478_ VGND VGND VPWR VPWR clknet_1_1__leaf__08478_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13930__91 clknet_1_1__leaf__08477_ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__inv_2
X_09707_ CPU.Iimm\[1\] _05758_ _05790_ CPU.cycles\[21\] _06048_ VGND VGND VPWR VPWR
+ _06049_ sky130_fd_sc_hd__a221o_1
X_13735__1105 clknet_1_1__leaf__08458_ VGND VGND VPWR VPWR net1161 sky130_fd_sc_hd__inv_2
X_09638_ CPU.PC\[14\] _05980_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__or2_1
X_09569_ _05547_ CPU.instr\[4\] VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__nand2b_2
X_11600_ net2219 _07318_ _07416_ VGND VGND VPWR VPWR _07420_ sky130_fd_sc_hd__mux2_1
X_12580_ _07980_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__clkbuf_1
X_11531_ net2294 _07318_ _07379_ VGND VGND VPWR VPWR _07383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11462_ _06105_ VGND VGND VPWR VPWR _07337_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13201_ _05300_ _05443_ _08313_ _08314_ VGND VGND VPWR VPWR _08315_ sky130_fd_sc_hd__or4_1
XFILLER_0_135_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10413_ _06667_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__05015_ clknet_0__05015_ VGND VGND VPWR VPWR clknet_1_0__leaf__05015_
+ sky130_fd_sc_hd__clkbuf_16
X_11393_ net1795 _06245_ _07285_ VGND VGND VPWR VPWR _07294_ sky130_fd_sc_hd__mux2_1
X_13132_ net2666 CPU.cycles\[5\] _08271_ VGND VGND VPWR VPWR _08273_ sky130_fd_sc_hd__and3_1
X_10344_ _06620_ net1847 _06618_ VGND VGND VPWR VPWR _06621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ CPU.registerFile\[4\]\[13\] net1388 _08228_ VGND VGND VPWR VPWR _08237_ sky130_fd_sc_hd__mux2_1
X_17940_ net951 _01468_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_10275_ _06577_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__clkbuf_1
X_12014_ _07640_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__clkbuf_1
X_17871_ clknet_leaf_24_clk _00020_ VGND VGND VPWR VPWR CPU.cycles\[14\] sky130_fd_sc_hd__dfxtp_1
X_16822_ _04484_ _04485_ CPU.registerFile\[25\]\[19\] VGND VGND VPWR VPWR _04530_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14168__305 clknet_1_0__leaf__08501_ VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__inv_2
X_16753_ CPU.registerFile\[8\]\[18\] _04101_ _04102_ _04461_ VGND VGND VPWR VPWR _04462_
+ sky130_fd_sc_hd__o211a_1
X_12916_ _08159_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__clkbuf_1
X_16684_ _04098_ _04378_ _04384_ _04394_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__a31o_2
XFILLER_0_158_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__08498_ clknet_0__08498_ VGND VGND VPWR VPWR clknet_1_0__leaf__08498_
+ sky130_fd_sc_hd__clkbuf_16
X_18423_ net244 _01951_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _06106_ net2332 _08120_ VGND VGND VPWR VPWR _08123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ net175 _01882_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_15566_ _08580_ _03614_ _03616_ _08418_ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__a211o_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _06634_ net2454 _08076_ VGND VGND VPWR VPWR _08085_ sky130_fd_sc_hd__mux2_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14517_ CPU.registerFile\[21\]\[5\] _08718_ VGND VGND VPWR VPWR _08758_ sky130_fd_sc_hd__or2_1
X_11729_ _05735_ _05736_ CPU.writeBack VGND VGND VPWR VPWR _07488_ sky130_fd_sc_hd__and3b_4
X_18285_ net1296 _01813_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15497_ _03548_ _03549_ _08541_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17236_ _03714_ _04928_ _04932_ _08403_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14448_ _08515_ _08677_ _08681_ _08690_ VGND VGND VPWR VPWR _08691_ sky130_fd_sc_hd__a31o_1
Xclkbuf_0__08501_ _08501_ VGND VGND VPWR VPWR clknet_0__08501_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_40_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13657__1035 clknet_1_0__leaf__08450_ VGND VGND VPWR VPWR net1091 sky130_fd_sc_hd__inv_2
XFILLER_0_101_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17167_ _04864_ _04865_ _03742_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14379_ _08520_ _08620_ _08623_ _08419_ VGND VGND VPWR VPWR _08624_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold905 CPU.registerFile\[21\]\[31\] VGND VGND VPWR VPWR net2202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 CPU.registerFile\[29\]\[5\] VGND VGND VPWR VPWR net2213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 CPU.registerFile\[20\]\[13\] VGND VGND VPWR VPWR net2224 sky130_fd_sc_hd__dlygate4sd3_1
X_16118_ CPU.registerFile\[22\]\[2\] CPU.registerFile\[23\]\[2\] _03759_ VGND VGND
+ VPWR VPWR _03843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold938 CPU.registerFile\[27\]\[16\] VGND VGND VPWR VPWR net2235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 CPU.registerFile\[9\]\[23\] VGND VGND VPWR VPWR net2246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17098_ CPU.registerFile\[16\]\[26\] _04656_ _04494_ _04798_ VGND VGND VPWR VPWR
+ _04799_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__08363_ _08363_ VGND VGND VPWR VPWR clknet_0__08363_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16049_ _03758_ _03764_ _03774_ _03775_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__o211a_1
X_08940_ _05269_ _05283_ _05286_ _05290_ _05291_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_86_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14034__184 clknet_1_0__leaf__08488_ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__inv_2
XFILLER_0_79_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13593__977 clknet_1_1__leaf__08444_ VGND VGND VPWR VPWR net1033 sky130_fd_sc_hd__inv_2
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09423_ _05408_ _05772_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09354_ _05585_ _05589_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09285_ CPU.PC\[21\] _05636_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15622__424 clknet_1_1__leaf__03640_ VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__inv_2
XFILLER_0_31_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14117__259 clknet_1_1__leaf__08496_ VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__inv_2
X_10060_ _06387_ VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10962_ _07008_ _07012_ VGND VGND VPWR VPWR _07013_ sky130_fd_sc_hd__or2_1
X_12701_ _08044_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__clkbuf_1
X_10893_ net2633 _06959_ _06868_ VGND VGND VPWR VPWR _06960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15420_ _08580_ _03472_ _03474_ _03218_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__a211o_1
X_13717__1089 clknet_1_1__leaf__08456_ VGND VGND VPWR VPWR net1145 sky130_fd_sc_hd__inv_2
X_12632_ _06624_ net1956 _08004_ VGND VGND VPWR VPWR _08008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15351_ CPU.registerFile\[15\]\[25\] CPU.registerFile\[14\]\[25\] _08560_ VGND VGND
+ VPWR VPWR _03408_ sky130_fd_sc_hd__mux2_1
X_12563_ _07971_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11514_ _06507_ VGND VGND VPWR VPWR _07372_ sky130_fd_sc_hd__clkbuf_4
X_14302_ _08546_ _08547_ CPU.registerFile\[25\]\[0\] VGND VGND VPWR VPWR _08548_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18070_ net1081 _01598_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12494_ _07934_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__clkbuf_1
X_15282_ _03138_ _03139_ CPU.registerFile\[9\]\[23\] VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17021_ CPU.registerFile\[22\]\[24\] CPU.registerFile\[23\]\[24\] _04362_ VGND VGND
+ VPWR VPWR _04724_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11445_ _07325_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__03690_ _03690_ VGND VGND VPWR VPWR clknet_0__03690_ sky130_fd_sc_hd__clkbuf_16
X_14164_ clknet_1_1__leaf__08495_ VGND VGND VPWR VPWR _08501_ sky130_fd_sc_hd__buf_1
XFILLER_0_151_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11376_ _07273_ VGND VGND VPWR VPWR _07285_ sky130_fd_sc_hd__buf_4
XFILLER_0_150_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10327_ _05852_ VGND VGND VPWR VPWR _06609_ sky130_fd_sc_hd__clkbuf_4
X_13115_ CPU.state\[2\] _08252_ VGND VGND VPWR VPWR _08264_ sky130_fd_sc_hd__nand2_1
X_18972_ net746 _02492_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _08216_ VGND VGND VPWR VPWR _08228_ sky130_fd_sc_hd__buf_4
X_17923_ clknet_leaf_23_clk _01451_ VGND VGND VPWR VPWR CPU.Bimm\[10\] sky130_fd_sc_hd__dfxtp_4
X_10258_ _06568_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__clkbuf_1
X_17854_ net934 _01416_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_10189_ _06140_ _06510_ _05724_ VGND VGND VPWR VPWR _06511_ sky130_fd_sc_hd__mux2_1
X_16805_ CPU.registerFile\[12\]\[19\] _04421_ _04422_ _04512_ VGND VGND VPWR VPWR
+ _04513_ sky130_fd_sc_hd__o211a_1
X_17785_ net865 _01347_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_18589__46 VGND VGND VPWR VPWR _18589__46/HI net46 sky130_fd_sc_hd__conb_1
X_14997_ _02728_ _03058_ _03062_ _02784_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__o211a_1
X_16736_ _06495_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__buf_4
XFILLER_0_158_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16667_ _04099_ _04375_ _04377_ _04105_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__a211o_1
XFILLER_0_159_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18406_ net227 _01934_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16598_ CPU.registerFile\[0\]\[14\] _04233_ _04068_ _04310_ VGND VGND VPWR VPWR _04311_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18337_ net158 _01865_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15549_ _08596_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_155_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13291__793 clknet_1_0__leaf__08361_ VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__inv_2
XFILLER_0_56_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09070_ CPU.instr\[5\] VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18268_ net1279 _01796_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17219_ _03766_ _04913_ _04915_ _03716_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__a211o_1
X_18199_ net1210 _01727_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold702 CPU.registerFile\[10\]\[15\] VGND VGND VPWR VPWR net1999 sky130_fd_sc_hd__dlygate4sd3_1
X_13734__1104 clknet_1_1__leaf__08458_ VGND VGND VPWR VPWR net1160 sky130_fd_sc_hd__inv_2
Xhold713 CPU.registerFile\[18\]\[24\] VGND VGND VPWR VPWR net2010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold724 CPU.registerFile\[15\]\[28\] VGND VGND VPWR VPWR net2021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 CPU.registerFile\[22\]\[2\] VGND VGND VPWR VPWR net2032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 CPU.registerFile\[3\]\[20\] VGND VGND VPWR VPWR net2043 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold757 CPU.registerFile\[18\]\[21\] VGND VGND VPWR VPWR net2054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 CPU.registerFile\[11\]\[17\] VGND VGND VPWR VPWR net2065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold779 CPU.registerFile\[5\]\[22\] VGND VGND VPWR VPWR net2076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09972_ _05261_ _05533_ _05536_ CPU.aluReg\[10\] _06302_ VGND VGND VPWR VPWR _06303_
+ sky130_fd_sc_hd__a221o_1
X_08923_ _05240_ _05241_ CPU.mem_wdata\[0\] _05243_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__a211o_1
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13601__984 clknet_1_0__leaf__08445_ VGND VGND VPWR VPWR net1040 sky130_fd_sc_hd__inv_2
XFILLER_0_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15847__594 clknet_1_0__leaf__03680_ VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__inv_2
X_13374__868 clknet_1_1__leaf__08369_ VGND VGND VPWR VPWR net924 sky130_fd_sc_hd__inv_2
XFILLER_0_138_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09406_ _05750_ _05751_ _05756_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__or3_2
XFILLER_0_48_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09337_ _05659_ _05678_ _05688_ _05683_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__a211o_4
XFILLER_0_118_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09268_ _05596_ _05597_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__and2b_1
XFILLER_0_161_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09199_ _05547_ CPU.instr\[2\] VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11230_ _07207_ VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11161_ _07163_ VGND VGND VPWR VPWR _07164_ sky130_fd_sc_hd__buf_2
X_10112_ _06434_ _06435_ _06437_ _05541_ VGND VGND VPWR VPWR _06438_ sky130_fd_sc_hd__o31a_1
X_11092_ net1669 _07114_ VGND VGND VPWR VPWR _07120_ sky130_fd_sc_hd__nor2_1
X_14920_ CPU.registerFile\[0\]\[14\] _02948_ _02987_ _02791_ VGND VGND VPWR VPWR _02988_
+ sky130_fd_sc_hd__o211a_1
X_10043_ _05296_ _05429_ _05447_ VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__nand3b_1
X_15592__397 clknet_1_1__leaf__08511_ VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__inv_2
Xhold40 mapped_spi_ram.snd_bitcount\[3\] VGND VGND VPWR VPWR net1337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 _08219_ VGND VGND VPWR VPWR net1348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 _08251_ VGND VGND VPWR VPWR net1359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 mapped_spi_flash.rcv_data\[19\] VGND VGND VPWR VPWR net1370 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ CPU.registerFile\[22\]\[13\] CPU.registerFile\[23\]\[13\] _08756_ VGND VGND
+ VPWR VPWR _02920_ sky130_fd_sc_hd__mux2_1
Xhold84 mapped_spi_flash.rcv_data\[5\] VGND VGND VPWR VPWR net1381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 _08247_ VGND VGND VPWR VPWR net1392 sky130_fd_sc_hd__dlygate4sd3_1
X_13656__1034 clknet_1_0__leaf__08450_ VGND VGND VPWR VPWR net1090 sky130_fd_sc_hd__inv_2
XFILLER_0_98_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17570_ _05133_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__clkbuf_4
X_14782_ CPU.registerFile\[27\]\[11\] CPU.registerFile\[26\]\[11\] _02768_ VGND VGND
+ VPWR VPWR _02853_ sky130_fd_sc_hd__mux2_1
X_11994_ _06655_ net2372 _07620_ VGND VGND VPWR VPWR _07629_ sky130_fd_sc_hd__mux2_1
X_16521_ _03943_ _04232_ _04235_ _04117_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__a211o_1
X_10945_ _06854_ VGND VGND VPWR VPWR _07001_ sky130_fd_sc_hd__buf_4
XFILLER_0_156_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16452_ _04075_ _04163_ _04168_ _04042_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__o211a_1
X_13664_ clknet_1_0__leaf__08340_ VGND VGND VPWR VPWR _08451_ sky130_fd_sc_hd__buf_1
XFILLER_0_85_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10876_ CPU.aluIn1\[8\] _06946_ _06880_ VGND VGND VPWR VPWR _06947_ sky130_fd_sc_hd__mux2_1
X_15403_ _03450_ _03458_ _03241_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12615_ _06607_ net2371 _07993_ VGND VGND VPWR VPWR _07999_ sky130_fd_sc_hd__mux2_1
X_19171_ clknet_leaf_5_clk _02691_ VGND VGND VPWR VPWR per_uart.uart0.rx_count16\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16383_ _08393_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18122_ net1133 _01650_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_15334_ CPU.registerFile\[19\]\[25\] CPU.registerFile\[18\]\[25\] _03157_ VGND VGND
+ VPWR VPWR _03391_ sky130_fd_sc_hd__mux2_1
X_12546_ _07962_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18053_ net1064 _01581_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15265_ CPU.registerFile\[22\]\[23\] CPU.registerFile\[23\]\[23\] _02998_ VGND VGND
+ VPWR VPWR _03324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12477_ _07925_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__clkbuf_1
X_17004_ CPU.registerFile\[6\]\[24\] CPU.registerFile\[7\]\[24\] _04426_ VGND VGND
+ VPWR VPWR _04707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_4 CPU.mem_wdata\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11428_ _05766_ VGND VGND VPWR VPWR _07314_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1__f__03642_ clknet_0__03642_ VGND VGND VPWR VPWR clknet_1_1__leaf__03642_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15196_ CPU.registerFile\[27\]\[21\] CPU.registerFile\[26\]\[21\] _03172_ VGND VGND
+ VPWR VPWR _03257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11359_ _07276_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__clkbuf_1
X_18955_ net729 _02475_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ net1348 VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__clkbuf_1
X_17906_ clknet_leaf_22_clk _01434_ VGND VGND VPWR VPWR CPU.Jimm\[13\] sky130_fd_sc_hd__dfxtp_4
X_18886_ net660 _02406_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_17837_ net917 _01399_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_17768_ net848 _01330_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16719_ CPU.registerFile\[5\]\[17\] CPU.registerFile\[4\]\[17\] _04428_ VGND VGND
+ VPWR VPWR _04429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17699_ _05207_ _05223_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14146__285 clknet_1_0__leaf__08499_ VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__inv_2
XFILLER_0_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09122_ _05455_ _05458_ _05467_ _05473_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__a211o_1
XFILLER_0_161_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09053_ _05399_ _05404_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold510 CPU.registerFile\[19\]\[28\] VGND VGND VPWR VPWR net1807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold521 CPU.registerFile\[15\]\[18\] VGND VGND VPWR VPWR net1818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 CPU.registerFile\[11\]\[6\] VGND VGND VPWR VPWR net1829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold543 CPU.registerFile\[15\]\[30\] VGND VGND VPWR VPWR net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 CPU.registerFile\[28\]\[31\] VGND VGND VPWR VPWR net1851 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold565 CPU.aluReg\[5\] VGND VGND VPWR VPWR net1862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold576 CPU.registerFile\[17\]\[20\] VGND VGND VPWR VPWR net1873 sky130_fd_sc_hd__dlygate4sd3_1
X_15734__525 clknet_1_0__leaf__03651_ VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__inv_2
Xhold587 CPU.registerFile\[7\]\[18\] VGND VGND VPWR VPWR net1884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 CPU.registerFile\[20\]\[28\] VGND VGND VPWR VPWR net1895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09955_ mapped_spi_ram.rcv_data\[19\] _05685_ _05698_ net1370 VGND VGND VPWR VPWR
+ _06287_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13716__1088 clknet_1_1__leaf__08456_ VGND VGND VPWR VPWR net1144 sky130_fd_sc_hd__inv_2
X_08906_ CPU.aluIn1\[28\] _05257_ VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__nand2_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _05889_ _06220_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__or2_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 CPU.registerFile\[31\]\[2\] VGND VGND VPWR VPWR net2507 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 CPU.registerFile\[24\]\[27\] VGND VGND VPWR VPWR net2518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1232 CPU.registerFile\[14\]\[11\] VGND VGND VPWR VPWR net2529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1243 CPU.aluIn1\[29\] VGND VGND VPWR VPWR net2540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1254 CPU.registerFile\[23\]\[23\] VGND VGND VPWR VPWR net2551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1265 CPU.registerFile\[9\]\[5\] VGND VGND VPWR VPWR net2562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 per_uart.rx_data\[6\] VGND VGND VPWR VPWR net2573 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1287 CPU.aluIn1\[27\] VGND VGND VPWR VPWR net2584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1298 CPU.registerFile\[12\]\[3\] VGND VGND VPWR VPWR net2595 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15628__430 clknet_1_0__leaf__03640_ VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__inv_2
X_10730_ _06815_ VGND VGND VPWR VPWR _06838_ sky130_fd_sc_hd__buf_4
XFILLER_0_138_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10661_ _06800_ VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12400_ net1696 _07309_ _07884_ VGND VGND VPWR VPWR _07885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10592_ net1923 _06316_ _06761_ VGND VGND VPWR VPWR _06763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12331_ _07847_ VGND VGND VPWR VPWR _07848_ sky130_fd_sc_hd__buf_4
XFILLER_0_133_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12262_ net1572 _07799_ _07804_ _07796_ VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15050_ _02750_ _03094_ _03114_ _02839_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__a211o_1
X_11213_ net1630 _07188_ _07195_ VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__a21o_1
Xoutput6 net6 VGND VGND VPWR VPWR TXD sky130_fd_sc_hd__clkbuf_4
X_12193_ net1314 _07692_ _07756_ _07755_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__o211a_1
X_11144_ net1599 _07149_ VGND VGND VPWR VPWR _07154_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18740_ net529 _02264_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[2\] sky130_fd_sc_hd__dfxtp_1
X_11075_ _06992_ _07106_ VGND VGND VPWR VPWR _07107_ sky130_fd_sc_hd__and2_1
X_14251__380 clknet_1_1__leaf__08509_ VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__inv_2
X_14903_ _08764_ _02968_ _02970_ _02814_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__a211o_1
X_10026_ _06354_ _05969_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__xnor2_1
X_18671_ net460 _02195_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_17622_ net1667 per_uart.uart0.rxd_reg\[1\] _05170_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__mux2_1
X_14834_ _08857_ _02900_ _02902_ _02903_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15863__609 clknet_1_1__leaf__03681_ VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__inv_2
XFILLER_0_156_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13733__1103 clknet_1_1__leaf__08458_ VGND VGND VPWR VPWR net1159 sky130_fd_sc_hd__inv_2
X_17553_ _05117_ _05120_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__or2_1
X_14765_ _05861_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__buf_2
XFILLER_0_98_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13357__852 clknet_1_0__leaf__08368_ VGND VGND VPWR VPWR net908 sky130_fd_sc_hd__inv_2
X_11977_ _07597_ VGND VGND VPWR VPWR _07620_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16504_ _04141_ _04200_ _04219_ _04096_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__a211o_1
X_17484_ _05016_ CPU.PC\[11\] _05063_ _05064_ _05053_ VGND VGND VPWR VPWR _02649_
+ sky130_fd_sc_hd__o221a_1
X_10928_ _06973_ _06988_ VGND VGND VPWR VPWR _06989_ sky130_fd_sc_hd__and2_1
X_14696_ CPU.registerFile\[27\]\[9\] CPU.registerFile\[26\]\[9\] _02768_ VGND VGND
+ VPWR VPWR _02769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16435_ CPU.registerFile\[5\]\[10\] CPU.registerFile\[4\]\[10\] _04024_ VGND VGND
+ VPWR VPWR _04152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10859_ CPU.aluIn1\[12\] _06933_ _06914_ VGND VGND VPWR VPWR _06934_ sky130_fd_sc_hd__mux2_1
X_13961__119 clknet_1_1__leaf__08480_ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__inv_2
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19154_ clknet_leaf_4_clk net1464 VGND VGND VPWR VPWR per_uart.uart0.txd_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16366_ _04075_ _04078_ _04084_ _04042_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18105_ net1116 _01633_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15317_ CPU.registerFile\[10\]\[24\] CPU.registerFile\[11\]\[24\] _03183_ VGND VGND
+ VPWR VPWR _03375_ sky130_fd_sc_hd__mux2_1
X_12529_ _07952_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__clkbuf_1
X_19085_ clknet_leaf_0_clk _02605_ VGND VGND VPWR VPWR per_uart.uart0.rxd_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16297_ _08393_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18036_ net1047 _01564_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15248_ _03098_ _03304_ _03306_ _03307_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__a211o_1
XFILLER_0_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15179_ _05861_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__buf_2
XFILLER_0_78_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__03656_ _03656_ VGND VGND VPWR VPWR clknet_0__03656_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09740_ _05912_ _06080_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__nor2_1
X_18938_ net712 _02458_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[19\] sky130_fd_sc_hd__dfxtp_1
.ends

